-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 17:10:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2068\ : std_logic;
signal \VGAClock.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \Pixel_1_RNOZ0Z_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_i\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_i\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_\ : std_logic;
signal \un13_beamx_6_cascade_\ : std_logic;
signal un13_beamx_5 : std_logic;
signal un1_beamylto9_4 : std_logic;
signal \un1_beamylto9_5_cascade_\ : std_logic;
signal \un1_beamy_cascade_\ : std_logic;
signal \VSync_c\ : std_logic;
signal \un11_beamx_3_cascade_\ : std_logic;
signal un11_beamx_6 : std_logic;
signal \un11_beamx_6_cascade_\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum\ : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_\ : std_logic;
signal un5_visiblex_i : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_i\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_axb_6 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\ : std_logic;
signal \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal un4_beamy_cry_1 : std_logic;
signal un4_beamy_cry_2 : std_logic;
signal un4_beamy_cry_3 : std_logic;
signal un4_beamy_cry_4 : std_logic;
signal un4_beamy_cry_5 : std_logic;
signal un4_beamy_cry_6 : std_logic;
signal un4_beamy_cry_7 : std_logic;
signal un4_beamy_cry_8 : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un16_beamx_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un16_beamx_cry_2 : std_logic;
signal un16_beamx_cry_3 : std_logic;
signal un16_beamx_cry_4 : std_logic;
signal un16_beamx_cry_5 : std_logic;
signal un16_beamx_cry_6 : std_logic;
signal un16_beamx_cry_7 : std_logic;
signal un16_beamx_cry_8 : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal un1_beamy : std_logic;
signal un4_beamxlt9 : std_logic;
signal \Pixel_0_sqmuxa_0_cascade_\ : std_logic;
signal un11_beamx_1 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un8_beamxlt9_0 : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \un1_beamxlto9_0_cascade_\ : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal \HSync_c\ : std_logic;
signal \un5_visiblex_cry_7_c_RNIVZ0Z952\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_c5_i\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_c5\ : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal un13_beamx : std_logic;
signal \beamX_RNIVEM1Z0Z_4\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal un5_visibley_cry_0 : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal un5_visibley_cry_1 : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un5_visibley_cry_2 : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal un5_visibley_cry_3 : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum : std_logic;
signal un5_visibley_cry_4 : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum : std_logic;
signal un5_visibley_cry_5 : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum : std_logic;
signal un5_visibley_cry_6 : std_logic;
signal un5_visibley_cry_7 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \un5_visibley_cry_7_c_RNI1L4CZ0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal un5_visibley_cry_8 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_axb_3 : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \un1_beamX_27\ : std_logic;
signal \Pixel_0_sqmuxa_1\ : std_logic;
signal \un13_0_1_cascade_\ : std_logic;
signal un12lt10 : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \Pixel_1_RNOZ0Z_9\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0\ : std_logic;
signal \N_11\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum : std_logic;
signal \un5_visibley_cry_0_c_RNIJVSBZ0\ : std_logic;
signal \G_7_i_a4_0_0\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \VGAClock.PixelClock_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1001010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \VGAClock.PixelClock\,
            REFERENCECLK => \N__2077\,
            RESETB => \N__3789\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4463\,
            DIN => \N__4462\,
            DOUT => \N__4461\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4463\,
            PADOUT => \N__4462\,
            PADIN => \N__4461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4454\,
            DIN => \N__4453\,
            DOUT => \N__4452\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4454\,
            PADOUT => \N__4453\,
            PADIN => \N__4452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4445\,
            DIN => \N__4444\,
            DOUT => \N__4443\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4445\,
            PADOUT => \N__4444\,
            PADIN => \N__4443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4436\,
            DIN => \N__4435\,
            DOUT => \N__4434\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4436\,
            PADOUT => \N__4435\,
            PADIN => \N__4434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3555\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4427\,
            DIN => \N__4426\,
            DOUT => \N__4425\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4427\,
            PADOUT => \N__4426\,
            PADIN => \N__4425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4418\,
            DIN => \N__4417\,
            DOUT => \N__4416\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4418\,
            PADOUT => \N__4417\,
            PADIN => \N__4416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4409\,
            DIN => \N__4408\,
            DOUT => \N__4407\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4409\,
            PADOUT => \N__4408\,
            PADIN => \N__4407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3007\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__957\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4386\
        );

    \I__956\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4383\,
            I => \N__4377\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__4380\,
            I => \N__4374\
        );

    \I__952\ : Span4Mux_s2_h
    port map (
            O => \N__4377\,
            I => \N__4371\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__4374\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum
        );

    \I__950\ : Odrv4
    port map (
            O => \N__4371\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4366\,
            I => \N__4363\
        );

    \I__948\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4360\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49\
        );

    \I__946\ : InMux
    port map (
            O => \N__4357\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__945\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4351\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4351\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4\
        );

    \I__943\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4345\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0\
        );

    \I__941\ : InMux
    port map (
            O => \N__4342\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4339\,
            I => \N__4335\
        );

    \I__939\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4326\
        );

    \I__938\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4326\
        );

    \I__937\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4326\
        );

    \I__936\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4323\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4326\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4323\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__932\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4312\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6\
        );

    \I__930\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4306\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4306\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0\
        );

    \I__928\ : InMux
    port map (
            O => \N__4303\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__927\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4297\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__924\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4288\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4288\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__921\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4279\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__919\ : InMux
    port map (
            O => \N__4276\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__918\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4270\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__916\ : InMux
    port map (
            O => \N__4267\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4264\,
            I => \N__4259\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__4263\,
            I => \N__4255\
        );

    \I__913\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4251\
        );

    \I__912\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4242\
        );

    \I__911\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4242\
        );

    \I__910\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4242\
        );

    \I__909\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4242\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4251\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4242\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0\
        );

    \I__906\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4230\
        );

    \I__904\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4227\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__4230\,
            I => \N__4224\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__901\ : Sp12to4
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__4218\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum
        );

    \I__898\ : Odrv4
    port map (
            O => \N__4215\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__896\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4204\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4201\,
            I => \N__4198\
        );

    \I__893\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__4192\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__890\ : InMux
    port map (
            O => \N__4189\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__889\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__4180\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1\
        );

    \I__886\ : InMux
    port map (
            O => \N__4177\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__884\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__4165\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2\
        );

    \I__881\ : InMux
    port map (
            O => \N__4162\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__880\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__4153\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3\
        );

    \I__877\ : InMux
    port map (
            O => \N__4150\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__876\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4141\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__873\ : InMux
    port map (
            O => \N__4138\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__4135\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__4132\,
            I => \N__4128\
        );

    \I__870\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4116\
        );

    \I__869\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4116\
        );

    \I__868\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4116\
        );

    \I__867\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4116\
        );

    \I__866\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4113\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4113\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__4110\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__861\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4099\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__859\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4093\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__4090\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__856\ : InMux
    port map (
            O => \N__4087\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__855\ : InMux
    port map (
            O => \N__4084\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__854\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4078\,
            I => \Pixel_1_RNOZ0Z_9\
        );

    \I__852\ : InMux
    port map (
            O => \N__4075\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__850\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4066\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4066\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__848\ : InMux
    port map (
            O => \N__4063\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__847\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4057\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11\
        );

    \I__845\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4050\
        );

    \I__844\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4047\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4050\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4047\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4042\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_\
        );

    \I__840\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4035\
        );

    \I__839\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4032\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4035\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4032\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0\
        );

    \I__836\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N_11\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__833\ : InMux
    port map (
            O => \N__4018\,
            I => \N__4015\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4015\,
            I => \N__4010\
        );

    \I__831\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4005\
        );

    \I__830\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4005\
        );

    \I__829\ : Span4Mux_s2_h
    port map (
            O => \N__4010\,
            I => \N__4002\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__3999\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__4002\,
            I => \N__3996\
        );

    \I__826\ : Span4Mux_s2_h
    port map (
            O => \N__3999\,
            I => \N__3993\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__3996\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum
        );

    \I__824\ : Odrv4
    port map (
            O => \N__3993\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum
        );

    \I__823\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3985\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3981\
        );

    \I__821\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3978\
        );

    \I__820\ : Span4Mux_s2_v
    port map (
            O => \N__3981\,
            I => \N__3975\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__3975\,
            I => \N__3969\
        );

    \I__817\ : Span4Mux_s2_h
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__3969\,
            I => \un5_visibley_cry_0_c_RNIJVSBZ0\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__3966\,
            I => \un5_visibley_cry_0_c_RNIJVSBZ0\
        );

    \I__814\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3958\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3958\,
            I => \G_7_i_a4_0_0\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__3955\,
            I => \N__3949\
        );

    \I__811\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3946\
        );

    \I__810\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3943\
        );

    \I__809\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3940\
        );

    \I__808\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3937\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__3946\,
            I => \beamYZ0Z_5\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__3943\,
            I => \beamYZ0Z_5\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3940\,
            I => \beamYZ0Z_5\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__3937\,
            I => \beamYZ0Z_5\
        );

    \I__803\ : InMux
    port map (
            O => \N__3928\,
            I => \N__3922\
        );

    \I__802\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3922\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__3922\,
            I => \N__3919\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__3919\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum
        );

    \I__799\ : InMux
    port map (
            O => \N__3916\,
            I => un5_visibley_cry_4
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__3913\,
            I => \N__3907\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__3912\,
            I => \N__3904\
        );

    \I__796\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3901\
        );

    \I__795\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3898\
        );

    \I__794\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3895\
        );

    \I__793\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3892\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3901\,
            I => \beamYZ0Z_6\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3898\,
            I => \beamYZ0Z_6\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3895\,
            I => \beamYZ0Z_6\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3892\,
            I => \beamYZ0Z_6\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__3883\,
            I => \N__3879\
        );

    \I__787\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3876\
        );

    \I__786\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3873\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3876\,
            I => \N__3868\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__3873\,
            I => \N__3868\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__3868\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum
        );

    \I__782\ : InMux
    port map (
            O => \N__3865\,
            I => un5_visibley_cry_5
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__3862\,
            I => \N__3857\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__3861\,
            I => \N__3853\
        );

    \I__779\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3850\
        );

    \I__778\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3845\
        );

    \I__777\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3845\
        );

    \I__776\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3842\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3850\,
            I => \beamYZ0Z_7\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3845\,
            I => \beamYZ0Z_7\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3842\,
            I => \beamYZ0Z_7\
        );

    \I__772\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3832\,
            I => \N__3828\
        );

    \I__770\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3825\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__3828\,
            I => \N__3822\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3825\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum
        );

    \I__767\ : Odrv4
    port map (
            O => \N__3822\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum
        );

    \I__766\ : InMux
    port map (
            O => \N__3817\,
            I => un5_visibley_cry_6
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__3814\,
            I => \N__3800\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__3813\,
            I => \N__3797\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__3812\,
            I => \N__3794\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__3811\,
            I => \N__3790\
        );

    \I__761\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3781\
        );

    \I__760\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3781\
        );

    \I__759\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3781\
        );

    \I__758\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3778\
        );

    \I__757\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3773\
        );

    \I__756\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3773\
        );

    \I__755\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3770\
        );

    \I__754\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3767\
        );

    \I__753\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3764\
        );

    \I__752\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3757\
        );

    \I__751\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3757\
        );

    \I__750\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3757\
        );

    \I__749\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3754\
        );

    \I__748\ : IoInMux
    port map (
            O => \N__3789\,
            I => \N__3751\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__3788\,
            I => \N__3748\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3781\,
            I => \N__3743\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3734\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3773\,
            I => \N__3734\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3734\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3767\,
            I => \N__3734\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3764\,
            I => \N__3727\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3757\,
            I => \N__3727\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3754\,
            I => \N__3727\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3751\,
            I => \N__3724\
        );

    \I__737\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3721\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__3747\,
            I => \N__3718\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__3746\,
            I => \N__3715\
        );

    \I__734\ : Span4Mux_v
    port map (
            O => \N__3743\,
            I => \N__3708\
        );

    \I__733\ : Span4Mux_v
    port map (
            O => \N__3734\,
            I => \N__3708\
        );

    \I__732\ : Span4Mux_s3_v
    port map (
            O => \N__3727\,
            I => \N__3708\
        );

    \I__731\ : IoSpan4Mux
    port map (
            O => \N__3724\,
            I => \N__3705\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3721\,
            I => \N__3702\
        );

    \I__729\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3697\
        );

    \I__728\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3697\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__3708\,
            I => \CONSTANT_ONE_NET\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__3705\,
            I => \CONSTANT_ONE_NET\
        );

    \I__725\ : Odrv4
    port map (
            O => \N__3702\,
            I => \CONSTANT_ONE_NET\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3697\,
            I => \CONSTANT_ONE_NET\
        );

    \I__723\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3682\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3687\,
            I => \N__3679\
        );

    \I__721\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3676\
        );

    \I__720\ : InMux
    port map (
            O => \N__3685\,
            I => \N__3673\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3682\,
            I => \N__3670\
        );

    \I__718\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3667\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3676\,
            I => \beamYZ0Z_8\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3673\,
            I => \beamYZ0Z_8\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__3670\,
            I => \beamYZ0Z_8\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3667\,
            I => \beamYZ0Z_8\
        );

    \I__713\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3652\
        );

    \I__712\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3652\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3652\,
            I => \N__3649\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__3649\,
            I => \un5_visibley_cry_7_c_RNI1L4CZ0\
        );

    \I__709\ : InMux
    port map (
            O => \N__3646\,
            I => \bfn_9_8_0_\
        );

    \I__708\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3639\
        );

    \I__707\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3634\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3639\,
            I => \N__3631\
        );

    \I__705\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3628\
        );

    \I__704\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3625\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3634\,
            I => \beamYZ0Z_9\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__3631\,
            I => \beamYZ0Z_9\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3628\,
            I => \beamYZ0Z_9\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3625\,
            I => \beamYZ0Z_9\
        );

    \I__699\ : InMux
    port map (
            O => \N__3616\,
            I => un5_visibley_cry_8
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__697\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3604\
        );

    \I__696\ : InMux
    port map (
            O => \N__3609\,
            I => \N__3604\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__3601\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_axb_3
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__3598\,
            I => \N_8_cascade_\
        );

    \I__692\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__690\ : Odrv12
    port map (
            O => \N__3589\,
            I => \un1_beamX_27\
        );

    \I__689\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3583\,
            I => \N__3580\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__3580\,
            I => \Pixel_0_sqmuxa_1\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3577\,
            I => \un13_0_1_cascade_\
        );

    \I__685\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3571\,
            I => \N__3568\
        );

    \I__683\ : Span4Mux_s2_v
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__3565\,
            I => un12lt10
        );

    \I__681\ : IoInMux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__679\ : Span4Mux_s3_v
    port map (
            O => \N__3556\,
            I => \N__3552\
        );

    \I__678\ : IoInMux
    port map (
            O => \N__3555\,
            I => \N__3549\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__3552\,
            I => \N__3546\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3549\,
            I => \N__3543\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__3546\,
            I => \N__3540\
        );

    \I__674\ : Span4Mux_s1_v
    port map (
            O => \N__3543\,
            I => \N__3537\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3540\,
            I => \Pixel_c\
        );

    \I__672\ : Odrv4
    port map (
            O => \N__3537\,
            I => \Pixel_c\
        );

    \I__671\ : ClkMux
    port map (
            O => \N__3532\,
            I => \N__3508\
        );

    \I__670\ : ClkMux
    port map (
            O => \N__3531\,
            I => \N__3508\
        );

    \I__669\ : ClkMux
    port map (
            O => \N__3530\,
            I => \N__3508\
        );

    \I__668\ : ClkMux
    port map (
            O => \N__3529\,
            I => \N__3508\
        );

    \I__667\ : ClkMux
    port map (
            O => \N__3528\,
            I => \N__3508\
        );

    \I__666\ : ClkMux
    port map (
            O => \N__3527\,
            I => \N__3508\
        );

    \I__665\ : ClkMux
    port map (
            O => \N__3526\,
            I => \N__3508\
        );

    \I__664\ : ClkMux
    port map (
            O => \N__3525\,
            I => \N__3508\
        );

    \I__663\ : GlobalMux
    port map (
            O => \N__3508\,
            I => \N__3505\
        );

    \I__662\ : gio2CtrlBuf
    port map (
            O => \N__3505\,
            I => \PixelClock_g\
        );

    \I__661\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3499\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__659\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3490\
        );

    \I__658\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3487\
        );

    \I__657\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3484\
        );

    \I__656\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3481\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3490\,
            I => \N__3476\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3476\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3473\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3481\,
            I => un13_beamx
        );

    \I__651\ : Odrv4
    port map (
            O => \N__3476\,
            I => un13_beamx
        );

    \I__650\ : Odrv4
    port map (
            O => \N__3473\,
            I => un13_beamx
        );

    \I__649\ : CEMux
    port map (
            O => \N__3466\,
            I => \N__3461\
        );

    \I__648\ : CEMux
    port map (
            O => \N__3465\,
            I => \N__3458\
        );

    \I__647\ : CEMux
    port map (
            O => \N__3464\,
            I => \N__3455\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3461\,
            I => \N__3452\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3458\,
            I => \N__3449\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3442\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__3452\,
            I => \N__3437\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__3449\,
            I => \N__3437\
        );

    \I__641\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3432\
        );

    \I__640\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3432\
        );

    \I__639\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3429\
        );

    \I__638\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3426\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__3442\,
            I => \N__3423\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__3437\,
            I => \N__3420\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3432\,
            I => \beamX_RNIVEM1Z0Z_4\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3429\,
            I => \beamX_RNIVEM1Z0Z_4\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3426\,
            I => \beamX_RNIVEM1Z0Z_4\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3423\,
            I => \beamX_RNIVEM1Z0Z_4\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3420\,
            I => \beamX_RNIVEM1Z0Z_4\
        );

    \I__630\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3403\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3408\,
            I => \N__3399\
        );

    \I__628\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3394\
        );

    \I__627\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3394\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3403\,
            I => \N__3391\
        );

    \I__625\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3388\
        );

    \I__624\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3385\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3394\,
            I => \beamYZ0Z_0\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__3391\,
            I => \beamYZ0Z_0\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3388\,
            I => \beamYZ0Z_0\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3385\,
            I => \beamYZ0Z_0\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3376\,
            I => \N__3371\
        );

    \I__618\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3368\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \N__3363\
        );

    \I__616\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3360\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3368\,
            I => \N__3357\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3367\,
            I => \N__3354\
        );

    \I__613\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3351\
        );

    \I__612\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3348\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3360\,
            I => \N__3343\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__3357\,
            I => \N__3343\
        );

    \I__609\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3340\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3351\,
            I => \beamYZ0Z_1\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3348\,
            I => \beamYZ0Z_1\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__3343\,
            I => \beamYZ0Z_1\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3340\,
            I => \beamYZ0Z_1\
        );

    \I__604\ : InMux
    port map (
            O => \N__3331\,
            I => un5_visibley_cry_0
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3328\,
            I => \N__3322\
        );

    \I__602\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3319\
        );

    \I__601\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3314\
        );

    \I__600\ : InMux
    port map (
            O => \N__3325\,
            I => \N__3314\
        );

    \I__599\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3311\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3319\,
            I => \beamYZ0Z_2\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3314\,
            I => \beamYZ0Z_2\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3311\,
            I => \beamYZ0Z_2\
        );

    \I__595\ : InMux
    port map (
            O => \N__3304\,
            I => un5_visibley_cry_1
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__3301\,
            I => \N__3295\
        );

    \I__593\ : InMux
    port map (
            O => \N__3300\,
            I => \N__3292\
        );

    \I__592\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3287\
        );

    \I__591\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3287\
        );

    \I__590\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3284\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3292\,
            I => \beamYZ0Z_3\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3287\,
            I => \beamYZ0Z_3\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3284\,
            I => \beamYZ0Z_3\
        );

    \I__586\ : InMux
    port map (
            O => \N__3277\,
            I => un5_visibley_cry_2
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__3274\,
            I => \N__3268\
        );

    \I__584\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3265\
        );

    \I__583\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3262\
        );

    \I__582\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3259\
        );

    \I__581\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3256\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3265\,
            I => \beamYZ0Z_4\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3262\,
            I => \beamYZ0Z_4\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3259\,
            I => \beamYZ0Z_4\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3256\,
            I => \beamYZ0Z_4\
        );

    \I__576\ : InMux
    port map (
            O => \N__3247\,
            I => un5_visibley_cry_3
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__3244\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\
        );

    \I__574\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3238\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\
        );

    \I__572\ : InMux
    port map (
            O => \N__3235\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__570\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3226\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1\
        );

    \I__568\ : InMux
    port map (
            O => \N__3223\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__567\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3217\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1\
        );

    \I__565\ : InMux
    port map (
            O => \N__3214\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__564\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3208\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3208\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1\
        );

    \I__562\ : InMux
    port map (
            O => \N__3205\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__561\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3199\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__559\ : InMux
    port map (
            O => \N__3196\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3193\,
            I => \N__3188\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3192\,
            I => \N__3184\
        );

    \I__556\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3180\
        );

    \I__555\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3171\
        );

    \I__554\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3171\
        );

    \I__553\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3171\
        );

    \I__552\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3171\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3180\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3171\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1\
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__3166\,
            I => \N__3163\
        );

    \I__548\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3160\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3160\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__3157\,
            I => \N__3152\
        );

    \I__545\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3147\
        );

    \I__544\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3140\
        );

    \I__543\ : InMux
    port map (
            O => \N__3152\,
            I => \N__3140\
        );

    \I__542\ : InMux
    port map (
            O => \N__3151\,
            I => \N__3140\
        );

    \I__541\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3137\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3147\,
            I => \beamXZ0Z_9\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3140\,
            I => \beamXZ0Z_9\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3137\,
            I => \beamXZ0Z_9\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__3130\,
            I => \N__3123\
        );

    \I__536\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3119\
        );

    \I__535\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3116\
        );

    \I__534\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3109\
        );

    \I__533\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3109\
        );

    \I__532\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3109\
        );

    \I__531\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3106\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3119\,
            I => \beamXZ0Z_7\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3116\,
            I => \beamXZ0Z_7\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3109\,
            I => \beamXZ0Z_7\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3106\,
            I => \beamXZ0Z_7\
        );

    \I__526\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3089\
        );

    \I__525\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3084\
        );

    \I__524\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3084\
        );

    \I__523\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3079\
        );

    \I__522\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3079\
        );

    \I__521\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3076\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3089\,
            I => \beamXZ0Z_6\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3084\,
            I => \beamXZ0Z_6\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3079\,
            I => \beamXZ0Z_6\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3076\,
            I => \beamXZ0Z_6\
        );

    \I__516\ : InMux
    port map (
            O => \N__3067\,
            I => \N__3060\
        );

    \I__515\ : InMux
    port map (
            O => \N__3066\,
            I => \N__3057\
        );

    \I__514\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3052\
        );

    \I__513\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3052\
        );

    \I__512\ : InMux
    port map (
            O => \N__3063\,
            I => \N__3049\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3060\,
            I => \beamXZ0Z_8\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3057\,
            I => \beamXZ0Z_8\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3052\,
            I => \beamXZ0Z_8\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3049\,
            I => \beamXZ0Z_8\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3040\,
            I => \un1_beamxlto9_0_cascade_\
        );

    \I__506\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3029\
        );

    \I__505\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3024\
        );

    \I__504\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3024\
        );

    \I__503\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3019\
        );

    \I__502\ : InMux
    port map (
            O => \N__3033\,
            I => \N__3019\
        );

    \I__501\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3016\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3029\,
            I => \beamXZ0Z_5\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3024\,
            I => \beamXZ0Z_5\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3019\,
            I => \beamXZ0Z_5\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3016\,
            I => \beamXZ0Z_5\
        );

    \I__496\ : IoInMux
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3004\,
            I => \N__3001\
        );

    \I__494\ : Span4Mux_s2_v
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__493\ : Span4Mux_v
    port map (
            O => \N__2998\,
            I => \N__2995\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__2995\,
            I => \N__2991\
        );

    \I__491\ : IoInMux
    port map (
            O => \N__2994\,
            I => \N__2988\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__2991\,
            I => \N__2985\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2982\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__2985\,
            I => \HSync_c\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__2982\,
            I => \HSync_c\
        );

    \I__486\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2973\
        );

    \I__485\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2970\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2973\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2970\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__482\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2962\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2962\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_c5_i\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__2959\,
            I => \N__2956\
        );

    \I__479\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2953\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__2953\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\
        );

    \I__477\ : InMux
    port map (
            O => \N__2950\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__2947\,
            I => \N__2944\
        );

    \I__475\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2941\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2941\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575\
        );

    \I__473\ : InMux
    port map (
            O => \N__2938\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__2935\,
            I => \N__2932\
        );

    \I__471\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2929\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\
        );

    \I__469\ : InMux
    port map (
            O => \N__2926\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__468\ : InMux
    port map (
            O => \N__2923\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\
        );

    \I__467\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2915\
        );

    \I__466\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2910\
        );

    \I__465\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2910\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2915\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_c5\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2910\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_c5\
        );

    \I__462\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2902\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\
        );

    \I__460\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2895\
        );

    \I__459\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2892\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2895\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2892\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__456\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2883\
        );

    \I__455\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2880\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2883\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2880\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\
        );

    \I__452\ : InMux
    port map (
            O => \N__2875\,
            I => un16_beamx_cry_4
        );

    \I__451\ : InMux
    port map (
            O => \N__2872\,
            I => un16_beamx_cry_5
        );

    \I__450\ : InMux
    port map (
            O => \N__2869\,
            I => un16_beamx_cry_6
        );

    \I__449\ : InMux
    port map (
            O => \N__2866\,
            I => un16_beamx_cry_7
        );

    \I__448\ : InMux
    port map (
            O => \N__2863\,
            I => \bfn_9_2_0_\
        );

    \I__447\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2857\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__445\ : Span4Mux_s2_v
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__444\ : Span4Mux_v
    port map (
            O => \N__2851\,
            I => \N__2848\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__2848\,
            I => un1_beamy
        );

    \I__442\ : InMux
    port map (
            O => \N__2845\,
            I => \N__2842\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2842\,
            I => un4_beamxlt9
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__2839\,
            I => \Pixel_0_sqmuxa_0_cascade_\
        );

    \I__439\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2832\
        );

    \I__438\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2829\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2832\,
            I => un11_beamx_1
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2829\,
            I => un11_beamx_1
        );

    \I__435\ : InMux
    port map (
            O => \N__2824\,
            I => \N__2816\
        );

    \I__434\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2811\
        );

    \I__433\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2811\
        );

    \I__432\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2808\
        );

    \I__431\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2803\
        );

    \I__430\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2803\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2816\,
            I => \beamXZ0Z_4\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2811\,
            I => \beamXZ0Z_4\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2808\,
            I => \beamXZ0Z_4\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2803\,
            I => \beamXZ0Z_4\
        );

    \I__425\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2791\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2791\,
            I => un8_beamxlt9_0
        );

    \I__423\ : InMux
    port map (
            O => \N__2788\,
            I => un4_beamy_cry_5
        );

    \I__422\ : InMux
    port map (
            O => \N__2785\,
            I => un4_beamy_cry_6
        );

    \I__421\ : InMux
    port map (
            O => \N__2782\,
            I => un4_beamy_cry_7
        );

    \I__420\ : InMux
    port map (
            O => \N__2779\,
            I => \bfn_8_8_0_\
        );

    \I__419\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2770\
        );

    \I__418\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2763\
        );

    \I__417\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2763\
        );

    \I__416\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2763\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2770\,
            I => \beamXZ0Z_0\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2763\,
            I => \beamXZ0Z_0\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__412\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2750\
        );

    \I__411\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2745\
        );

    \I__410\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2745\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2750\,
            I => \beamXZ0Z_1\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2745\,
            I => \beamXZ0Z_1\
        );

    \I__407\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2736\
        );

    \I__406\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2733\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2736\,
            I => \beamXZ0Z_2\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2733\,
            I => \beamXZ0Z_2\
        );

    \I__403\ : InMux
    port map (
            O => \N__2728\,
            I => un16_beamx_cry_1
        );

    \I__402\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2722\,
            I => \N__2718\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__2721\,
            I => \N__2714\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__2718\,
            I => \N__2711\
        );

    \I__398\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2708\
        );

    \I__397\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2705\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__2711\,
            I => \beamXZ0Z_3\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2708\,
            I => \beamXZ0Z_3\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2705\,
            I => \beamXZ0Z_3\
        );

    \I__393\ : InMux
    port map (
            O => \N__2698\,
            I => un16_beamx_cry_2
        );

    \I__392\ : InMux
    port map (
            O => \N__2695\,
            I => un16_beamx_cry_3
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__2692\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__2689\,
            I => \N__2684\
        );

    \I__389\ : InMux
    port map (
            O => \N__2688\,
            I => \N__2681\
        );

    \I__388\ : InMux
    port map (
            O => \N__2687\,
            I => \N__2678\
        );

    \I__387\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2675\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2681\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2678\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2675\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__383\ : InMux
    port map (
            O => \N__2668\,
            I => \N__2665\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2665\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__381\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2659\,
            I => \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__2656\,
            I => \N__2653\
        );

    \I__378\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2650\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2650\,
            I => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\
        );

    \I__376\ : InMux
    port map (
            O => \N__2647\,
            I => un4_beamy_cry_1
        );

    \I__375\ : InMux
    port map (
            O => \N__2644\,
            I => un4_beamy_cry_2
        );

    \I__374\ : InMux
    port map (
            O => \N__2641\,
            I => un4_beamy_cry_3
        );

    \I__373\ : InMux
    port map (
            O => \N__2638\,
            I => un4_beamy_cry_4
        );

    \I__372\ : InMux
    port map (
            O => \N__2635\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__371\ : CascadeMux
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__370\ : InMux
    port map (
            O => \N__2629\,
            I => \N__2626\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2626\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0\
        );

    \I__368\ : InMux
    port map (
            O => \N__2623\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__367\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2617\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2617\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0\
        );

    \I__365\ : InMux
    port map (
            O => \N__2614\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__364\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2607\
        );

    \I__363\ : InMux
    port map (
            O => \N__2610\,
            I => \N__2604\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2607\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2604\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__359\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2593\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2593\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1\
        );

    \I__357\ : InMux
    port map (
            O => \N__2590\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__356\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2584\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2581\,
            I => \N__2576\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2580\,
            I => \N__2573\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2579\,
            I => \N__2569\
        );

    \I__351\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2560\
        );

    \I__350\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2560\
        );

    \I__349\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2560\
        );

    \I__348\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2560\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2560\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0\
        );

    \I__346\ : InMux
    port map (
            O => \N__2557\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__345\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2551\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2551\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\
        );

    \I__343\ : InMux
    port map (
            O => \N__2548\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__342\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2542\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\
        );

    \I__340\ : InMux
    port map (
            O => \N__2539\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__339\ : InMux
    port map (
            O => \N__2536\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__338\ : InMux
    port map (
            O => \N__2533\,
            I => \N__2530\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2530\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__336\ : InMux
    port map (
            O => \N__2527\,
            I => \N__2524\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2524\,
            I => \N__2520\
        );

    \I__334\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2517\
        );

    \I__333\ : Span4Mux_v
    port map (
            O => \N__2520\,
            I => \N__2514\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2517\,
            I => \N__2511\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__2514\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__2511\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum\
        );

    \I__329\ : InMux
    port map (
            O => \N__2506\,
            I => \N__2503\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2503\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__2500\,
            I => \N__2497\
        );

    \I__326\ : InMux
    port map (
            O => \N__2497\,
            I => \N__2494\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2494\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_i\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2491\,
            I => \N__2488\
        );

    \I__323\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2485\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2485\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731\
        );

    \I__321\ : InMux
    port map (
            O => \N__2482\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__320\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2476\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2476\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__2473\,
            I => \N__2470\
        );

    \I__317\ : InMux
    port map (
            O => \N__2470\,
            I => \N__2467\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2467\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1\
        );

    \I__315\ : InMux
    port map (
            O => \N__2464\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__314\ : InMux
    port map (
            O => \N__2461\,
            I => \N__2458\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2458\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\
        );

    \I__312\ : InMux
    port map (
            O => \N__2455\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__311\ : InMux
    port map (
            O => \N__2452\,
            I => \N__2449\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2449\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\
        );

    \I__309\ : InMux
    port map (
            O => \N__2446\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\
        );

    \I__308\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2439\
        );

    \I__307\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2436\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2439\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2436\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2431\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_\
        );

    \I__303\ : InMux
    port map (
            O => \N__2428\,
            I => \N__2422\
        );

    \I__302\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2422\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2422\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2419\,
            I => \N__2415\
        );

    \I__299\ : InMux
    port map (
            O => \N__2418\,
            I => \N__2410\
        );

    \I__298\ : InMux
    port map (
            O => \N__2415\,
            I => \N__2410\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2410\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\
        );

    \I__296\ : CascadeMux
    port map (
            O => \N__2407\,
            I => \N__2403\
        );

    \I__295\ : InMux
    port map (
            O => \N__2406\,
            I => \N__2399\
        );

    \I__294\ : InMux
    port map (
            O => \N__2403\,
            I => \N__2394\
        );

    \I__293\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2394\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2399\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2394\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0\
        );

    \I__290\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2386\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2386\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2383\,
            I => \N__2379\
        );

    \I__287\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2374\
        );

    \I__286\ : InMux
    port map (
            O => \N__2379\,
            I => \N__2371\
        );

    \I__285\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2366\
        );

    \I__284\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2366\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2374\,
            I => un5_visiblex_i
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2371\,
            I => un5_visiblex_i
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2366\,
            I => un5_visiblex_i
        );

    \I__280\ : InMux
    port map (
            O => \N__2359\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__279\ : InMux
    port map (
            O => \N__2356\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__278\ : InMux
    port map (
            O => \N__2353\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__277\ : InMux
    port map (
            O => \N__2350\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__2347\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_\
        );

    \I__275\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2338\
        );

    \I__274\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2338\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2338\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__271\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2329\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2329\,
            I => un5_visiblex_i_24
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2326\,
            I => \N__2323\
        );

    \I__268\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2319\
        );

    \I__267\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2316\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2313\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2316\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum\
        );

    \I__264\ : Odrv4
    port map (
            O => \N__2313\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum\
        );

    \I__263\ : InMux
    port map (
            O => \N__2308\,
            I => un5_visiblex_cry_4
        );

    \I__262\ : InMux
    port map (
            O => \N__2305\,
            I => un5_visiblex_cry_5
        );

    \I__261\ : InMux
    port map (
            O => \N__2302\,
            I => un5_visiblex_cry_6
        );

    \I__260\ : InMux
    port map (
            O => \N__2299\,
            I => un5_visiblex_cry_7
        );

    \I__259\ : InMux
    port map (
            O => \N__2296\,
            I => un5_visiblex_cry_8
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__2293\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2290\,
            I => \un13_beamx_6_cascade_\
        );

    \I__256\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2284\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2284\,
            I => un13_beamx_5
        );

    \I__254\ : InMux
    port map (
            O => \N__2281\,
            I => \N__2278\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2278\,
            I => un1_beamylto9_4
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2275\,
            I => \un1_beamylto9_5_cascade_\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2272\,
            I => \un1_beamy_cascade_\
        );

    \I__250\ : IoInMux
    port map (
            O => \N__2269\,
            I => \N__2266\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2266\,
            I => \N__2263\
        );

    \I__248\ : Span4Mux_s2_v
    port map (
            O => \N__2263\,
            I => \N__2259\
        );

    \I__247\ : IoInMux
    port map (
            O => \N__2262\,
            I => \N__2256\
        );

    \I__246\ : Span4Mux_h
    port map (
            O => \N__2259\,
            I => \N__2253\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2256\,
            I => \N__2250\
        );

    \I__244\ : Span4Mux_v
    port map (
            O => \N__2253\,
            I => \N__2247\
        );

    \I__243\ : Span4Mux_s2_v
    port map (
            O => \N__2250\,
            I => \N__2244\
        );

    \I__242\ : Odrv4
    port map (
            O => \N__2247\,
            I => \VSync_c\
        );

    \I__241\ : Odrv4
    port map (
            O => \N__2244\,
            I => \VSync_c\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2239\,
            I => \un11_beamx_3_cascade_\
        );

    \I__239\ : InMux
    port map (
            O => \N__2236\,
            I => \N__2233\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2233\,
            I => un11_beamx_6
        );

    \I__237\ : CascadeMux
    port map (
            O => \N__2230\,
            I => \un11_beamx_6_cascade_\
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__2227\,
            I => \N__2224\
        );

    \I__235\ : InMux
    port map (
            O => \N__2224\,
            I => \N__2221\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2221\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_i\
        );

    \I__233\ : InMux
    port map (
            O => \N__2218\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__232\ : InMux
    port map (
            O => \N__2215\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__231\ : InMux
    port map (
            O => \N__2212\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__230\ : InMux
    port map (
            O => \N__2209\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__229\ : InMux
    port map (
            O => \N__2206\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__2203\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_\
        );

    \I__227\ : InMux
    port map (
            O => \N__2200\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\
        );

    \I__226\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2194\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2194\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57\
        );

    \I__224\ : CascadeMux
    port map (
            O => \N__2191\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_\
        );

    \I__223\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2184\
        );

    \I__222\ : InMux
    port map (
            O => \N__2187\,
            I => \N__2181\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2184\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2181\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__2176\,
            I => \N__2173\
        );

    \I__218\ : InMux
    port map (
            O => \N__2173\,
            I => \N__2170\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2170\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_i\
        );

    \I__216\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2164\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2164\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1\
        );

    \I__214\ : InMux
    port map (
            O => \N__2161\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__213\ : CascadeMux
    port map (
            O => \N__2158\,
            I => \N__2155\
        );

    \I__212\ : InMux
    port map (
            O => \N__2155\,
            I => \N__2152\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2152\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2\
        );

    \I__210\ : InMux
    port map (
            O => \N__2149\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__209\ : InMux
    port map (
            O => \N__2146\,
            I => \N__2143\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__2143\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\
        );

    \I__207\ : InMux
    port map (
            O => \N__2140\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__206\ : InMux
    port map (
            O => \N__2137\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\
        );

    \I__205\ : CascadeMux
    port map (
            O => \N__2134\,
            I => \N__2130\
        );

    \I__204\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2126\
        );

    \I__203\ : InMux
    port map (
            O => \N__2130\,
            I => \N__2121\
        );

    \I__202\ : InMux
    port map (
            O => \N__2129\,
            I => \N__2121\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2126\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2121\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3\
        );

    \I__199\ : InMux
    port map (
            O => \N__2116\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__198\ : InMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2110\,
            I => \Pixel_1_RNOZ0Z_6\
        );

    \I__196\ : InMux
    port map (
            O => \N__2107\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\
        );

    \I__195\ : InMux
    port map (
            O => \N__2104\,
            I => \N__2098\
        );

    \I__194\ : InMux
    port map (
            O => \N__2103\,
            I => \N__2098\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__2098\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\
        );

    \I__192\ : IoInMux
    port map (
            O => \N__2095\,
            I => \N__2092\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__2092\,
            I => \N__2089\
        );

    \I__190\ : Span4Mux_s1_h
    port map (
            O => \N__2089\,
            I => \N__2086\
        );

    \I__189\ : Span4Mux_h
    port map (
            O => \N__2086\,
            I => \N__2083\
        );

    \I__188\ : Sp12to4
    port map (
            O => \N__2083\,
            I => \N__2080\
        );

    \I__187\ : Odrv12
    port map (
            O => \N__2080\,
            I => \VGAClock.PixelClock\
        );

    \I__186\ : IoInMux
    port map (
            O => \N__2077\,
            I => \N__2074\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__2074\,
            I => \N__2071\
        );

    \I__184\ : IoSpan4Mux
    port map (
            O => \N__2071\,
            I => \N__2068\
        );

    \I__183\ : Odrv4
    port map (
            O => \N__2068\,
            I => \Clock12MHz_c\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visibley_cry_7,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_beamy_cry_8,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un16_beamx_cry_8,
            carryinitout => \bfn_9_2_0_\
        );

    \VGAClock.PLLOUTCORE_derived_clock_RNIE579\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2095\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__2187\,
            in1 => \N__2113\,
            in2 => \N__2383\,
            in3 => \N__2197\,
            lcout => \un1_beamX_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2377\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2103\,
            in2 => \N__2176\,
            in3 => \N__2116\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_6_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2167\,
            in2 => \N__2134\,
            in3 => \N__2107\,
            lcout => \Pixel_1_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2104\,
            in2 => \N__2158\,
            in3 => \N__2129\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCR57_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2146\,
            in2 => \_gnd_net_\,
            in3 => \N__2200\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57\,
            ltout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_2_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110101000000"
        )
    port map (
            in0 => \N__2378\,
            in1 => \N__2725\,
            in2 => \N__2191\,
            in3 => \N__2188\,
            lcout => un12lt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2322\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2326\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRM1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2427\,
            in2 => \N__2227\,
            in3 => \N__2161\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1O2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2443\,
            in2 => \N__2491\,
            in3 => \N__2149\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIG1IT6_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2133\,
            in1 => \N__2428\,
            in2 => \N__2473\,
            in3 => \N__2140\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3P3_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2461\,
            in2 => \_gnd_net_\,
            in3 => \N__2137\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2527\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3835\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6O_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2662\,
            in2 => \N__3746\,
            in3 => \N__2218\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3U_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2554\,
            in2 => \N__3788\,
            in3 => \N__2215\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5U_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2545\,
            in2 => \N__3747\,
            in3 => \N__2212\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2689\,
            in3 => \N__2209\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883I_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2533\,
            in2 => \_gnd_net_\,
            in3 => \N__2206\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0\,
            ltout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29G1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__2611\,
            in1 => \_gnd_net_\,
            in2 => \N__2203\,
            in3 => \_gnd_net_\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIB625_9_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3953\,
            in1 => \N__3272\,
            in2 => \N__3376\,
            in3 => \N__3643\,
            lcout => OPEN,
            ltout => \un13_beamx_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2287\,
            in1 => \N__3409\,
            in2 => \N__2290\,
            in3 => \N__3685\,
            lcout => un13_beamx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIA525_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3326\,
            in1 => \N__3910\,
            in2 => \N__3862\,
            in3 => \N__3299\,
            lcout => un13_beamx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJNP3_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3688\,
            in1 => \N__3856\,
            in2 => \_gnd_net_\,
            in3 => \N__3325\,
            lcout => un1_beamylto9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3271\,
            in1 => \N__3298\,
            in2 => \N__3913\,
            in3 => \N__3375\,
            lcout => OPEN,
            ltout => \un1_beamylto9_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0DB_9_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2281\,
            in1 => \N__3638\,
            in2 => \N__2275\,
            in3 => \N__3952\,
            lcout => un1_beamy,
            ltout => \un1_beamy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2272\,
            in3 => \_gnd_net_\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIG3M_5_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3036\,
            in1 => \N__2835\,
            in2 => \_gnd_net_\,
            in3 => \N__3096\,
            lcout => OPEN,
            ltout => \un11_beamx_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_4_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2236\,
            in1 => \N__3128\,
            in2 => \N__2239\,
            in3 => \N__2823\,
            lcout => \beamX_RNIVEM1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2739\,
            in1 => \N__2753\,
            in2 => \N__2721\,
            in3 => \N__2773\,
            lcout => un11_beamx_6,
            ltout => \un11_beamx_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_5_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010101"
        )
    port map (
            in0 => \N__3095\,
            in1 => \N__3035\,
            in2 => \N__2230\,
            in3 => \N__2822\,
            lcout => un4_beamxlt9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2754\,
            in2 => \_gnd_net_\,
            in3 => \N__2775\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3529\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2819\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3032\,
            in2 => \N__3814\,
            in3 => \N__2308\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3092\,
            in2 => \N__3812\,
            in3 => \N__2305\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3122\,
            in2 => \_gnd_net_\,
            in3 => \N__2302\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3063\,
            in2 => \N__3813\,
            in3 => \N__2299\,
            lcout => \un5_visiblex_cry_7_c_RNIVZ0Z952\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_7,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3150\,
            in2 => \_gnd_net_\,
            in3 => \N__2296\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_c5\,
            ltout => \un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2293\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_c5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2820\,
            in1 => \N__3793\,
            in2 => \_gnd_net_\,
            in3 => \N__2382\,
            lcout => un5_visiblex_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2343\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2899\,
            in2 => \N__2335\,
            in3 => \N__2359\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2886\,
            in2 => \N__2959\,
            in3 => \N__2356\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6C831_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2406\,
            in1 => \N__3241\,
            in2 => \N__2947\,
            in3 => \N__2353\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2887\,
            in1 => \N__2920\,
            in2 => \N__2935\,
            in3 => \N__2350\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0\,
            ltout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2347\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2344\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2523\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISM731_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2506\,
            in2 => \N__2500\,
            in3 => \N__2482\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJF1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2479\,
            in2 => \N__2407\,
            in3 => \N__2464\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5E1N3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2442\,
            in1 => \N__2389\,
            in2 => \N__2419\,
            in3 => \N__2455\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2452\,
            in2 => \_gnd_net_\,
            in3 => \N__2446\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1\,
            ltout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2431\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI48631_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__2418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2402\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453A1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2668\,
            in2 => \N__2579\,
            in3 => \N__2635\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTO1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2572\,
            in2 => \N__2632\,
            in3 => \N__2623\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRU1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2620\,
            in2 => \N__2580\,
            in3 => \N__2614\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNI894A4_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3191\,
            in1 => \N__2610\,
            in2 => \N__2599\,
            in3 => \N__2590\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2587\,
            in1 => \N__2687\,
            in2 => \N__2581\,
            in3 => \N__2557\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3657\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3803\,
            in2 => \N__2656\,
            in3 => \N__2548\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3804\,
            in2 => \N__3613\,
            in3 => \N__2539\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2536\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2692\,
            in3 => \N__2688\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3831\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_7_c_RNI1L4C_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3658\,
            lcout => \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3609\,
            lcout => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_beamy_cry_1_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3402\,
            in2 => \N__3374\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => un4_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3493\,
            in1 => \N__3327\,
            in2 => \_gnd_net_\,
            in3 => \N__2647\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => un4_beamy_cry_1,
            carryout => un4_beamy_cry_2,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3300\,
            in2 => \_gnd_net_\,
            in3 => \N__2644\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => un4_beamy_cry_2,
            carryout => un4_beamy_cry_3,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3273\,
            in2 => \_gnd_net_\,
            in3 => \N__2641\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un4_beamy_cry_3,
            carryout => un4_beamy_cry_4,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3954\,
            in2 => \_gnd_net_\,
            in3 => \N__2638\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un4_beamy_cry_4,
            carryout => un4_beamy_cry_5,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3911\,
            in2 => \_gnd_net_\,
            in3 => \N__2788\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un4_beamy_cry_5,
            carryout => un4_beamy_cry_6,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3496\,
            in1 => \N__3860\,
            in2 => \_gnd_net_\,
            in3 => \N__2785\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => un4_beamy_cry_6,
            carryout => un4_beamy_cry_7,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3686\,
            in2 => \_gnd_net_\,
            in3 => \N__2782\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un4_beamy_cry_7,
            carryout => un4_beamy_cry_8,
            clk => \N__3527\,
            ce => \N__3466\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3642\,
            in1 => \N__3495\,
            in2 => \_gnd_net_\,
            in3 => \N__2779\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3526\,
            ce => \N__3465\,
            sr => \_gnd_net_\
        );

    \un16_beamx_cry_1_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2776\,
            in2 => \N__2758\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => un16_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2740\,
            in2 => \_gnd_net_\,
            in3 => \N__2728\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un16_beamx_cry_1,
            carryout => un16_beamx_cry_2,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2717\,
            in2 => \_gnd_net_\,
            in3 => \N__2698\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un16_beamx_cry_2,
            carryout => un16_beamx_cry_3,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2824\,
            in2 => \_gnd_net_\,
            in3 => \N__2695\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un16_beamx_cry_3,
            carryout => un16_beamx_cry_4,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3037\,
            in2 => \_gnd_net_\,
            in3 => \N__2875\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un16_beamx_cry_4,
            carryout => un16_beamx_cry_5,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3447\,
            in1 => \N__3097\,
            in2 => \_gnd_net_\,
            in3 => \N__2872\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un16_beamx_cry_5,
            carryout => un16_beamx_cry_6,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3445\,
            in1 => \N__3129\,
            in2 => \_gnd_net_\,
            in3 => \N__2869\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un16_beamx_cry_6,
            carryout => un16_beamx_cry_7,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3448\,
            in1 => \N__3066\,
            in2 => \_gnd_net_\,
            in3 => \N__2866\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un16_beamx_cry_7,
            carryout => un16_beamx_cry_8,
            clk => \N__3531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3156\,
            in1 => \N__3446\,
            in2 => \_gnd_net_\,
            in3 => \N__2863\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_4_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__3065\,
            in1 => \N__2794\,
            in2 => \N__3157\,
            in3 => \N__2860\,
            lcout => OPEN,
            ltout => \Pixel_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__2845\,
            in1 => \N__2836\,
            in2 => \N__2839\,
            in3 => \N__3126\,
            lcout => \Pixel_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3151\,
            in2 => \_gnd_net_\,
            in3 => \N__3064\,
            lcout => un11_beamx_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_10_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__3093\,
            in1 => \N__3033\,
            in2 => \N__3130\,
            in3 => \N__2821\,
            lcout => un8_beamxlt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_RNO_0_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3155\,
            in2 => \_gnd_net_\,
            in3 => \N__3127\,
            lcout => OPEN,
            ltout => \un1_beamxlto9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__3094\,
            in1 => \N__3067\,
            in2 => \N__3040\,
            in3 => \N__3034\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2976\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2965\,
            in2 => \_gnd_net_\,
            in3 => \N__2950\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNI1575_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2905\,
            in2 => \N__3811\,
            in3 => \N__2938\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2919\,
            in2 => \_gnd_net_\,
            in3 => \N__2926\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2923\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2918\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2898\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\,
            ltout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3244\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3927\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQ1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3502\,
            in2 => \N__3192\,
            in3 => \N__3235\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTR2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3187\,
            in2 => \N__3232\,
            in3 => \N__3223\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPA3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3220\,
            in2 => \N__3193\,
            in3 => \N__3214\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMVQV7_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4125\,
            in1 => \N__3211\,
            in2 => \N__3166\,
            in3 => \N__3205\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3202\,
            in2 => \_gnd_net_\,
            in3 => \N__3196\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_0_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3882\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3494\,
            in2 => \_gnd_net_\,
            in3 => \N__3406\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3528\,
            ce => \N__3464\,
            sr => \_gnd_net_\
        );

    \beamY_1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3366\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3528\,
            ce => \N__3464\,
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_0_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3408\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => un5_visibley_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_0_c_RNIJVSB_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3367\,
            in3 => \N__3331\,
            lcout => \un5_visibley_cry_0_c_RNIJVSBZ0\,
            ltout => OPEN,
            carryin => un5_visibley_cry_0,
            carryout => un5_visibley_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_1_c_RNIL2UB_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3808\,
            in2 => \N__3328\,
            in3 => \N__3304\,
            lcout => un1_visibley_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_1,
            carryout => un5_visibley_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_2_c_RNIN5VB_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3805\,
            in2 => \N__3301\,
            in3 => \N__3277\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_2,
            carryout => un5_visibley_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_3_c_RNIP80C_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3809\,
            in2 => \N__3274\,
            in3 => \N__3247\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_3,
            carryout => un5_visibley_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_4_c_RNIRB1C_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3955\,
            in3 => \N__3916\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_4,
            carryout => un5_visibley_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_5_c_RNITE2C_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3810\,
            in2 => \N__3912\,
            in3 => \N__3865\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_5,
            carryout => un5_visibley_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_6_c_RNIVH3C_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3806\,
            in2 => \N__3861\,
            in3 => \N__3817\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_6,
            carryout => un5_visibley_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_7_c_RNI1L4C_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3807\,
            in2 => \N__3687\,
            in3 => \N__3646\,
            lcout => \un5_visibley_cry_7_c_RNI1L4CZ0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => un5_visibley_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3637\,
            in2 => \_gnd_net_\,
            in3 => \N__3616\,
            lcout => un1_visibley_if_generate_plus_mult1_un33_sum_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_7_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4053\,
            in1 => \N__4038\,
            in2 => \N__4021\,
            in3 => \N__4060\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_3_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__3988\,
            in1 => \N__4081\,
            in2 => \N__3598\,
            in3 => \N__4027\,
            lcout => OPEN,
            ltout => \un13_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000100"
        )
    port map (
            in0 => \N__3595\,
            in1 => \N__3586\,
            in2 => \N__3577\,
            in3 => \N__3574\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4013\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCH_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4096\,
            in2 => \N__4263\,
            in3 => \N__4087\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6Q_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4258\,
            in2 => \N__4366\,
            in3 => \N__4084\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_9_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4348\,
            in2 => \N__4264\,
            in3 => \N__4075\,
            lcout => \Pixel_1_RNOZ0Z_9\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4309\,
            in2 => \N__4072\,
            in3 => \N__4254\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDG11_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4285\,
            in3 => \N__4063\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11\,
            ltout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_8_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3961\,
            in1 => \N__4054\,
            in2 => \N__4042\,
            in3 => \N__4039\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_11_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3984\,
            lcout => \G_7_i_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4233\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGS4_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4127\,
            in2 => \N__4201\,
            in3 => \N__4189\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEK6_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4186\,
            in2 => \N__4132\,
            in3 => \N__4177\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3M7_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4131\,
            in2 => \N__4174\,
            in3 => \N__4162\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNI2S0GG_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__4159\,
            in2 => \N__4105\,
            in3 => \N__4150\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4147\,
            in2 => \_gnd_net_\,
            in3 => \N__4138\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8\,
            ltout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_0_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4135\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_0_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4126\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4390\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4389\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMR49_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4334\,
            in2 => \N__4210\,
            in3 => \N__4357\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LD_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4354\,
            in2 => \N__4339\,
            in3 => \N__4342\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DF_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4338\,
            in2 => \N__4318\,
            in3 => \N__4303\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIG8GC11_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4262\,
            in1 => \N__4300\,
            in2 => \N__4294\,
            in3 => \N__4276\,
            lcout => un1_visibley_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTG_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4273\,
            in2 => \_gnd_net_\,
            in3 => \N__4267\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4237\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
