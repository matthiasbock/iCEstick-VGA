-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 23 2015 21:38:03

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal r_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal r_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal r_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal r_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal r_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s_0 : std_logic;
signal r_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \r_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal r_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal r_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s_0 : std_logic;
signal r_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \r_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal r_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal r_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal if_generate_plus_mult1_un47_sum_cry_3_s : std_logic;
signal r_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \r_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal r_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal r_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \visibleYZ0Z_6\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_\ : std_logic;
signal \visibleYZ0Z_7\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal \visibleY_RNINQ3DZ0Z_8\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \G_251\ : std_logic;
signal r_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal \G_252\ : std_logic;
signal r_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal r_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal \G_250\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal r_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal r_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal r_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s_0 : std_logic;
signal \r_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal r_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \r_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal r_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal r_if_generate_plus_mult1_un75_sum : std_logic;
signal un5_vy_cry_0 : std_logic;
signal r_if_generate_plus_mult1_un68_sum : std_logic;
signal un5_vy_cry_1 : std_logic;
signal r_if_generate_plus_mult1_un61_sum : std_logic;
signal un5_vy_cry_2 : std_logic;
signal un5_vy_cry_3 : std_logic;
signal un5_vy_cry_4 : std_logic;
signal un5_vy_cry_5 : std_logic;
signal un5_vy_cry_6 : std_logic;
signal if_generate_plus_mult1_un61_sum_s_5 : std_logic;
signal if_generate_plus_mult1_un68_sum_s_5 : std_logic;
signal r_if_generate_plus_mult1_un54_sum : std_logic;
signal r_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal r_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5_0 : std_logic;
signal un7_r_1 : std_logic;
signal r_if_generate_plus_mult1_un47_sum : std_logic;
signal r_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \un5_vy_cry_6_c_RNIG9KKZ0\ : std_logic;
signal if_generate_plus_mult1_un47_sum_axb_4_l_ofx : std_logic;
signal \un5_vy_cry_6_c_RNI9MAAZ0\ : std_logic;
signal \N_7_i\ : std_logic;
signal if_generate_plus_mult1_un47_sum_s_5 : std_logic;
signal r_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal \un5_vy_cry_5_c_RNI7J9AZ0\ : std_logic;
signal un5_vy_i_24 : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_\ : std_logic;
signal \visibleYZ0Z_4\ : std_logic;
signal \visibleYZ0Z_5\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal \visibleYZ0Z_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6 : std_logic;
signal \visibleYZ0Z_9\ : std_logic;
signal \visibleY_RNIOR3DZ0Z_9\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \c_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal c_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal c_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal c_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal c_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal c_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal c_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \c_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal c_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal c_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_0_THRU_CO\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_1_THRU_CO\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_2_THRU_CO\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_3_THRU_CO\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_5_THRU_CO\ : std_logic;
signal \un21_beamy_cry_1_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal if_generate_plus_mult1_un82_sum_s_5 : std_logic;
signal un7_r_4 : std_logic;
signal if_generate_plus_mult1_un75_sum_s_5 : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11\ : std_logic;
signal \Pixel_RNOZ0Z_7\ : std_logic;
signal \visibleYZ0Z_3\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97\ : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal un5_vx_cry_0 : std_logic;
signal un5_vx_cry_1 : std_logic;
signal un5_vx_cry_2 : std_logic;
signal c_if_generate_plus_mult1_un61_sum : std_logic;
signal un5_vx_cry_3 : std_logic;
signal un5_vx_cry_4 : std_logic;
signal un5_vx_cry_5 : std_logic;
signal un5_vx_cry_6 : std_logic;
signal un5_vx_cry_7 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal un5_vx_cry_8 : std_logic;
signal \CO3_0_cascade_\ : std_logic;
signal \N_14\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal c_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal c_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal c_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \G_253\ : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal c_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal un9_r_0lto2 : std_logic;
signal \c_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal c_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un9_r_1lt6_0 : std_logic;
signal c_if_generate_plus_mult1_un68_sum : std_logic;
signal \c_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal un9_r_0lto3 : std_logic;
signal un9_r_0lto3_i : std_logic;
signal \N_404_i\ : std_logic;
signal c_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal \beamY_RNI9DLCZ0Z_2\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal un5_beamx_5 : std_logic;
signal \un1_beamy_4_cascade_\ : std_logic;
signal un5_beamx_3 : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal un1_beamy_4 : std_logic;
signal un8_beamy_2 : std_logic;
signal \un1_beamylto9_2_cascade_\ : std_logic;
signal \VSync_c\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \un4_beamylt8_0_cascade_\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un5_vy : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal un8_beamylto9_1 : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41\ : std_logic;
signal \Pixel_RNOZ0Z_5_cascade_\ : std_logic;
signal \N_45_cascade_\ : std_logic;
signal \N_76\ : std_logic;
signal \TextOutputEnabledZ0\ : std_logic;
signal \N_74_i_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \INVPixelZ0C_net\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0\ : std_logic;
signal \visibleYZ0Z_1\ : std_logic;
signal \visibleYZ0Z_2\ : std_logic;
signal \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0\ : std_logic;
signal \Pixel_RNOZ0Z_6\ : std_logic;
signal \un13_beamylt7_cascade_\ : std_logic;
signal \OutputEnabledZ0\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \un18_beamylto9_2_cascade_\ : std_logic;
signal un8_beamy : std_logic;
signal \un18_beamylt10_0_cascade_\ : std_logic;
signal un4_beamy_0 : std_logic;
signal un15_beamy_2 : std_logic;
signal un13_beamylt7 : std_logic;
signal \un15_beamy_2_cascade_\ : std_logic;
signal \beamX_RNISO4TZ0Z_7\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \un5_vx_i_25_cascade_\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal un5_vx_i_0_25 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_1_cry_1 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_axb_5_i : std_logic;
signal \N_13_0_i\ : std_logic;
signal c_if_generate_plus_mult1_un47_sum_1_cry_2 : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx : std_logic;
signal c_if_generate_plus_mult1_un47_sum_1_cry_3 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_1_cry_4 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_0 : std_logic;
signal c_if_generate_plus_mult1_un47_sum1_4 : std_logic;
signal \N_18_cascade_\ : std_logic;
signal c_if_generate_plus_mult1_un47_sum1_3 : std_logic;
signal c_if_generate_plus_mult1_un47_sum1_5 : std_logic;
signal c_if_generate_plus_mult1_un47_sum1_0 : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_2_l_fx : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal c_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_3_l_fx : std_logic;
signal if_generate_plus_mult1_un47_sum_m_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal c_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \N_18\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_4_l_fx : std_logic;
signal \c_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal c_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \c_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal c_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5 : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \N_84\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_\ : std_logic;
signal \N_53\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0\ : std_logic;
signal \Pixel_RNOZ0Z_8\ : std_logic;
signal \visibleXZ0Z_4\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0\ : std_logic;
signal \N_81\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \un3_beamx_5_cascade_\ : std_logic;
signal un5_vx : std_logic;
signal \un3_beamx_7_cascade_\ : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal c_if_generate_plus_mult1_un47_sum_1 : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx : std_logic;
signal un5_vx_i_25 : std_logic;
signal c_if_generate_plus_mult1_un47_sum0_2 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_cry_1 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_cry_3_ma : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx : std_logic;
signal c_if_generate_plus_mult1_un47_sum0_3 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_cry_2 : std_logic;
signal \N_186_0_i\ : std_logic;
signal c_if_generate_plus_mult1_un47_sum0_4 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_cry_3 : std_logic;
signal c_if_generate_plus_mult1_un47_sum_0_cry_4 : std_logic;
signal c_if_generate_plus_mult1_un47_sum0_5 : std_logic;
signal \un5_vx_cry_6_c_RNI59BZ0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \N_3_0\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx : std_logic;
signal \visibleXZ0Z_8\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \visibleXZ0Z_5\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08\ : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un1_beamx_2 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \HSync_c\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \visibleXZ0Z_6\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \visibleXZ0Z_7\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \CO3_0\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal un15_beamy_g : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7 : std_logic;
signal \visibleXZ0Z_9\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0\ : std_logic;
signal \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_\ : std_logic;
signal chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8 : std_logic;
signal \G_255_cascade_\ : std_logic;
signal \G_256\ : std_logic;
signal \CharacterDisplay__decfrac8\ : std_logic;
signal \G_255\ : std_logic;
signal \G_254\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__3688\,
            RESETB => \N__7752\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7874\,
            DIN => \N__7873\,
            DOUT => \N__7872\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7874\,
            PADOUT => \N__7873\,
            PADIN => \N__7872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7533\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7865\,
            DIN => \N__7864\,
            DOUT => \N__7863\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7865\,
            PADOUT => \N__7864\,
            PADIN => \N__7863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7856\,
            DIN => \N__7855\,
            DOUT => \N__7854\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7856\,
            PADOUT => \N__7855\,
            PADIN => \N__7854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7092\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7847\,
            DIN => \N__7846\,
            DOUT => \N__7845\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7847\,
            PADOUT => \N__7846\,
            PADIN => \N__7845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7838\,
            DIN => \N__7837\,
            DOUT => \N__7836\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7838\,
            PADOUT => \N__7837\,
            PADIN => \N__7836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7099\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7829\,
            DIN => \N__7828\,
            DOUT => \N__7827\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7829\,
            PADOUT => \N__7828\,
            PADIN => \N__7827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5386\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7820\,
            DIN => \N__7819\,
            DOUT => \N__7818\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7820\,
            PADOUT => \N__7819\,
            PADIN => \N__7818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1699\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7795\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7795\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7795\,
            I => \visibleXZ0Z_9\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7786\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__7783\,
            I => \N__7775\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__7782\,
            I => \N__7771\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__7781\,
            I => \N__7763\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__7780\,
            I => \N__7760\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__7779\,
            I => \N__7757\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__7778\,
            I => \N__7754\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7749\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7774\,
            I => \N__7744\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7744\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7741\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__7769\,
            I => \N__7737\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__7768\,
            I => \N__7732\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__7767\,
            I => \N__7728\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__7766\,
            I => \N__7724\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7720\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7715\
        );

    \I__1677\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7715\
        );

    \I__1676\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7710\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7710\
        );

    \I__1674\ : IoInMux
    port map (
            O => \N__7752\,
            I => \N__7707\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7749\,
            I => \N__7697\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7744\,
            I => \N__7697\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7741\,
            I => \N__7694\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7691\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7686\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7686\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7671\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7671\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7671\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7671\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7727\,
            I => \N__7671\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7671\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7671\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7720\,
            I => \N__7664\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7715\,
            I => \N__7664\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7664\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7707\,
            I => \N__7661\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7658\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__7705\,
            I => \N__7655\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__7704\,
            I => \N__7652\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__7703\,
            I => \N__7649\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__7702\,
            I => \N__7646\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__7697\,
            I => \N__7643\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__7694\,
            I => \N__7636\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7636\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7686\,
            I => \N__7636\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7633\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__7664\,
            I => \N__7630\
        );

    \I__1645\ : IoSpan4Mux
    port map (
            O => \N__7661\,
            I => \N__7625\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7658\,
            I => \N__7625\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7620\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7620\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7615\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7615\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7643\,
            I => \N__7612\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__7636\,
            I => \N__7607\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__7633\,
            I => \N__7607\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__7630\,
            I => \N__7598\
        );

    \I__1635\ : Span4Mux_s3_v
    port map (
            O => \N__7625\,
            I => \N__7598\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7620\,
            I => \N__7598\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7615\,
            I => \N__7598\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__7612\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__7607\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__7598\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__7591\,
            I => \N__7588\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7585\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7582\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__1625\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7573\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7573\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__7570\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7561\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7561\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7561\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__7558\,
            I => \G_255_cascade_\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7549\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7549\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7549\,
            I => \G_256\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__7534\,
            I => \N__7530\
        );

    \I__1609\ : IoInMux
    port map (
            O => \N__7533\,
            I => \N__7527\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__7530\,
            I => \CharacterDisplay__decfrac8\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7527\,
            I => \CharacterDisplay__decfrac8\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7513\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7513\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7513\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7513\,
            I => \G_255\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7501\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7501\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7501\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7501\,
            I => \G_254\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__7498\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7492\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7492\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__1595\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7485\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7482\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7485\,
            I => \visibleXZ0Z_7\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7482\,
            I => \visibleXZ0Z_7\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7471\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__1588\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7463\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7460\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__7466\,
            I => \N__7451\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7444\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7460\,
            I => \N__7444\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7441\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7423\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7423\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7423\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7423\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7423\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7420\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7415\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7415\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__7444\,
            I => \N__7410\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7410\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7405\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7405\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7398\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7398\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7398\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7395\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7392\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7423\,
            I => \CO3_0\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7420\,
            I => \CO3_0\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7415\,
            I => \CO3_0\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__7410\,
            I => \CO3_0\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7405\,
            I => \CO3_0\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7398\,
            I => \CO3_0\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7395\,
            I => \CO3_0\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7392\,
            I => \CO3_0\
        );

    \I__1557\ : ClkMux
    port map (
            O => \N__7375\,
            I => \N__7306\
        );

    \I__1556\ : ClkMux
    port map (
            O => \N__7374\,
            I => \N__7306\
        );

    \I__1555\ : ClkMux
    port map (
            O => \N__7373\,
            I => \N__7306\
        );

    \I__1554\ : ClkMux
    port map (
            O => \N__7372\,
            I => \N__7306\
        );

    \I__1553\ : ClkMux
    port map (
            O => \N__7371\,
            I => \N__7306\
        );

    \I__1552\ : ClkMux
    port map (
            O => \N__7370\,
            I => \N__7306\
        );

    \I__1551\ : ClkMux
    port map (
            O => \N__7369\,
            I => \N__7306\
        );

    \I__1550\ : ClkMux
    port map (
            O => \N__7368\,
            I => \N__7306\
        );

    \I__1549\ : ClkMux
    port map (
            O => \N__7367\,
            I => \N__7306\
        );

    \I__1548\ : ClkMux
    port map (
            O => \N__7366\,
            I => \N__7306\
        );

    \I__1547\ : ClkMux
    port map (
            O => \N__7365\,
            I => \N__7306\
        );

    \I__1546\ : ClkMux
    port map (
            O => \N__7364\,
            I => \N__7306\
        );

    \I__1545\ : ClkMux
    port map (
            O => \N__7363\,
            I => \N__7306\
        );

    \I__1544\ : ClkMux
    port map (
            O => \N__7362\,
            I => \N__7306\
        );

    \I__1543\ : ClkMux
    port map (
            O => \N__7361\,
            I => \N__7306\
        );

    \I__1542\ : ClkMux
    port map (
            O => \N__7360\,
            I => \N__7306\
        );

    \I__1541\ : ClkMux
    port map (
            O => \N__7359\,
            I => \N__7306\
        );

    \I__1540\ : ClkMux
    port map (
            O => \N__7358\,
            I => \N__7306\
        );

    \I__1539\ : ClkMux
    port map (
            O => \N__7357\,
            I => \N__7306\
        );

    \I__1538\ : ClkMux
    port map (
            O => \N__7356\,
            I => \N__7306\
        );

    \I__1537\ : ClkMux
    port map (
            O => \N__7355\,
            I => \N__7306\
        );

    \I__1536\ : ClkMux
    port map (
            O => \N__7354\,
            I => \N__7306\
        );

    \I__1535\ : ClkMux
    port map (
            O => \N__7353\,
            I => \N__7306\
        );

    \I__1534\ : GlobalMux
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__1533\ : gio2CtrlBuf
    port map (
            O => \N__7303\,
            I => \PixelClock_g\
        );

    \I__1532\ : CEMux
    port map (
            O => \N__7300\,
            I => \N__7258\
        );

    \I__1531\ : CEMux
    port map (
            O => \N__7299\,
            I => \N__7258\
        );

    \I__1530\ : CEMux
    port map (
            O => \N__7298\,
            I => \N__7258\
        );

    \I__1529\ : CEMux
    port map (
            O => \N__7297\,
            I => \N__7258\
        );

    \I__1528\ : CEMux
    port map (
            O => \N__7296\,
            I => \N__7258\
        );

    \I__1527\ : CEMux
    port map (
            O => \N__7295\,
            I => \N__7258\
        );

    \I__1526\ : CEMux
    port map (
            O => \N__7294\,
            I => \N__7258\
        );

    \I__1525\ : CEMux
    port map (
            O => \N__7293\,
            I => \N__7258\
        );

    \I__1524\ : CEMux
    port map (
            O => \N__7292\,
            I => \N__7258\
        );

    \I__1523\ : CEMux
    port map (
            O => \N__7291\,
            I => \N__7258\
        );

    \I__1522\ : CEMux
    port map (
            O => \N__7290\,
            I => \N__7258\
        );

    \I__1521\ : CEMux
    port map (
            O => \N__7289\,
            I => \N__7258\
        );

    \I__1520\ : CEMux
    port map (
            O => \N__7288\,
            I => \N__7258\
        );

    \I__1519\ : CEMux
    port map (
            O => \N__7287\,
            I => \N__7258\
        );

    \I__1518\ : GlobalMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1517\ : gio2CtrlBuf
    port map (
            O => \N__7255\,
            I => un15_beamy_g
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7246\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7243\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7234\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7234\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7231\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__1508\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7225\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7222\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__1505\ : InMux
    port map (
            O => \N__7219\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7
        );

    \I__1504\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7213\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7213\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7207\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7206\,
            I => \N__7198\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7195\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7192\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__7201\,
            I => \N__7189\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7186\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7183\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7192\,
            I => \beamXZ0Z_10\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__7189\,
            I => \beamXZ0Z_10\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7186\,
            I => \beamXZ0Z_10\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__7183\,
            I => \beamXZ0Z_10\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7171\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__1488\ : Span4Mux_h
    port map (
            O => \N__7168\,
            I => \N__7162\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7159\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7154\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7154\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__7162\,
            I => un1_beamx_2
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7159\,
            I => un1_beamx_2
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7154\,
            I => un1_beamx_2
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7132\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7129\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7126\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7119\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7119\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7119\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7116\
        );

    \I__1472\ : Odrv12
    port map (
            O => \N__7132\,
            I => \beamXZ0Z_7\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7129\,
            I => \beamXZ0Z_7\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7126\,
            I => \beamXZ0Z_7\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7119\,
            I => \beamXZ0Z_7\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7116\,
            I => \beamXZ0Z_7\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7105\,
            I => \N__7102\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7102\,
            I => un1_beamxlt10_0
        );

    \I__1465\ : IoInMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1463\ : IoSpan4Mux
    port map (
            O => \N__7093\,
            I => \N__7089\
        );

    \I__1462\ : IoInMux
    port map (
            O => \N__7092\,
            I => \N__7086\
        );

    \I__1461\ : Span4Mux_s2_v
    port map (
            O => \N__7089\,
            I => \N__7083\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7080\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7083\,
            I => \N__7075\
        );

    \I__1458\ : Span12Mux_s1_v
    port map (
            O => \N__7080\,
            I => \N__7075\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__7075\,
            I => \HSync_c\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7066\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__1453\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7059\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7056\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7059\,
            I => \visibleXZ0Z_6\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7056\,
            I => \visibleXZ0Z_6\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7048\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7045\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1446\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7038\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7035\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7038\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7035\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7024\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__7021\,
            I => \N__7017\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7012\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7012\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7012\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7009\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__1434\ : InMux
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7005\,
            I => \N__7000\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7000\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6991\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6985\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6985\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__1426\ : InMux
    port map (
            O => \N__6982\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__1425\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6976\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__1423\ : InMux
    port map (
            O => \N__6973\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__6970\,
            I => \N__6966\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6962\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6957\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6957\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6962\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6957\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__6952\,
            I => \N__6949\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6946\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6946\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6943\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__1412\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6937\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6937\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__1410\ : InMux
    port map (
            O => \N__6934\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__1409\ : InMux
    port map (
            O => \N__6931\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__1408\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6923\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6918\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6918\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6923\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6918\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6907\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6907\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__1400\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6900\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6897\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6892\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6897\,
            I => \N__6892\
        );

    \I__1396\ : Span4Mux_h
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__6889\,
            I => \visibleXZ0Z_5\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6883\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__6880\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6877\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__6874\,
            I => \N__6871\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6868\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6868\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6865\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__1386\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6859\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__1384\ : InMux
    port map (
            O => \N__6856\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__1383\ : InMux
    port map (
            O => \N__6853\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__6850\,
            I => \N__6846\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6842\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6837\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6837\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6842\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6837\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6832\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1375\ : InMux
    port map (
            O => \N__6829\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__1374\ : InMux
    port map (
            O => \N__6826\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__1373\ : InMux
    port map (
            O => \N__6823\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__6820\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__6817\,
            I => \N__6814\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__6811\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__1368\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6804\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6797\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6794\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6785\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6785\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6801\,
            I => \N__6785\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6785\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N_3_0\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__6794\,
            I => \N_3_0\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N_3_0\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6775\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6775\,
            I => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx
        );

    \I__1356\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6768\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6765\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6768\,
            I => \visibleXZ0Z_8\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6765\,
            I => \visibleXZ0Z_8\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__6760\,
            I => \N__6757\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6754\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6754\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6751\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__6748\,
            I => \N__6740\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6737\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6732\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6732\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6727\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6727\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6724\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6737\,
            I => \beamXZ0Z_6\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6732\,
            I => \beamXZ0Z_6\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6727\,
            I => \beamXZ0Z_6\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6724\,
            I => \beamXZ0Z_6\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6707\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6702\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6702\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6697\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6711\,
            I => \N__6697\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6694\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6707\,
            I => \beamXZ0Z_4\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6702\,
            I => \beamXZ0Z_4\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6697\,
            I => \beamXZ0Z_4\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6694\,
            I => \beamXZ0Z_4\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__6685\,
            I => \N__6680\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__6684\,
            I => \N__6675\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6683\,
            I => \N__6671\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6666\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6666\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6661\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6661\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6658\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6671\,
            I => \beamXZ0Z_5\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6666\,
            I => \beamXZ0Z_5\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6661\,
            I => \beamXZ0Z_5\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6658\,
            I => \beamXZ0Z_5\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \N__6643\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6639\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6634\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6634\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6631\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6628\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6639\,
            I => \beamXZ0Z_3\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6634\,
            I => \beamXZ0Z_3\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6631\,
            I => \beamXZ0Z_3\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6628\,
            I => \beamXZ0Z_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6611\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6611\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6605\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6605\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6611\,
            I => \N__6602\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6599\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6605\,
            I => \N__6596\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__6602\,
            I => c_if_generate_plus_mult1_un47_sum_1
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6599\,
            I => c_if_generate_plus_mult1_un47_sum_1
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__6596\,
            I => c_if_generate_plus_mult1_un47_sum_1
        );

    \I__1295\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6586\,
            I => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6577\,
            I => un5_vx_i_25
        );

    \I__1290\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1288\ : Span4Mux_h
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6565\,
            I => c_if_generate_plus_mult1_un47_sum0_2
        );

    \I__1286\ : InMux
    port map (
            O => \N__6562\,
            I => c_if_generate_plus_mult1_un47_sum_0_cry_1
        );

    \I__1285\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6556\,
            I => if_generate_plus_mult1_un47_sum_0_cry_3_ma
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__6553\,
            I => \N__6550\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6547\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6547\,
            I => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx
        );

    \I__1280\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6541\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6541\,
            I => \N__6538\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__6538\,
            I => c_if_generate_plus_mult1_un47_sum0_3
        );

    \I__1277\ : InMux
    port map (
            O => \N__6535\,
            I => c_if_generate_plus_mult1_un47_sum_0_cry_2
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__6532\,
            I => \N__6529\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6526\,
            I => \N_186_0_i\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6517\,
            I => c_if_generate_plus_mult1_un47_sum0_4
        );

    \I__1270\ : InMux
    port map (
            O => \N__6514\,
            I => c_if_generate_plus_mult1_un47_sum_0_cry_3
        );

    \I__1269\ : InMux
    port map (
            O => \N__6511\,
            I => c_if_generate_plus_mult1_un47_sum_0_cry_4
        );

    \I__1268\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6505\,
            I => \N__6500\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6495\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6495\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__6500\,
            I => \N__6492\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6489\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__6492\,
            I => c_if_generate_plus_mult1_un47_sum0_5
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__6489\,
            I => c_if_generate_plus_mult1_un47_sum0_5
        );

    \I__1260\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6471\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6468\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6465\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6460\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6460\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6453\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6453\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6453\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__6471\,
            I => \un5_vx_cry_6_c_RNI59BZ0\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6468\,
            I => \un5_vx_cry_6_c_RNI59BZ0\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6465\,
            I => \un5_vx_cry_6_c_RNI59BZ0\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6460\,
            I => \un5_vx_cry_6_c_RNI59BZ0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6453\,
            I => \un5_vx_cry_6_c_RNI59BZ0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6436\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6436\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6436\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__1243\ : InMux
    port map (
            O => \N__6433\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__1242\ : InMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6427\,
            I => \N__6424\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__6421\,
            I => \N_84\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__6418\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N_53\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6405\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6402\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6405\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6402\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6394\,
            I => \Pixel_RNOZ0Z_8\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6379\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6379\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6379\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6370\,
            I => \visibleXZ0Z_4\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6364\,
            I => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N_81\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6349\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__1214\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6340\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6337\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6334\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6331\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6340\,
            I => \beamXZ0Z_2\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6337\,
            I => \beamXZ0Z_2\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6334\,
            I => \beamXZ0Z_2\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6331\,
            I => \beamXZ0Z_2\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6315\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6310\
        );

    \I__1203\ : Span4Mux_v
    port map (
            O => \N__6315\,
            I => \N__6307\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6304\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6301\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6310\,
            I => \beamXZ0Z_1\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__6307\,
            I => \beamXZ0Z_1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6304\,
            I => \beamXZ0Z_1\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6301\,
            I => \beamXZ0Z_1\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__6292\,
            I => \un3_beamx_5_cascade_\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__6289\,
            I => \N__6285\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6278\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6275\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6272\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6269\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6264\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6281\,
            I => \N__6264\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6278\,
            I => un5_vx
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6275\,
            I => un5_vx
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6272\,
            I => un5_vx
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6269\,
            I => un5_vx
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6264\,
            I => un5_vx
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__6253\,
            I => \un3_beamx_7_cascade_\
        );

    \I__1182\ : CEMux
    port map (
            O => \N__6250\,
            I => \N__6245\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6240\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6240\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6245\,
            I => \N__6236\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6231\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6228\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__6236\,
            I => \N__6225\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6220\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6220\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6231\,
            I => \N__6217\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6228\,
            I => \N__6212\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__6225\,
            I => \N__6212\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6220\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__6217\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__6212\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6199\,
            I => if_generate_plus_mult1_un54_sum_axb_2_l_fx
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6190\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__6187\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__1160\ : InMux
    port map (
            O => \N__6184\,
            I => c_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__1159\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6178\,
            I => if_generate_plus_mult1_un54_sum_axb_3_l_fx
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6168\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6165\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6162\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6165\,
            I => if_generate_plus_mult1_un47_sum_m_2
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6162\,
            I => if_generate_plus_mult1_un47_sum_m_2
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__6148\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__1147\ : InMux
    port map (
            O => \N__6145\,
            I => c_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__6142\,
            I => \N__6138\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__6141\,
            I => \N__6135\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6130\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6127\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6122\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6122\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N_18\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6127\,
            I => \N_18\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N_18\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6109\,
            I => if_generate_plus_mult1_un54_sum_axb_4_l_fx
        );

    \I__1134\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__6100\,
            I => \c_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6097\,
            I => c_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__1130\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6091\,
            I => \c_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6088\,
            I => c_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1127\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__1125\ : Span4Mux_v
    port map (
            O => \N__6079\,
            I => \N__6075\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6072\
        );

    \I__1123\ : Span4Mux_v
    port map (
            O => \N__6075\,
            I => \N__6065\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6072\,
            I => \N__6065\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6062\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6059\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6065\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6062\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6059\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1116\ : InMux
    port map (
            O => \N__6052\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1115\ : InMux
    port map (
            O => \N__6049\,
            I => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__1114\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6043\,
            I => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx
        );

    \I__1112\ : InMux
    port map (
            O => \N__6040\,
            I => c_if_generate_plus_mult1_un47_sum_1_cry_3
        );

    \I__1111\ : InMux
    port map (
            O => \N__6037\,
            I => c_if_generate_plus_mult1_un47_sum_1_cry_4
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__6034\,
            I => \N__6030\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6021\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6021\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6018\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6011\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6011\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6011\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6021\,
            I => c_if_generate_plus_mult1_un47_sum_0_0
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6018\,
            I => c_if_generate_plus_mult1_un47_sum_0_0
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6011\,
            I => c_if_generate_plus_mult1_un47_sum_0_0
        );

    \I__1100\ : InMux
    port map (
            O => \N__6004\,
            I => \N__6001\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6001\,
            I => c_if_generate_plus_mult1_un47_sum1_4
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__5998\,
            I => \N_18_cascade_\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5995\,
            I => \N__5992\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5992\,
            I => c_if_generate_plus_mult1_un47_sum1_3
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5989\,
            I => \N__5985\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5981\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5976\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5976\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5981\,
            I => c_if_generate_plus_mult1_un47_sum1_5
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5976\,
            I => c_if_generate_plus_mult1_un47_sum1_5
        );

    \I__1089\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5966\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5961\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5961\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5956\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5956\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__5956\,
            I => c_if_generate_plus_mult1_un47_sum1_0
        );

    \I__1083\ : InMux
    port map (
            O => \N__5953\,
            I => un8_beamx_cry_9
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__5950\,
            I => \un5_vx_i_25_cascade_\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5941\,
            I => un5_vx_i_0_25
        );

    \I__1078\ : InMux
    port map (
            O => \N__5938\,
            I => c_if_generate_plus_mult1_un47_sum_1_cry_1
        );

    \I__1077\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5932\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5932\,
            I => c_if_generate_plus_mult1_un47_sum_0_axb_5_i
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5923\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5923\,
            I => \N_13_0_i\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5920\,
            I => c_if_generate_plus_mult1_un47_sum_1_cry_2
        );

    \I__1071\ : InMux
    port map (
            O => \N__5917\,
            I => un8_beamx_cry_1
        );

    \I__1070\ : InMux
    port map (
            O => \N__5914\,
            I => un8_beamx_cry_2
        );

    \I__1069\ : InMux
    port map (
            O => \N__5911\,
            I => un8_beamx_cry_3
        );

    \I__1068\ : InMux
    port map (
            O => \N__5908\,
            I => un8_beamx_cry_4
        );

    \I__1067\ : InMux
    port map (
            O => \N__5905\,
            I => un8_beamx_cry_5
        );

    \I__1066\ : InMux
    port map (
            O => \N__5902\,
            I => un8_beamx_cry_6
        );

    \I__1065\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5890\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5885\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5885\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5893\,
            I => \N__5882\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5890\,
            I => \beamXZ0Z_8\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5885\,
            I => \beamXZ0Z_8\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__5882\,
            I => \beamXZ0Z_8\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5875\,
            I => un8_beamx_cry_7
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5872\,
            I => \N__5868\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5862\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5862\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5858\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5862\,
            I => \N__5855\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5852\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5858\,
            I => \beamXZ0Z_9\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__5855\,
            I => \beamXZ0Z_9\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5852\,
            I => \beamXZ0Z_9\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5845\,
            I => \bfn_7_9_0_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5837\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5832\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5832\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5837\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5832\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5818\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1037\ : Span4Mux_v
    port map (
            O => \N__5815\,
            I => \N__5812\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__5812\,
            I => \visibleYZ0Z_1\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__5809\,
            I => \N__5803\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5798\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5807\,
            I => \N__5798\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5806\,
            I => \N__5795\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5792\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5789\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5795\,
            I => \visibleYZ0Z_2\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5792\,
            I => \visibleYZ0Z_2\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__5789\,
            I => \visibleYZ0Z_2\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5777\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5774\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5771\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5768\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5774\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5771\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5768\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5758\,
            I => \Pixel_RNOZ0Z_6\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \un13_beamylt7_cascade_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5749\,
            I => \OutputEnabledZ0\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5740\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__5737\,
            I => un18_beamylt4
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__5734\,
            I => \un18_beamylto9_2_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__5725\,
            I => un8_beamy
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__5722\,
            I => \un18_beamylt10_0_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__5713\,
            I => un4_beamy_0
        );

    \I__1002\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5707\,
            I => un15_beamy_2
        );

    \I__1000\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5701\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5701\,
            I => un13_beamylt7
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__5698\,
            I => \un15_beamy_2_cascade_\
        );

    \I__997\ : IoInMux
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__995\ : Span4Mux_s2_h
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__5683\,
            I => \beamX_RNISO4TZ0Z_7\
        );

    \I__992\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__991\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5671\
        );

    \I__990\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5668\
        );

    \I__989\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5665\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5674\,
            I => \beamYZ0Z_6\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5671\,
            I => \beamYZ0Z_6\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5668\,
            I => \beamYZ0Z_6\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5665\,
            I => \beamYZ0Z_6\
        );

    \I__984\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5650\
        );

    \I__983\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5647\
        );

    \I__982\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5644\
        );

    \I__981\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5641\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5650\,
            I => \beamYZ0Z_5\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5647\,
            I => \beamYZ0Z_5\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5644\,
            I => \beamYZ0Z_5\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5641\,
            I => \beamYZ0Z_5\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \un4_beamylt6_cascade_\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5629\,
            I => \N__5624\
        );

    \I__974\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5619\
        );

    \I__973\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5616\
        );

    \I__972\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5611\
        );

    \I__971\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5611\
        );

    \I__970\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5608\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5619\,
            I => \beamYZ0Z_9\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5616\,
            I => \beamYZ0Z_9\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5611\,
            I => \beamYZ0Z_9\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5608\,
            I => \beamYZ0Z_9\
        );

    \I__965\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5592\
        );

    \I__964\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5589\
        );

    \I__963\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5584\
        );

    \I__962\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5584\
        );

    \I__961\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5581\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5592\,
            I => \beamYZ0Z_8\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5589\,
            I => \beamYZ0Z_8\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5584\,
            I => \beamYZ0Z_8\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5581\,
            I => \beamYZ0Z_8\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__5572\,
            I => \un4_beamylt8_0_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5561\
        );

    \I__954\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5558\
        );

    \I__953\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5555\
        );

    \I__952\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5550\
        );

    \I__951\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5550\
        );

    \I__950\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5547\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5561\,
            I => \beamYZ0Z_7\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5558\,
            I => \beamYZ0Z_7\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5555\,
            I => \beamYZ0Z_7\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5550\,
            I => \beamYZ0Z_7\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5547\,
            I => \beamYZ0Z_7\
        );

    \I__944\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5529\
        );

    \I__943\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5523\
        );

    \I__942\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5518\
        );

    \I__941\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5518\
        );

    \I__940\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5515\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5529\,
            I => \N__5512\
        );

    \I__938\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5507\
        );

    \I__937\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5507\
        );

    \I__936\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5504\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5523\,
            I => un5_vy
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5518\,
            I => un5_vy
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5515\,
            I => un5_vy
        );

    \I__932\ : Odrv4
    port map (
            O => \N__5512\,
            I => un5_vy
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5507\,
            I => un5_vy
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5504\,
            I => un5_vy
        );

    \I__929\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5483\
        );

    \I__928\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5480\
        );

    \I__927\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5477\
        );

    \I__926\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5472\
        );

    \I__925\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5472\
        );

    \I__924\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5469\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5483\,
            I => \beamYZ0Z_4\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5480\,
            I => \beamYZ0Z_4\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5477\,
            I => \beamYZ0Z_4\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5472\,
            I => \beamYZ0Z_4\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5469\,
            I => \beamYZ0Z_4\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__917\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5452\,
            I => un8_beamylto9_1
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5449\,
            I => \N__5445\
        );

    \I__914\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5438\
        );

    \I__913\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5433\
        );

    \I__912\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5433\
        );

    \I__911\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5430\
        );

    \I__910\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5427\
        );

    \I__909\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5424\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5438\,
            I => \beamYZ0Z_3\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5433\,
            I => \beamYZ0Z_3\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5430\,
            I => \beamYZ0Z_3\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5427\,
            I => \beamYZ0Z_3\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5424\,
            I => \beamYZ0Z_3\
        );

    \I__903\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5410\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \Pixel_RNOZ0Z_5_cascade_\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5404\,
            I => \N_45_cascade_\
        );

    \I__899\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N_76\
        );

    \I__897\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5392\,
            I => \TextOutputEnabledZ0\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \N_74_i_cascade_\
        );

    \I__894\ : IoInMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__892\ : IoSpan4Mux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__891\ : Span4Mux_s2_v
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__5374\,
            I => \Pixel_c\
        );

    \I__889\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__888\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5365\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5358\
        );

    \I__886\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5355\
        );

    \I__885\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5352\
        );

    \I__884\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5347\
        );

    \I__883\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5347\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__5358\,
            I => \beamY_RNI9DLCZ0Z_2\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5355\,
            I => \beamY_RNI9DLCZ0Z_2\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5352\,
            I => \beamY_RNI9DLCZ0Z_2\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5347\,
            I => \beamY_RNI9DLCZ0Z_2\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__5338\,
            I => \N__5332\
        );

    \I__877\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5327\
        );

    \I__876\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5327\
        );

    \I__875\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5324\
        );

    \I__874\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5321\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5327\,
            I => \beamYZ0Z_0\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5324\,
            I => \beamYZ0Z_0\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5321\,
            I => \beamYZ0Z_0\
        );

    \I__870\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5311\,
            I => un5_beamx_5
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__5308\,
            I => \un1_beamy_4_cascade_\
        );

    \I__867\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5302\,
            I => un5_beamx_3
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__864\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5289\
        );

    \I__863\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5284\
        );

    \I__862\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5284\
        );

    \I__861\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5279\
        );

    \I__860\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5279\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5289\,
            I => \beamYZ0Z_1\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5284\,
            I => \beamYZ0Z_1\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5279\,
            I => \beamYZ0Z_1\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__5272\,
            I => \N__5268\
        );

    \I__855\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5265\
        );

    \I__854\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5262\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5265\,
            I => un1_beamy_4
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5262\,
            I => un1_beamy_4
        );

    \I__851\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__850\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5251\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5251\,
            I => un8_beamy_2
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__5248\,
            I => \un1_beamylto9_2_cascade_\
        );

    \I__847\ : IoInMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__845\ : IoSpan4Mux
    port map (
            O => \N__5239\,
            I => \N__5235\
        );

    \I__844\ : IoInMux
    port map (
            O => \N__5238\,
            I => \N__5232\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5226\
        );

    \I__841\ : Span12Mux_v
    port map (
            O => \N__5229\,
            I => \N__5223\
        );

    \I__840\ : Span4Mux_s2_v
    port map (
            O => \N__5226\,
            I => \N__5220\
        );

    \I__839\ : Odrv12
    port map (
            O => \N__5223\,
            I => \VSync_c\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5220\,
            I => \VSync_c\
        );

    \I__837\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5212\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__835\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5203\
        );

    \I__834\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5203\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5203\,
            I => \G_253\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__831\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5194\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5191\,
            I => \N__5186\
        );

    \I__828\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5182\
        );

    \I__827\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5175\
        );

    \I__826\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5175\
        );

    \I__825\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5175\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5182\,
            I => un9_r_0lto2
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5175\,
            I => un9_r_0lto2
        );

    \I__822\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5167\,
            I => \c_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__820\ : InMux
    port map (
            O => \N__5164\,
            I => c_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__819\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__5155\,
            I => un9_r_1lt6_0
        );

    \I__816\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5145\
        );

    \I__815\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5145\
        );

    \I__814\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5142\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5145\,
            I => \N__5139\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5142\,
            I => \N__5136\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__5139\,
            I => \N__5133\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5136\,
            I => c_if_generate_plus_mult1_un68_sum
        );

    \I__809\ : Odrv4
    port map (
            O => \N__5133\,
            I => c_if_generate_plus_mult1_un68_sum
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__807\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5122\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5122\,
            I => \c_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5119\,
            I => \N__5115\
        );

    \I__804\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5111\
        );

    \I__803\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5107\
        );

    \I__802\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5104\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5101\
        );

    \I__800\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5098\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5107\,
            I => un9_r_0lto3
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5104\,
            I => un9_r_0lto3
        );

    \I__797\ : Odrv4
    port map (
            O => \N__5101\,
            I => un9_r_0lto3
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5098\,
            I => un9_r_0lto3
        );

    \I__795\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5083\
        );

    \I__794\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5083\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5083\,
            I => un9_r_0lto3_i
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__791\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N_404_i\
        );

    \I__789\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5065\
        );

    \I__788\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5065\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5065\,
            I => c_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__786\ : InMux
    port map (
            O => \N__5062\,
            I => \bfn_6_10_0_\
        );

    \I__785\ : InMux
    port map (
            O => \N__5059\,
            I => un5_vx_cry_8
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__5056\,
            I => \CO3_0_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__5044\,
            I => \N_14\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__5041\,
            I => \N_3_0_cascade_\
        );

    \I__778\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5035\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__5032\,
            I => c_if_generate_plus_mult1_un75_sum
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__5029\,
            I => \N__5024\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5028\,
            I => \N__5019\
        );

    \I__773\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5016\
        );

    \I__772\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5007\
        );

    \I__771\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5007\
        );

    \I__770\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5007\
        );

    \I__769\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5007\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5016\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5007\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0\
        );

    \I__766\ : InMux
    port map (
            O => \N__5002\,
            I => un5_vx_cry_1
        );

    \I__765\ : InMux
    port map (
            O => \N__4999\,
            I => un5_vx_cry_2
        );

    \I__764\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4990\
        );

    \I__763\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4990\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4990\,
            I => \N__4986\
        );

    \I__761\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4983\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__4986\,
            I => \N__4980\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4983\,
            I => c_if_generate_plus_mult1_un61_sum
        );

    \I__758\ : Odrv4
    port map (
            O => \N__4980\,
            I => c_if_generate_plus_mult1_un61_sum
        );

    \I__757\ : InMux
    port map (
            O => \N__4975\,
            I => un5_vx_cry_3
        );

    \I__756\ : InMux
    port map (
            O => \N__4972\,
            I => un5_vx_cry_4
        );

    \I__755\ : InMux
    port map (
            O => \N__4969\,
            I => un5_vx_cry_5
        );

    \I__754\ : InMux
    port map (
            O => \N__4966\,
            I => un5_vx_cry_6
        );

    \I__753\ : InMux
    port map (
            O => \N__4963\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__4960\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_\
        );

    \I__751\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4951\
        );

    \I__750\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4951\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4951\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11\
        );

    \I__748\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4945\,
            I => \Pixel_RNOZ0Z_7\
        );

    \I__746\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4938\
        );

    \I__745\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4938\,
            I => \N__4930\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4930\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__4927\,
            I => \visibleYZ0Z_3\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__739\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4918\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__736\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4909\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0\
        );

    \I__734\ : InMux
    port map (
            O => \N__4906\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__733\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4900\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4900\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94\
        );

    \I__731\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4894\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0\
        );

    \I__729\ : InMux
    port map (
            O => \N__4891\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4888\,
            I => \N__4884\
        );

    \I__727\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4875\
        );

    \I__726\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4875\
        );

    \I__725\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4875\
        );

    \I__724\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4872\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4875\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4872\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__720\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4861\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4861\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56\
        );

    \I__718\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4855\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4855\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0\
        );

    \I__716\ : InMux
    port map (
            O => \N__4852\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__715\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4846\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4846\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__712\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4837\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__710\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4831\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__708\ : InMux
    port map (
            O => \N__4828\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__707\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4822\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__705\ : InMux
    port map (
            O => \N__4819\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__704\ : InMux
    port map (
            O => \N__4816\,
            I => un21_beamy_cry_8
        );

    \I__703\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4810\,
            I => \N__4807\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__4807\,
            I => if_generate_plus_mult1_un82_sum_s_5
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__4804\,
            I => \N__4801\
        );

    \I__699\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4798\,
            I => un7_r_4
        );

    \I__697\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4791\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__4794\,
            I => \N__4787\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4791\,
            I => \N__4783\
        );

    \I__694\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4780\
        );

    \I__693\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4775\
        );

    \I__692\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4775\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__4783\,
            I => if_generate_plus_mult1_un75_sum_s_5
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4780\,
            I => if_generate_plus_mult1_un75_sum_s_5
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4775\,
            I => if_generate_plus_mult1_un75_sum_s_5
        );

    \I__688\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4765\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__686\ : InMux
    port map (
            O => \N__4762\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__685\ : InMux
    port map (
            O => \N__4759\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__684\ : InMux
    port map (
            O => \N__4756\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__4753\,
            I => \N__4750\
        );

    \I__682\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4747\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__680\ : InMux
    port map (
            O => \N__4744\,
            I => \bfn_6_4_0_\
        );

    \I__679\ : InMux
    port map (
            O => \N__4741\,
            I => un21_beamy_cry_2
        );

    \I__678\ : InMux
    port map (
            O => \N__4738\,
            I => un21_beamy_cry_3
        );

    \I__677\ : InMux
    port map (
            O => \N__4735\,
            I => un21_beamy_cry_4
        );

    \I__676\ : InMux
    port map (
            O => \N__4732\,
            I => un21_beamy_cry_5
        );

    \I__675\ : InMux
    port map (
            O => \N__4729\,
            I => un21_beamy_cry_6
        );

    \I__674\ : InMux
    port map (
            O => \N__4726\,
            I => un21_beamy_cry_7
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__672\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4717\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__670\ : InMux
    port map (
            O => \N__4714\,
            I => c_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__669\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4708\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4708\,
            I => \c_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__667\ : InMux
    port map (
            O => \N__4705\,
            I => c_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__666\ : InMux
    port map (
            O => \N__4702\,
            I => c_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__665\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__664\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4693\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4693\,
            I => \visibleYZ0Z_9\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__661\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4684\,
            I => \visibleY_RNIOR3DZ0Z_9\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__658\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4675\,
            I => \c_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__656\ : InMux
    port map (
            O => \N__4672\,
            I => c_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__655\ : InMux
    port map (
            O => \N__4669\,
            I => c_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__654\ : InMux
    port map (
            O => \N__4666\,
            I => c_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__653\ : InMux
    port map (
            O => \N__4663\,
            I => c_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4660\,
            I => \N__4657\
        );

    \I__651\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4654\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__649\ : InMux
    port map (
            O => \N__4651\,
            I => c_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__648\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4644\
        );

    \I__647\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4641\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4644\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4641\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__643\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4630\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3\
        );

    \I__641\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4624\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__639\ : InMux
    port map (
            O => \N__4621\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__638\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4615\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__636\ : InMux
    port map (
            O => \N__4612\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__4609\,
            I => \N__4605\
        );

    \I__634\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4596\
        );

    \I__633\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4596\
        );

    \I__632\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4596\
        );

    \I__631\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4593\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4596\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4593\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__4588\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__626\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4579\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__624\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4572\
        );

    \I__623\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4572\,
            I => \visibleYZ0Z_8\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4569\,
            I => \visibleYZ0Z_8\
        );

    \I__620\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4561\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0\
        );

    \I__618\ : InMux
    port map (
            O => \N__4558\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__617\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4552\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0\
        );

    \I__615\ : InMux
    port map (
            O => \N__4549\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__614\ : InMux
    port map (
            O => \N__4546\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__613\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4540\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__4537\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__4534\,
            I => \N__4529\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__4533\,
            I => \N__4526\
        );

    \I__608\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4523\
        );

    \I__607\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4520\
        );

    \I__606\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4517\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4523\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4520\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4517\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__602\ : InMux
    port map (
            O => \N__4510\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__601\ : InMux
    port map (
            O => \N__4507\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__4504\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_\
        );

    \I__599\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4495\
        );

    \I__598\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4495\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__4489\,
            I => \visibleYZ0Z_4\
        );

    \I__594\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4482\
        );

    \I__593\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4479\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4482\,
            I => \N__4476\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4479\,
            I => \N__4471\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__4476\,
            I => \N__4471\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__4471\,
            I => \visibleYZ0Z_5\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__587\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4462\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__585\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4456\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1\
        );

    \I__583\ : InMux
    port map (
            O => \N__4453\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__582\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4447\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__579\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4438\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33\
        );

    \I__577\ : InMux
    port map (
            O => \N__4435\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4432\,
            I => \N__4428\
        );

    \I__575\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4419\
        );

    \I__574\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4419\
        );

    \I__573\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4419\
        );

    \I__572\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4416\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4419\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4416\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__568\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4405\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1\
        );

    \I__566\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4399\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3\
        );

    \I__564\ : InMux
    port map (
            O => \N__4396\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__563\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4390\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4390\,
            I => \un5_vy_cry_6_c_RNIG9KKZ0\
        );

    \I__561\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4384\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4384\,
            I => if_generate_plus_mult1_un47_sum_axb_4_l_ofx
        );

    \I__559\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__557\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4365\
        );

    \I__556\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4365\
        );

    \I__555\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4365\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__4372\,
            I => \N__4362\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4365\,
            I => \N__4359\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4362\,
            I => \un5_vy_cry_6_c_RNI9MAAZ0\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__4359\,
            I => \un5_vy_cry_6_c_RNI9MAAZ0\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__4354\,
            I => \N__4351\
        );

    \I__549\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4348\,
            I => \N_7_i\
        );

    \I__547\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4339\
        );

    \I__546\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4336\
        );

    \I__545\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4333\
        );

    \I__544\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4330\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4339\,
            I => if_generate_plus_mult1_un47_sum_s_5
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4336\,
            I => if_generate_plus_mult1_un47_sum_s_5
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4333\,
            I => if_generate_plus_mult1_un47_sum_s_5
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4330\,
            I => if_generate_plus_mult1_un47_sum_s_5
        );

    \I__539\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4318\,
            I => r_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__537\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4307\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__4311\,
            I => \N__4304\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__4310\,
            I => \N__4301\
        );

    \I__533\ : Span4Mux_h
    port map (
            O => \N__4307\,
            I => \N__4296\
        );

    \I__532\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4287\
        );

    \I__531\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4287\
        );

    \I__530\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4287\
        );

    \I__529\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4287\
        );

    \I__528\ : Span4Mux_v
    port map (
            O => \N__4296\,
            I => \N__4282\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4287\,
            I => \N__4282\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__4282\,
            I => \un5_vy_cry_5_c_RNI7J9AZ0\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4279\,
            I => \N__4276\
        );

    \I__524\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4273\,
            I => un5_vy_i_24
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__521\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4264\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__519\ : InMux
    port map (
            O => \N__4261\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__518\ : InMux
    port map (
            O => \N__4258\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__517\ : InMux
    port map (
            O => \N__4255\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__516\ : InMux
    port map (
            O => \N__4252\,
            I => un5_vy_cry_4
        );

    \I__515\ : InMux
    port map (
            O => \N__4249\,
            I => un5_vy_cry_5
        );

    \I__514\ : InMux
    port map (
            O => \N__4246\,
            I => un5_vy_cry_6
        );

    \I__513\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4239\
        );

    \I__512\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4234\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4239\,
            I => \N__4231\
        );

    \I__510\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4228\
        );

    \I__509\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4225\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4234\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4231\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4228\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4225\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__504\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__502\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4204\
        );

    \I__501\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4201\
        );

    \I__500\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4198\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4207\,
            I => if_generate_plus_mult1_un68_sum_s_5
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4204\,
            I => if_generate_plus_mult1_un68_sum_s_5
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4201\,
            I => if_generate_plus_mult1_un68_sum_s_5
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4198\,
            I => if_generate_plus_mult1_un68_sum_s_5
        );

    \I__495\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4182\
        );

    \I__494\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4182\
        );

    \I__493\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4179\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4182\,
            I => \N__4176\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4179\,
            I => r_if_generate_plus_mult1_un54_sum
        );

    \I__490\ : Odrv4
    port map (
            O => \N__4176\,
            I => r_if_generate_plus_mult1_un54_sum
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__488\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4165\,
            I => r_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__486\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4159\,
            I => r_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__484\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4150\
        );

    \I__483\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4147\
        );

    \I__482\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4144\
        );

    \I__481\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4141\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4150\,
            I => if_generate_plus_mult1_un54_sum_s_5_0
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4147\,
            I => if_generate_plus_mult1_un54_sum_s_5_0
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4144\,
            I => if_generate_plus_mult1_un54_sum_s_5_0
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4141\,
            I => if_generate_plus_mult1_un54_sum_s_5_0
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__475\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4126\,
            I => un7_r_1
        );

    \I__473\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4116\
        );

    \I__472\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4116\
        );

    \I__471\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4113\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4113\,
            I => \N__4105\
        );

    \I__468\ : Span4Mux_h
    port map (
            O => \N__4110\,
            I => \N__4105\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__4105\,
            I => r_if_generate_plus_mult1_un47_sum
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__465\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4096\,
            I => r_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__462\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4087\,
            I => r_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__459\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4078\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__457\ : InMux
    port map (
            O => \N__4075\,
            I => r_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__456\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4069\,
            I => r_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__453\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4060\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s_0
        );

    \I__451\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4054\,
            I => \r_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__449\ : InMux
    port map (
            O => \N__4051\,
            I => r_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__448\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4045\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4045\,
            I => \r_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__446\ : InMux
    port map (
            O => \N__4042\,
            I => r_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__445\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4035\
        );

    \I__444\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4032\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4035\,
            I => \N__4028\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4032\,
            I => \N__4025\
        );

    \I__441\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4022\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__4028\,
            I => r_if_generate_plus_mult1_un75_sum
        );

    \I__439\ : Odrv4
    port map (
            O => \N__4025\,
            I => r_if_generate_plus_mult1_un75_sum
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4022\,
            I => r_if_generate_plus_mult1_un75_sum
        );

    \I__437\ : InMux
    port map (
            O => \N__4015\,
            I => un5_vy_cry_0
        );

    \I__436\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4009\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4009\,
            I => \N__4004\
        );

    \I__434\ : InMux
    port map (
            O => \N__4008\,
            I => \N__3999\
        );

    \I__433\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3999\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__4004\,
            I => r_if_generate_plus_mult1_un68_sum
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3999\,
            I => r_if_generate_plus_mult1_un68_sum
        );

    \I__430\ : InMux
    port map (
            O => \N__3994\,
            I => un5_vy_cry_1
        );

    \I__429\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3986\
        );

    \I__428\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3981\
        );

    \I__427\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3981\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3986\,
            I => r_if_generate_plus_mult1_un61_sum
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3981\,
            I => r_if_generate_plus_mult1_un61_sum
        );

    \I__424\ : InMux
    port map (
            O => \N__3976\,
            I => un5_vy_cry_2
        );

    \I__423\ : InMux
    port map (
            O => \N__3973\,
            I => un5_vy_cry_3
        );

    \I__422\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3967\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3967\,
            I => \visibleY_RNINQ3DZ0Z_8\
        );

    \I__420\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3961\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3961\,
            I => \G_251\
        );

    \I__418\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3955\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3955\,
            I => \G_252\
        );

    \I__416\ : InMux
    port map (
            O => \N__3952\,
            I => r_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__415\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3943\
        );

    \I__414\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3943\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3943\,
            I => \G_250\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__3940\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_\
        );

    \I__411\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3933\
        );

    \I__410\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3930\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3933\,
            I => \N__3927\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3930\,
            I => \visibleYZ0Z_7\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__3927\,
            I => \visibleYZ0Z_7\
        );

    \I__406\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3919\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3919\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0\
        );

    \I__404\ : InMux
    port map (
            O => \N__3916\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__3913\,
            I => \N__3910\
        );

    \I__402\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3907\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3907\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01\
        );

    \I__400\ : InMux
    port map (
            O => \N__3904\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__399\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3898\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01\
        );

    \I__397\ : InMux
    port map (
            O => \N__3895\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__396\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3889\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3889\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__394\ : InMux
    port map (
            O => \N__3886\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__393\ : InMux
    port map (
            O => \N__3883\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__3880\,
            I => \N__3875\
        );

    \I__391\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3865\
        );

    \I__390\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3865\
        );

    \I__389\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3865\
        );

    \I__388\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3865\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3865\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3862\,
            I => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3859\,
            I => \N__3856\
        );

    \I__384\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3853\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3853\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__382\ : InMux
    port map (
            O => \N__3850\,
            I => r_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__381\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3843\
        );

    \I__380\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3840\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3843\,
            I => \N__3835\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3835\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__3835\,
            I => \visibleYZ0Z_6\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__3832\,
            I => \N__3829\
        );

    \I__375\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3826\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3826\,
            I => \N__3823\
        );

    \I__373\ : Odrv4
    port map (
            O => \N__3823\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__372\ : InMux
    port map (
            O => \N__3820\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__371\ : InMux
    port map (
            O => \N__3817\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__370\ : InMux
    port map (
            O => \N__3814\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__369\ : InMux
    port map (
            O => \N__3811\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__368\ : InMux
    port map (
            O => \N__3808\,
            I => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__367\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__3802\,
            I => \N__3799\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__3799\,
            I => \r_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__364\ : InMux
    port map (
            O => \N__3796\,
            I => r_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__363\ : InMux
    port map (
            O => \N__3793\,
            I => r_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__361\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3784\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3784\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s_0
        );

    \I__359\ : InMux
    port map (
            O => \N__3781\,
            I => r_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__358\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3775\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3775\,
            I => \r_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__356\ : InMux
    port map (
            O => \N__3772\,
            I => r_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__355\ : InMux
    port map (
            O => \N__3769\,
            I => r_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__3766\,
            I => \N__3763\
        );

    \I__353\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3760\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3760\,
            I => if_generate_plus_mult1_un47_sum_cry_3_s
        );

    \I__351\ : InMux
    port map (
            O => \N__3757\,
            I => r_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__350\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3751\,
            I => \r_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__348\ : InMux
    port map (
            O => \N__3748\,
            I => r_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__347\ : InMux
    port map (
            O => \N__3745\,
            I => r_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__346\ : InMux
    port map (
            O => \N__3742\,
            I => r_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__345\ : InMux
    port map (
            O => \N__3739\,
            I => r_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__344\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3733\,
            I => r_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__341\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3724\,
            I => r_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__338\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__336\ : Odrv4
    port map (
            O => \N__3712\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s_0
        );

    \I__335\ : InMux
    port map (
            O => \N__3709\,
            I => r_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__334\ : IoInMux
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__332\ : Span4Mux_s1_h
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__331\ : Span4Mux_h
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__3694\,
            I => \N__3691\
        );

    \I__329\ : Odrv4
    port map (
            O => \N__3691\,
            I => \Clock50MHz.PixelClock\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__3688\,
            I => \N__3685\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3685\,
            I => \N__3682\
        );

    \I__326\ : IoSpan4Mux
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__3679\,
            I => \Clock12MHz_c\
        );

    \INVPixelZ0C\ : INV
    port map (
            O => \INVPixelZ0C_net\,
            I => \N__7367\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_vx_cry_7,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un21_beamy_cry_1_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3706\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \beamX_RNISO4T_0_7\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5695\,
            GLOBALBUFFEROUTPUT => un15_beamy_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \visibleY_4_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4007\,
            in2 => \_gnd_net_\,
            in3 => \N__4008\,
            lcout => \visibleYZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => r_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \N__7363\,
            ce => \N__7295\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un68_sum_cry_3_s_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4243\,
            in2 => \N__3730\,
            in3 => \N__3745\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s_0,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un75_sum_axb_5_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4211\,
            in1 => \N__3736\,
            in2 => \N__3721\,
            in3 => \N__3742\,
            lcout => \r_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un68_sum_s_5_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3805\,
            in2 => \_gnd_net_\,
            in3 => \N__3739\,
            lcout => if_generate_plus_mult1_un68_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4237\,
            lcout => r_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3991\,
            lcout => r_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un68_sum_sbtinv_5_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4210\,
            lcout => r_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_5_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3989\,
            in2 => \_gnd_net_\,
            in3 => \N__3990\,
            lcout => \visibleYZ0Z_5\,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => r_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \N__7357\,
            ce => \N__7292\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4155\,
            in2 => \N__4171\,
            in3 => \N__3709\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s_0,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un68_sum_axb_5_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4238\,
            in1 => \N__4162\,
            in2 => \N__3790\,
            in3 => \N__3796\,
            lcout => \r_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un61_sum_s_5_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3778\,
            in2 => \_gnd_net_\,
            in3 => \N__3793\,
            lcout => if_generate_plus_mult1_un61_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_6_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4188\,
            in2 => \_gnd_net_\,
            in3 => \N__4189\,
            lcout => \visibleYZ0Z_6\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => r_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \N__7354\,
            ce => \N__7289\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4344\,
            in2 => \N__4102\,
            in3 => \N__3781\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s_0,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un61_sum_axb_5_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4154\,
            in1 => \N__4321\,
            in2 => \N__3766\,
            in3 => \N__3772\,
            lcout => \r_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un54_sum_s_5_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3754\,
            in2 => \_gnd_net_\,
            in3 => \N__3769\,
            lcout => if_generate_plus_mult1_un54_sum_s_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_7_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4122\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => \visibleYZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => r_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \N__7353\,
            ce => \N__7288\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4393\,
            in2 => \N__4279\,
            in3 => \N__3757\,
            lcout => if_generate_plus_mult1_un47_sum_cry_3_s,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un54_sum_axb_5_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4343\,
            in1 => \N__4387\,
            in2 => \N__4354\,
            in3 => \N__3748\,
            lcout => \r_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un47_sum_s_5_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3850\,
            lcout => if_generate_plus_mult1_un47_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3936\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3847\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3846\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71E1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3874\,
            in2 => \N__3832\,
            in3 => \N__3820\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5T1_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3922\,
            in2 => \N__3880\,
            in3 => \N__3817\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4T32_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3878\,
            in2 => \N__3913\,
            in3 => \N__3814\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQP8K3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4426\,
            in1 => \N__3901\,
            in2 => \N__3859\,
            in3 => \N__3811\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8G1_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3892\,
            in1 => \N__3879\,
            in2 => \N__4534\,
            in3 => \N__3808\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5K3_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__4648\,
            in1 => \_gnd_net_\,
            in2 => \N__3940\,
            in3 => \_gnd_net_\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3937\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450Q_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3970\,
            in2 => \N__7779\,
            in3 => \N__3916\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9M01_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4564\,
            in2 => \N__7781\,
            in3 => \N__3904\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDO01_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4555\,
            in2 => \N__7780\,
            in3 => \N__3895\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4533\,
            in3 => \N__3886\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4543\,
            in2 => \_gnd_net_\,
            in3 => \N__3883\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3862\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_RNINQ3D_8_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4576\,
            lcout => \visibleY_RNINQ3DZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_8_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4315\,
            lcout => \visibleYZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7356\,
            ce => \N__7287\,
            sr => \_gnd_net_\
        );

    \visibleY_9_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4381\,
            lcout => \visibleYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7356\,
            ce => \N__7287\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3948\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => r_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_cry_3_c_inv_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3964\,
            in2 => \N__4794\,
            in3 => \N__4038\,
            lcout => \G_251\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3958\,
            in2 => \N__4084\,
            in3 => \N__4786\,
            lcout => \G_252\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_s_5_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4057\,
            in2 => \_gnd_net_\,
            in3 => \N__3952\,
            lcout => if_generate_plus_mult1_un82_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__7706\,
            in1 => \N__3949\,
            in2 => \_gnd_net_\,
            in3 => \N__5536\,
            lcout => \G_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un68_sum_sbtinv_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4012\,
            lcout => r_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_3_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4031\,
            in2 => \_gnd_net_\,
            in3 => \N__4039\,
            lcout => \visibleYZ0Z_3\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => r_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \N__7369\,
            ce => \N__7299\,
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4212\,
            in2 => \N__4093\,
            in3 => \N__4075\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => r_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un82_sum_axb_5_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4790\,
            in1 => \N__4072\,
            in2 => \N__4066\,
            in3 => \N__4051\,
            lcout => \r_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => r_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => r_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un75_sum_s_5_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4048\,
            in2 => \_gnd_net_\,
            in3 => \N__4042\,
            lcout => if_generate_plus_mult1_un75_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_0_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => un5_vy_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_0_c_RNIT34A_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5441\,
            in2 => \_gnd_net_\,
            in3 => \N__4015\,
            lcout => r_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_vy_cry_0,
            carryout => un5_vy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_1_c_RNIV65A_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5486\,
            in2 => \_gnd_net_\,
            in3 => \N__3994\,
            lcout => r_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_vy_cry_1,
            carryout => un5_vy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_2_c_RNI1A6A_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5653\,
            in2 => \N__7702\,
            in3 => \N__3976\,
            lcout => r_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_vy_cry_2,
            carryout => un5_vy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_3_c_RNI3D7A_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5677\,
            in2 => \N__7704\,
            in3 => \N__3973\,
            lcout => r_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_vy_cry_3,
            carryout => un5_vy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_4_c_RNI5G8A_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5564\,
            in2 => \N__7703\,
            in3 => \N__4252\,
            lcout => r_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_vy_cry_4,
            carryout => un5_vy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_5_c_RNI7J9A_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5595\,
            in2 => \N__7705\,
            in3 => \N__4249\,
            lcout => \un5_vy_cry_5_c_RNI7J9AZ0\,
            ltout => OPEN,
            carryin => un5_vy_cry_5,
            carryout => un5_vy_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_6_c_RNI9MAA_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5622\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \un5_vy_cry_6_c_RNI9MAAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TextOutputEnabled_RNO_0_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6085\,
            in1 => \N__4242\,
            in2 => \N__4132\,
            in3 => \N__4216\,
            lcout => un7_r_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4187\,
            lcout => r_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4153\,
            lcout => r_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TextOutputEnabled_RNO_2_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5053\,
            in1 => \N__4156\,
            in2 => \_gnd_net_\,
            in3 => \N__4345\,
            lcout => un7_r_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un47_sum_sbtinv_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4121\,
            lcout => r_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4485\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_6_c_RNIG9KK_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4300\,
            in2 => \_gnd_net_\,
            in3 => \N__4375\,
            lcout => \un5_vy_cry_6_c_RNIG9KKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un47_sum_axb_4_l_ofx_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4376\,
            in1 => \_gnd_net_\,
            in2 => \N__4310\,
            in3 => \_gnd_net_\,
            lcout => if_generate_plus_mult1_un47_sum_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_6_c_RNIG9KK_0_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__4377\,
            in1 => \_gnd_net_\,
            in2 => \N__4311\,
            in3 => \_gnd_net_\,
            lcout => \N_7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_if_generate_plus_mult1_un47_sum_sbtinv_5_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4342\,
            lcout => r_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vy_cry_5_c_RNI7J9A_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4299\,
            lcout => un5_vy_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4500\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73P94_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4604\,
            in2 => \N__4270\,
            in3 => \N__4261\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQ56_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4459\,
            in2 => \N__4609\,
            in3 => \N__4258\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUT97_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4608\,
            in2 => \N__4444\,
            in3 => \N__4255\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIP00TH_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4882\,
            in1 => \N__4402\,
            in2 => \N__4585\,
            in3 => \N__4510\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4627\,
            in2 => \_gnd_net_\,
            in3 => \N__4507\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4504\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4501\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSV1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4427\,
            in2 => \N__4468\,
            in3 => \N__4453\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0V33_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4450\,
            in2 => \N__4432\,
            in3 => \N__4435\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4J3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4431\,
            in2 => \N__4411\,
            in3 => \N__4396\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI9FRN9_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4603\,
            in1 => \N__4647\,
            in2 => \N__4636\,
            in3 => \N__4621\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4618\,
            in2 => \_gnd_net_\,
            in3 => \N__4612\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_0_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4588\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4575\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJ_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7753\,
            in2 => \N__4690\,
            in3 => \N__4558\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJ_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4699\,
            in2 => \N__7778\,
            in3 => \N__4549\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4546\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4537\,
            in3 => \N__4532\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_RNIOR3D_9_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4698\,
            lcout => \visibleY_RNIOR3DZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un61_sum_i_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4989\,
            lcout => \c_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5151\,
            in2 => \_gnd_net_\,
            in3 => \N__5152\,
            lcout => \N_84\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => c_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \N__7359\,
            ce => \N__7290\,
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un68_sum_cry_2_s_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5088\,
            in2 => \N__4681\,
            in3 => \N__4672\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => c_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5114\,
            in2 => \N__4660\,
            in3 => \N__4669\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => c_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un75_sum_axb_5_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5190\,
            in1 => \N__5089\,
            in2 => \N__4723\,
            in3 => \N__4666\,
            lcout => \c_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => c_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un68_sum_s_5_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4711\,
            in2 => \_gnd_net_\,
            in3 => \N__4663\,
            lcout => un9_r_0lto2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_4_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4995\,
            in2 => \_gnd_net_\,
            in3 => \N__4996\,
            lcout => \visibleXZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => c_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \N__7364\,
            ce => \N__7293\,
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5070\,
            in2 => \N__5080\,
            in3 => \N__4651\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => c_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6078\,
            in2 => \N__6196\,
            in3 => \N__4714\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => c_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un68_sum_axb_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5118\,
            in1 => \N__5071\,
            in2 => \N__6157\,
            in3 => \N__4705\,
            lcout => \c_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => c_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un61_sum_s_5_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6106\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => un9_r_0lto3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleY_1_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5292\,
            in2 => \N__5338\,
            in3 => \N__5293\,
            lcout => \visibleYZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => un21_beamy_cry_1,
            clk => \N__7371\,
            ce => \N__7300\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7723\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => \un21_beamy_cry_1_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__7766\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_0_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_2_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7727\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_1_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_3_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__7767\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_2_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_4_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7731\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_3_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_5_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__7768\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_4_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_THRU_CRY_6_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7735\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un21_beamy_cry_1_THRU_CRY_5_THRU_CO\,
            carryout => \un21_beamy_cry_1_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5532\,
            in2 => \_gnd_net_\,
            in3 => \N__4744\,
            lcout => un5_vy,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => un21_beamy_cry_2,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5370\,
            in1 => \N__5448\,
            in2 => \_gnd_net_\,
            in3 => \N__4741\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5361\,
            in1 => \N__5490\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5656\,
            in2 => \_gnd_net_\,
            in3 => \N__4735\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5680\,
            in2 => \_gnd_net_\,
            in3 => \N__4732\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5371\,
            in1 => \N__5568\,
            in2 => \_gnd_net_\,
            in3 => \N__4729\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5599\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__5628\,
            in1 => \N__5362\,
            in2 => \_gnd_net_\,
            in3 => \N__4816\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7370\,
            ce => \N__6250\,
            sr => \_gnd_net_\
        );

    \visibleY_2_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5535\,
            lcout => \visibleYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7365\,
            ce => \N__7296\,
            sr => \_gnd_net_\
        );

    \TextOutputEnabled_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5161\,
            in1 => \N__4813\,
            in2 => \N__4804\,
            in3 => \N__4795\,
            lcout => \TextOutputEnabledZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7365\,
            ce => \N__7296\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5807\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSI_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4768\,
            in2 => \N__5028\,
            in3 => \N__4762\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GT_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5022\,
            in2 => \N__4915\,
            in3 => \N__4759\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7C11_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4897\,
            in2 => \N__5029\,
            in3 => \N__4756\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4858\,
            in2 => \N__4753\,
            in3 => \N__5023\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGC41_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4834\,
            in2 => \_gnd_net_\,
            in3 => \N__4963\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41\,
            ltout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_3_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__4957\,
            in1 => \_gnd_net_\,
            in2 => \N__4960\,
            in3 => \N__4948\,
            lcout => \N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_7_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000010"
        )
    port map (
            in0 => \N__5808\,
            in1 => \N__5842\,
            in2 => \N__5782\,
            in3 => \N__4956\,
            lcout => \Pixel_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4941\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000B_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4883\,
            in2 => \N__4924\,
            in3 => \N__4906\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SE_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4903\,
            in2 => \N__4888\,
            in3 => \N__4891\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OG_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4887\,
            in2 => \N__4867\,
            in3 => \N__4852\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI2VO741_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5027\,
            in1 => \N__4849\,
            in2 => \N__4843\,
            in3 => \N__4828\,
            lcout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBI_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__4819\,
            lcout => \chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__6344\,
            in1 => \N__6314\,
            in2 => \N__6649\,
            in3 => \N__6283\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_0_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6281\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => un5_vx_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6282\,
            in1 => \N__6313\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => un5_vx_cry_0,
            carryout => un5_vx_cry_1,
            clk => \N__7358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_1_c_RNIRP5_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6343\,
            in2 => \_gnd_net_\,
            in3 => \N__5002\,
            lcout => c_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_vx_cry_1,
            carryout => un5_vx_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_2_c_RNITS6_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6642\,
            in2 => \N__7782\,
            in3 => \N__4999\,
            lcout => c_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_vx_cry_2,
            carryout => un5_vx_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_3_c_RNIVV7_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6710\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => c_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_vx_cry_3,
            carryout => un5_vx_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_4_c_RNI139_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6674\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => c_if_generate_plus_mult1_un47_sum1_0,
            ltout => OPEN,
            carryin => un5_vx_cry_4,
            carryout => un5_vx_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_5_c_RNI36A_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7774\,
            in2 => \N__6748\,
            in3 => \N__4969\,
            lcout => c_if_generate_plus_mult1_un47_sum_1,
            ltout => OPEN,
            carryin => un5_vx_cry_5,
            carryout => un5_vx_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_6_c_RNI59B_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7135\,
            in2 => \_gnd_net_\,
            in3 => \N__4966\,
            lcout => \un5_vx_cry_6_c_RNI59BZ0\,
            ltout => OPEN,
            carryin => un5_vx_cry_6,
            carryout => un5_vx_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_7_c_RNI7CC_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5899\,
            in2 => \N__7783\,
            in3 => \N__5062\,
            lcout => c_if_generate_plus_mult1_un47_sum_0_0,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => un5_vx_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_8_c_RNI9FD_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5861\,
            in2 => \_gnd_net_\,
            in3 => \N__5059\,
            lcout => \CO3_0\,
            ltout => \CO3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TextOutputEnabled_RNO_3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__5988\,
            in1 => \N__6807\,
            in2 => \N__5056\,
            in3 => \N__6508\,
            lcout => \N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_7_c_RNIL451_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__7439\,
            in1 => \N__6476\,
            in2 => \_gnd_net_\,
            in3 => \N__6027\,
            lcout => \N_13_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_6_c_RNI59B_1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_vx_i_0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_7_c_RNICLN_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6474\,
            in2 => \_gnd_net_\,
            in3 => \N__6026\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__6028\,
            in1 => \N__7440\,
            in2 => \N__5041\,
            in3 => \N__6479\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_axb_5_sbtinv_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7435\,
            lcout => c_if_generate_plus_mult1_un47_sum_0_axb_5_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5038\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => c_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5208\,
            in2 => \N__5128\,
            in3 => \N__5185\,
            lcout => \G_253\,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => c_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un75_sum_cry_3_c_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5215\,
            in2 => \N__5191\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => c_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5209\,
            in2 => \N__5200\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => c_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TextOutputEnabled_RNO_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000111"
        )
    port map (
            in0 => \N__5189\,
            in1 => \N__5170\,
            in2 => \N__5119\,
            in3 => \N__5164\,
            lcout => un9_r_1lt6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un68_sum_i_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5150\,
            lcout => \c_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un9_r_0lto3_sbtinv_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5110\,
            lcout => un9_r_0lto3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_N_404_i_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5971\,
            lcout => \N_404_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6070\,
            lcout => c_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__5336\,
            in1 => \N__5363\,
            in2 => \_gnd_net_\,
            in3 => \N__6249\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001001110000"
        )
    port map (
            in0 => \N__6248\,
            in1 => \N__5364\,
            in2 => \N__5299\,
            in3 => \N__5337\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5305\,
            in1 => \N__5533\,
            in2 => \N__5272\,
            in3 => \N__5314\,
            lcout => \beamY_RNI9DLCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC725_0_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__5335\,
            in2 => \N__5629\,
            in3 => \N__5444\,
            lcout => un5_beamx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4H2_5_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5678\,
            in2 => \_gnd_net_\,
            in3 => \N__5654\,
            lcout => un1_beamy_4,
            ltout => \un1_beamy_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIH3B6_7_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5256\,
            in2 => \N__5308\,
            in3 => \N__5565\,
            lcout => un8_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITAH2_9_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5623\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => un8_beamy_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEIP3_1_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5489\,
            in1 => \N__5566\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => un5_beamx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_RNO_0_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__5295\,
            in1 => \N__5569\,
            in2 => \N__5449\,
            in3 => \N__5534\,
            lcout => OPEN,
            ltout => \un1_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__5271\,
            in1 => \N__5257\,
            in2 => \N__5248\,
            in3 => \N__5491\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5442\,
            in2 => \_gnd_net_\,
            in3 => \N__5527\,
            lcout => OPEN,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_5_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5679\,
            in1 => \N__5655\,
            in2 => \N__5632\,
            in3 => \N__5487\,
            lcout => OPEN,
            ltout => \un4_beamylt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_9_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__5627\,
            in1 => \N__5598\,
            in2 => \N__5572\,
            in3 => \N__5567\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5528\,
            in1 => \N__5488\,
            in2 => \N__5458\,
            in3 => \N__5443\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__5806\,
            in1 => \N__5840\,
            in2 => \N__5827\,
            in3 => \N__5781\,
            lcout => OPEN,
            ltout => \Pixel_RNOZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5413\,
            in2 => \N__5407\,
            in3 => \N__5761\,
            lcout => OPEN,
            ltout => \N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010110100"
        )
    port map (
            in0 => \N__6361\,
            in1 => \N__6415\,
            in2 => \N__5404\,
            in3 => \N__5401\,
            lcout => OPEN,
            ltout => \N_74_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__7546\,
            in1 => \N__5395\,
            in2 => \N__5389\,
            in3 => \N__5752\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVPixelZ0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_6_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__5823\,
            in2 => \N__5809\,
            in3 => \N__5780\,
            lcout => \Pixel_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI8P51_4_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__6712\,
            in1 => \N__6743\,
            in2 => \N__6684\,
            in3 => \N__5746\,
            lcout => un13_beamylt7,
            ltout => \un13_beamylt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \OutputEnabled_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__7138\,
            in1 => \N__7166\,
            in2 => \N__5755\,
            in3 => \N__5710\,
            lcout => \OutputEnabledZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5871\,
            in2 => \_gnd_net_\,
            in3 => \N__5897\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNII5M_9_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5896\,
            in1 => \N__7136\,
            in2 => \N__5872\,
            in3 => \N__6744\,
            lcout => OPEN,
            ltout => \un18_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_4_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__5745\,
            in1 => \N__6678\,
            in2 => \N__5734\,
            in3 => \N__6711\,
            lcout => OPEN,
            ltout => \un18_beamylt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIT9ER_10_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__7205\,
            in2 => \N__5722\,
            in3 => \N__5719\,
            lcout => un15_beamy_2,
            ltout => \un15_beamy_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNISO4T_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110000"
        )
    port map (
            in0 => \N__7137\,
            in1 => \N__5704\,
            in2 => \N__5698\,
            in3 => \N__7165\,
            lcout => \beamX_RNISO4TZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6318\,
            in2 => \N__6289\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6346\,
            in2 => \_gnd_net_\,
            in3 => \N__5917\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6648\,
            in2 => \_gnd_net_\,
            in3 => \N__5914\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6239\,
            in1 => \N__6715\,
            in2 => \_gnd_net_\,
            in3 => \N__5911\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6683\,
            in2 => \_gnd_net_\,
            in3 => \N__5908\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6747\,
            in2 => \_gnd_net_\,
            in3 => \N__5905\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7140\,
            in2 => \_gnd_net_\,
            in3 => \N__5902\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5898\,
            in2 => \_gnd_net_\,
            in3 => \N__5875\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__7355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5867\,
            in2 => \_gnd_net_\,
            in3 => \N__5845\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6234\,
            in1 => \N__7204\,
            in2 => \_gnd_net_\,
            in3 => \N__5953\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6235\,
            in2 => \_gnd_net_\,
            in3 => \N__6288\,
            lcout => un5_vx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_6_c_RNI59B_0_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6477\,
            lcout => un5_vx_i_25,
            ltout => \un5_vx_i_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__7438\,
            in1 => \N__6803\,
            in2 => \N__5950\,
            in3 => \N__6029\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7436\,
            lcout => if_generate_plus_mult1_un47_sum_0_cry_3_ma,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__6478\,
            in1 => \N__7434\,
            in2 => \_gnd_net_\,
            in3 => \N__6800\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_vx_cry_8_c_RNIL451_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7437\,
            lcout => \N_186_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6610\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => c_if_generate_plus_mult1_un47_sum_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_m_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__6574\,
            in1 => \N__7449\,
            in2 => \N__5947\,
            in3 => \N__5938\,
            lcout => if_generate_plus_mult1_un47_sum_m_2,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_1_cry_1,
            carryout => c_if_generate_plus_mult1_un47_sum_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5935\,
            in2 => \N__5929\,
            in3 => \N__5920\,
            lcout => c_if_generate_plus_mult1_un47_sum1_3,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_1_cry_2,
            carryout => c_if_generate_plus_mult1_un47_sum_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6046\,
            in2 => \N__7466\,
            in3 => \N__6040\,
            lcout => c_if_generate_plus_mult1_un47_sum1_4,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_1_cry_3,
            carryout => c_if_generate_plus_mult1_un47_sum_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__7450\,
            in1 => \N__6480\,
            in2 => \N__6034\,
            in3 => \N__6037\,
            lcout => c_if_generate_plus_mult1_un47_sum1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_8_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6033\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \visibleXZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7366\,
            ce => \N__7294\,
            sr => \_gnd_net_\
        );

    \un5_vx_cry_8_c_RNI24IE_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__7454\,
            in1 => \N__5984\,
            in2 => \_gnd_net_\,
            in3 => \N__6503\,
            lcout => \N_18\,
            ltout => \N_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_axb_5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__6523\,
            in2 => \N__5998\,
            in3 => \N__7458\,
            lcout => \c_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__7455\,
            in1 => \N__6618\,
            in2 => \N__6141\,
            in3 => \N__6619\,
            lcout => if_generate_plus_mult1_un54_sum_axb_2_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5995\,
            in1 => \N__7457\,
            in2 => \N__6142\,
            in3 => \N__6544\,
            lcout => if_generate_plus_mult1_un54_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__6504\,
            in1 => \N__6171\,
            in2 => \N__5989\,
            in3 => \N__7456\,
            lcout => if_generate_plus_mult1_un54_sum_axb_3_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_5_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5969\,
            in2 => \_gnd_net_\,
            in3 => \N__5970\,
            lcout => \visibleXZ0Z_5\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => c_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \N__7372\,
            ce => \N__7297\,
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6133\,
            in2 => \N__6205\,
            in3 => \N__6184\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => c_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6181\,
            in2 => \N__6175\,
            in3 => \N__6145\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => c_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6071\,
            in1 => \N__6134\,
            in2 => \N__6115\,
            in3 => \N__6097\,
            lcout => \c_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => c_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6094\,
            in2 => \_gnd_net_\,
            in3 => \N__6088\,
            lcout => if_generate_plus_mult1_un54_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6386\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HC_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6441\,
            in2 => \N__6355\,
            in3 => \N__6052\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_8_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6886\,
            in2 => \N__6850\,
            in3 => \N__6049\,
            lcout => \Pixel_RNOZ0Z_8\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6442\,
            in2 => \N__6874\,
            in3 => \N__6845\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53L_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6862\,
            in2 => \_gnd_net_\,
            in3 => \N__6433\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0\,
            ltout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001010111111"
        )
    port map (
            in0 => \N__6387\,
            in1 => \N__6430\,
            in2 => \N__6418\,
            in3 => \N__6408\,
            lcout => \N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_4_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__6409\,
            in1 => \N__6397\,
            in2 => \N__6391\,
            in3 => \N__6367\,
            lcout => \N_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_RNIJK0C_5_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6904\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6713\,
            in1 => \N__6345\,
            in2 => \N__7206\,
            in3 => \N__6322\,
            lcout => OPEN,
            ltout => \un3_beamx_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6745\,
            in1 => \N__6646\,
            in2 => \N__6292\,
            in3 => \N__6284\,
            lcout => OPEN,
            ltout => \un3_beamx_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7167\,
            in1 => \N__7139\,
            in2 => \N__6253\,
            in3 => \N__6679\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_RNO_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6746\,
            in1 => \N__6714\,
            in2 => \N__6685\,
            in3 => \N__6647\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_6_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6616\,
            in2 => \_gnd_net_\,
            in3 => \N__6617\,
            lcout => \visibleXZ0Z_6\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => c_if_generate_plus_mult1_un47_sum_0_cry_1,
            clk => \N__7368\,
            ce => \N__7291\,
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6589\,
            in2 => \N__6583\,
            in3 => \N__6562\,
            lcout => c_if_generate_plus_mult1_un47_sum0_2,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_0_cry_1,
            carryout => c_if_generate_plus_mult1_un47_sum_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6559\,
            in2 => \N__6553\,
            in3 => \N__6535\,
            lcout => c_if_generate_plus_mult1_un47_sum0_3,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_0_cry_2,
            carryout => c_if_generate_plus_mult1_un47_sum_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6778\,
            in2 => \N__6532\,
            in3 => \N__6514\,
            lcout => c_if_generate_plus_mult1_un47_sum0_4,
            ltout => OPEN,
            carryin => c_if_generate_plus_mult1_un47_sum_0_cry_3,
            carryout => c_if_generate_plus_mult1_un47_sum_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7467\,
            in2 => \_gnd_net_\,
            in3 => \N__6511\,
            lcout => c_if_generate_plus_mult1_un47_sum0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6484\,
            lcout => \visibleXZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7368\,
            ce => \N__7291\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7488\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BD1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6912\,
            in2 => \N__6817\,
            in3 => \N__6832\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMK642_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6928\,
            in2 => \N__6760\,
            in3 => \N__6829\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3O524_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__6913\,
            in2 => \N__6952\,
            in3 => \N__6826\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__6823\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412\,
            ltout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6820\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_RNIMN0C_8_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__7459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6808\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6771\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29R21_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7566\,
            in2 => \N__7792\,
            in3 => \N__6751\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKV_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7578\,
            in2 => \N__7252\,
            in3 => \N__6943\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIS2GV1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6927\,
            in1 => \N__7567\,
            in2 => \N__7240\,
            in3 => \N__6934\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__7228\,
            in1 => \N__7579\,
            in2 => \_gnd_net_\,
            in3 => \N__6931\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6926\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6903\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56B05_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7495\,
            in2 => \N__7072\,
            in3 => \N__6877\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIC7997_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7051\,
            in2 => \N__6970\,
            in3 => \N__6865\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI25I2L_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6849\,
            in1 => \N__7216\,
            in2 => \N__7021\,
            in3 => \N__6856\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJ19_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6988\,
            in2 => \_gnd_net_\,
            in3 => \N__6853\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEA08_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__7020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6965\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__7210\,
            in1 => \N__7174\,
            in2 => \N__7147\,
            in3 => \N__7105\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_RNIKL0C_6_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7063\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7062\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTK2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7005\,
            in2 => \N__7477\,
            in3 => \N__7045\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19M3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7042\,
            in2 => \N__7030\,
            in3 => \N__7009\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNI547N8_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6969\,
            in1 => \N__7006\,
            in2 => \N__6997\,
            in3 => \N__6982\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6979\,
            in2 => \_gnd_net_\,
            in3 => \N__6973\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4\,
            ltout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7498\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_RNILM0C_7_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7489\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_9_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7468\,
            lcout => \visibleXZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7374\,
            ce => \N__7298\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7800\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8P8_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7736\,
            in2 => \_gnd_net_\,
            in3 => \N__7243\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQ8_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7740\,
            in2 => \N__7769\,
            in3 => \N__7231\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7222\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7219\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \visibleX_RNINO0C_9_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7770\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7591\,
            in3 => \N__7582\,
            lcout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0\,
            ltout => \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7570\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \N_75_i_i_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__7555\,
            in1 => \N__7509\,
            in2 => \_gnd_net_\,
            in3 => \N__7521\,
            lcout => \G_256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \N_555_i_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7520\,
            lcout => \G_255\,
            ltout => \G_255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CharacterDisplay.Z_decfrac15_0_a2_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__7508\,
            in1 => \_gnd_net_\,
            in2 => \N__7558\,
            in3 => \N__7554\,
            lcout => \CharacterDisplay__decfrac8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SUM1_3_0_x2_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7510\,
            in2 => \_gnd_net_\,
            in3 => \N__7522\,
            lcout => \G_254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
