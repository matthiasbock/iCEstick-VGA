// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 17:51:28

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__4782;
    wire N__4781;
    wire N__4780;
    wire N__4773;
    wire N__4772;
    wire N__4771;
    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4746;
    wire N__4745;
    wire N__4744;
    wire N__4737;
    wire N__4736;
    wire N__4735;
    wire N__4728;
    wire N__4727;
    wire N__4726;
    wire N__4709;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4645;
    wire N__4644;
    wire N__4643;
    wire N__4636;
    wire N__4633;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4576;
    wire N__4573;
    wire N__4572;
    wire N__4571;
    wire N__4564;
    wire N__4561;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4540;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4453;
    wire N__4450;
    wire N__4441;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4347;
    wire N__4340;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4273;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4258;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4184;
    wire N__4183;
    wire N__4182;
    wire N__4181;
    wire N__4180;
    wire N__4179;
    wire N__4178;
    wire N__4177;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4150;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4032;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4020;
    wire N__4017;
    wire N__4012;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4002;
    wire N__4001;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3986;
    wire N__3979;
    wire N__3972;
    wire N__3971;
    wire N__3970;
    wire N__3969;
    wire N__3966;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3946;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3883;
    wire N__3882;
    wire N__3877;
    wire N__3874;
    wire N__3873;
    wire N__3872;
    wire N__3867;
    wire N__3862;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3784;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3776;
    wire N__3773;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3757;
    wire N__3754;
    wire N__3753;
    wire N__3752;
    wire N__3745;
    wire N__3742;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3724;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3706;
    wire N__3705;
    wire N__3700;
    wire N__3697;
    wire N__3692;
    wire N__3689;
    wire N__3688;
    wire N__3687;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3616;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3586;
    wire N__3585;
    wire N__3578;
    wire N__3575;
    wire N__3574;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3544;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3536;
    wire N__3533;
    wire N__3528;
    wire N__3525;
    wire N__3524;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3514;
    wire N__3509;
    wire N__3504;
    wire N__3497;
    wire N__3496;
    wire N__3495;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3489;
    wire N__3486;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3461;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3455;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3428;
    wire N__3427;
    wire N__3424;
    wire N__3423;
    wire N__3422;
    wire N__3421;
    wire N__3418;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3398;
    wire N__3397;
    wire N__3394;
    wire N__3393;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3378;
    wire N__3371;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3346;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3295;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3256;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3244;
    wire N__3239;
    wire N__3238;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3202;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3142;
    wire N__3141;
    wire N__3134;
    wire N__3133;
    wire N__3132;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3101;
    wire N__3098;
    wire N__3097;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3089;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3065;
    wire N__3062;
    wire N__3053;
    wire N__3050;
    wire N__3049;
    wire N__3046;
    wire N__3045;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3008;
    wire N__3005;
    wire N__3004;
    wire N__3003;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2966;
    wire N__2963;
    wire N__2962;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2954;
    wire N__2953;
    wire N__2950;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2921;
    wire N__2918;
    wire N__2917;
    wire N__2916;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2898;
    wire N__2895;
    wire N__2888;
    wire N__2885;
    wire N__2884;
    wire N__2883;
    wire N__2882;
    wire N__2881;
    wire N__2878;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2862;
    wire N__2859;
    wire N__2852;
    wire N__2849;
    wire N__2848;
    wire N__2847;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2836;
    wire N__2833;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2782;
    wire N__2779;
    wire N__2774;
    wire N__2771;
    wire N__2770;
    wire N__2769;
    wire N__2766;
    wire N__2765;
    wire N__2764;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2746;
    wire N__2743;
    wire N__2732;
    wire N__2731;
    wire N__2730;
    wire N__2729;
    wire N__2728;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2696;
    wire N__2693;
    wire N__2692;
    wire N__2691;
    wire N__2690;
    wire N__2687;
    wire N__2682;
    wire N__2679;
    wire N__2672;
    wire N__2671;
    wire N__2670;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2648;
    wire N__2647;
    wire N__2646;
    wire N__2645;
    wire N__2644;
    wire N__2641;
    wire N__2632;
    wire N__2629;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2591;
    wire N__2588;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2524;
    wire N__2523;
    wire N__2520;
    wire N__2515;
    wire N__2510;
    wire N__2509;
    wire N__2508;
    wire N__2507;
    wire N__2504;
    wire N__2497;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2467;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2419;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2353;
    wire N__2350;
    wire N__2349;
    wire N__2348;
    wire N__2347;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2335;
    wire N__2330;
    wire N__2327;
    wire N__2322;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2263;
    wire N__2262;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2225;
    wire VCCG0;
    wire \Clock50MHz.PixelClock ;
    wire Clock12MHz_c;
    wire GNDG0;
    wire bfn_7_1_0_;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0;
    wire bfn_7_2_0_;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_i;
    wire un5_beamx_0_a2_3_cascade_;
    wire un5_beamx_0_a2_5_cascade_;
    wire bfn_7_7_0_;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire un5_beamx;
    wire bfn_7_8_0_;
    wire bfn_8_1_0_;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_i;
    wire bfn_8_2_0_;
    wire un5_visiblex_cry_4;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un47_sum;
    wire un5_visiblex_cry_7;
    wire un5_visiblex_cry_8;
    wire un1_beamX_if_generate_plus_mult1_un40_sum;
    wire bfn_8_3_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_8_4_0_;
    wire un8_beamx_cry_9;
    wire beamXZ0Z_2;
    wire beamXZ0Z_1;
    wire beamXZ0Z_0;
    wire beamXZ0Z_7;
    wire beamXZ0Z_8;
    wire beamXZ0Z_9;
    wire Pixel_0_sqmuxa_i_2_1_cascade_;
    wire un1_beamylto9_0_a2_1_cascade_;
    wire VSync_c;
    wire N_84_cascade_;
    wire N_132;
    wire Pixel_0_sqmuxa_i_2;
    wire N_101_cascade_;
    wire Pixel_0_sqmuxa_i_1;
    wire un1_beamylto9_0_a2_1;
    wire Pixel_0_sqmuxa_i_4_cascade_;
    wire N_99;
    wire bfn_8_6_0_;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_;
    wire N_98;
    wire beamYZ0Z_0;
    wire bfn_8_7_0_;
    wire beamYZ0Z_1;
    wire un5_visibley_cry_0;
    wire beamYZ0Z_2;
    wire un5_visibley_cry_1;
    wire beamYZ0Z_3;
    wire un5_visibley_cry_2;
    wire beamYZ0Z_4;
    wire un5_visibley_cry_3;
    wire beamYZ0Z_5;
    wire un5_visibley_cry_4;
    wire beamYZ0Z_6;
    wire un5_visibley_cry_5;
    wire beamYZ0Z_7;
    wire un5_visibley_cry_6;
    wire un5_visibley_cry_7;
    wire beamYZ0Z_8;
    wire bfn_8_8_0_;
    wire beamYZ0Z_9;
    wire un5_visibley_cry_8;
    wire bfn_9_1_0_;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un54_sum;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_i;
    wire bfn_9_2_0_;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un61_sum;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_i;
    wire un1_beamX_if_generate_plus_mult1_un68_sum;
    wire bfn_9_3_0_;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_i;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_;
    wire Pixel_1_RNOZ0Z_7;
    wire un5_visiblex_i;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0;
    wire un5_visiblex_i_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6;
    wire un3_beamx_i_i_a2_4;
    wire un3_beamx_i_i_a2_5_cascade_;
    wire beamX_RNI5457Z0Z_1;
    wire beamXZ0Z_4;
    wire beamXZ0Z_6;
    wire beamXZ0Z_5;
    wire N_97;
    wire N_87;
    wire N_130_cascade_;
    wire beamXZ0Z_10;
    wire HSync_c;
    wire bfn_9_5_0_;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un47_sum;
    wire bfn_9_6_0_;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un40_sum;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_i_0;
    wire bfn_9_7_0_;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0;
    wire CONSTANT_ONE_NET;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_axb_6;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO;
    wire un1_visibley_if_generate_plus_mult1_un26_sum;
    wire un5_visibley_cry_8_c_RNI3O5CZ0Z_0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_i_0;
    wire un5_visibley_cry_0_c_RNIJVSBZ0;
    wire N_8_cascade_;
    wire Pixel_0_sqmuxa_i_5;
    wire N_94;
    wire N_49_cascade_;
    wire N_59;
    wire Pixel_c;
    wire PixelClock_g;
    wire un1_visibley_if_generate_plus_mult1_un75_sum;
    wire bfn_11_4_0_;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_3;
    wire Pixel_1_RNOZ0Z_6;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32;
    wire G_7_0_a4_0_0;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1;
    wire N_11;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_i_0;
    wire bfn_11_5_0_;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_i_0;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un54_sum;
    wire un1_visibley_if_generate_plus_mult1_un68_sum;
    wire bfn_12_4_0_;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_i_0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum;
    wire bfn_12_5_0_;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_i_0;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_i_7;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__2234),
            .RESETB(N__4061),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__4782),
            .DIN(N__4781),
            .DOUT(N__4780),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__4782),
            .PADOUT(N__4781),
            .PADIN(N__4780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4217),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__4773),
            .DIN(N__4772),
            .DOUT(N__4771),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__4773),
            .PADOUT(N__4772),
            .PADIN(N__4771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__4764),
            .DIN(N__4763),
            .DOUT(N__4762),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__4764),
            .PADOUT(N__4763),
            .PADIN(N__4762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__4755),
            .DIN(N__4754),
            .DOUT(N__4753),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__4755),
            .PADOUT(N__4754),
            .PADIN(N__4753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__4746),
            .DIN(N__4745),
            .DOUT(N__4744),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__4746),
            .PADOUT(N__4745),
            .PADIN(N__4744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__4737),
            .DIN(N__4736),
            .DOUT(N__4735),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__4737),
            .PADOUT(N__4736),
            .PADIN(N__4735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__4728),
            .DIN(N__4727),
            .DOUT(N__4726),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__4728),
            .PADOUT(N__4727),
            .PADIN(N__4726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1025 (
            .O(N__4709),
            .I(N__4705));
    InMux I__1024 (
            .O(N__4708),
            .I(N__4702));
    LocalMux I__1023 (
            .O(N__4705),
            .I(N__4699));
    LocalMux I__1022 (
            .O(N__4702),
            .I(N__4696));
    Span4Mux_v I__1021 (
            .O(N__4699),
            .I(N__4693));
    Span4Mux_s3_h I__1020 (
            .O(N__4696),
            .I(N__4690));
    Odrv4 I__1019 (
            .O(N__4693),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1018 (
            .O(N__4690),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1017 (
            .O(N__4685),
            .I(N__4682));
    InMux I__1016 (
            .O(N__4682),
            .I(N__4679));
    LocalMux I__1015 (
            .O(N__4679),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__1014 (
            .O(N__4676),
            .I(N__4673));
    LocalMux I__1013 (
            .O(N__4673),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8));
    InMux I__1012 (
            .O(N__4670),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__1011 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__1010 (
            .O(N__4664),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4));
    CascadeMux I__1009 (
            .O(N__4661),
            .I(N__4658));
    InMux I__1008 (
            .O(N__4658),
            .I(N__4655));
    LocalMux I__1007 (
            .O(N__4655),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0));
    InMux I__1006 (
            .O(N__4652),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__1005 (
            .O(N__4649),
            .I(N__4645));
    InMux I__1004 (
            .O(N__4648),
            .I(N__4636));
    InMux I__1003 (
            .O(N__4645),
            .I(N__4636));
    InMux I__1002 (
            .O(N__4644),
            .I(N__4636));
    InMux I__1001 (
            .O(N__4643),
            .I(N__4633));
    LocalMux I__1000 (
            .O(N__4636),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8));
    LocalMux I__999 (
            .O(N__4633),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8));
    CascadeMux I__998 (
            .O(N__4628),
            .I(N__4625));
    InMux I__997 (
            .O(N__4625),
            .I(N__4622));
    LocalMux I__996 (
            .O(N__4622),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117));
    InMux I__995 (
            .O(N__4619),
            .I(N__4616));
    LocalMux I__994 (
            .O(N__4616),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0));
    InMux I__993 (
            .O(N__4613),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__992 (
            .O(N__4610),
            .I(N__4607));
    LocalMux I__991 (
            .O(N__4607),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78));
    CascadeMux I__990 (
            .O(N__4604),
            .I(N__4601));
    InMux I__989 (
            .O(N__4601),
            .I(N__4598));
    LocalMux I__988 (
            .O(N__4598),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__987 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__986 (
            .O(N__4592),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__985 (
            .O(N__4589),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__984 (
            .O(N__4586),
            .I(N__4583));
    LocalMux I__983 (
            .O(N__4583),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__982 (
            .O(N__4580),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__981 (
            .O(N__4577),
            .I(N__4573));
    InMux I__980 (
            .O(N__4576),
            .I(N__4564));
    InMux I__979 (
            .O(N__4573),
            .I(N__4564));
    InMux I__978 (
            .O(N__4572),
            .I(N__4564));
    InMux I__977 (
            .O(N__4571),
            .I(N__4561));
    LocalMux I__976 (
            .O(N__4564),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0));
    LocalMux I__975 (
            .O(N__4561),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0));
    CascadeMux I__974 (
            .O(N__4556),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_));
    CascadeMux I__973 (
            .O(N__4553),
            .I(N__4550));
    InMux I__972 (
            .O(N__4550),
            .I(N__4547));
    LocalMux I__971 (
            .O(N__4547),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_i_7));
    CascadeMux I__970 (
            .O(N__4544),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_));
    InMux I__969 (
            .O(N__4541),
            .I(N__4535));
    InMux I__968 (
            .O(N__4540),
            .I(N__4535));
    LocalMux I__967 (
            .O(N__4535),
            .I(N__4532));
    Span4Mux_s3_h I__966 (
            .O(N__4532),
            .I(N__4529));
    Odrv4 I__965 (
            .O(N__4529),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum));
    InMux I__964 (
            .O(N__4526),
            .I(N__4522));
    InMux I__963 (
            .O(N__4525),
            .I(N__4519));
    LocalMux I__962 (
            .O(N__4522),
            .I(N__4514));
    LocalMux I__961 (
            .O(N__4519),
            .I(N__4514));
    Span4Mux_s3_h I__960 (
            .O(N__4514),
            .I(N__4511));
    Odrv4 I__959 (
            .O(N__4511),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum));
    CascadeMux I__958 (
            .O(N__4508),
            .I(N__4505));
    InMux I__957 (
            .O(N__4505),
            .I(N__4502));
    LocalMux I__956 (
            .O(N__4502),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0));
    InMux I__955 (
            .O(N__4499),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__954 (
            .O(N__4496),
            .I(N__4493));
    LocalMux I__953 (
            .O(N__4493),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0));
    InMux I__952 (
            .O(N__4490),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__951 (
            .O(N__4487),
            .I(N__4484));
    LocalMux I__950 (
            .O(N__4484),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0));
    InMux I__949 (
            .O(N__4481),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__948 (
            .O(N__4478),
            .I(N__4475));
    InMux I__947 (
            .O(N__4475),
            .I(N__4472));
    LocalMux I__946 (
            .O(N__4472),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__945 (
            .O(N__4469),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__944 (
            .O(N__4466),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__943 (
            .O(N__4463),
            .I(N__4458));
    CascadeMux I__942 (
            .O(N__4462),
            .I(N__4454));
    InMux I__941 (
            .O(N__4461),
            .I(N__4450));
    InMux I__940 (
            .O(N__4458),
            .I(N__4441));
    InMux I__939 (
            .O(N__4457),
            .I(N__4441));
    InMux I__938 (
            .O(N__4454),
            .I(N__4441));
    InMux I__937 (
            .O(N__4453),
            .I(N__4441));
    LocalMux I__936 (
            .O(N__4450),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21));
    LocalMux I__935 (
            .O(N__4441),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21));
    CascadeMux I__934 (
            .O(N__4436),
            .I(N__4433));
    InMux I__933 (
            .O(N__4433),
            .I(N__4430));
    LocalMux I__932 (
            .O(N__4430),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__931 (
            .O(N__4427),
            .I(N__4424));
    LocalMux I__930 (
            .O(N__4424),
            .I(N__4421));
    Odrv12 I__929 (
            .O(N__4421),
            .I(G_7_0_a4_0_0));
    InMux I__928 (
            .O(N__4418),
            .I(N__4414));
    InMux I__927 (
            .O(N__4417),
            .I(N__4411));
    LocalMux I__926 (
            .O(N__4414),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21));
    LocalMux I__925 (
            .O(N__4411),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21));
    CascadeMux I__924 (
            .O(N__4406),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_));
    InMux I__923 (
            .O(N__4403),
            .I(N__4399));
    InMux I__922 (
            .O(N__4402),
            .I(N__4396));
    LocalMux I__921 (
            .O(N__4399),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1));
    LocalMux I__920 (
            .O(N__4396),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1));
    InMux I__919 (
            .O(N__4391),
            .I(N__4388));
    LocalMux I__918 (
            .O(N__4388),
            .I(N_11));
    InMux I__917 (
            .O(N__4385),
            .I(N__4382));
    LocalMux I__916 (
            .O(N__4382),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_i_0));
    CascadeMux I__915 (
            .O(N__4379),
            .I(N__4376));
    InMux I__914 (
            .O(N__4376),
            .I(N__4373));
    LocalMux I__913 (
            .O(N__4373),
            .I(N__4370));
    Odrv12 I__912 (
            .O(N__4370),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__911 (
            .O(N__4367),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__910 (
            .O(N__4364),
            .I(N__4361));
    LocalMux I__909 (
            .O(N__4361),
            .I(N__4358));
    Odrv4 I__908 (
            .O(N__4358),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2));
    InMux I__907 (
            .O(N__4355),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__906 (
            .O(N__4352),
            .I(N__4348));
    InMux I__905 (
            .O(N__4351),
            .I(N__4340));
    InMux I__904 (
            .O(N__4348),
            .I(N__4340));
    InMux I__903 (
            .O(N__4347),
            .I(N__4340));
    LocalMux I__902 (
            .O(N__4340),
            .I(N__4336));
    InMux I__901 (
            .O(N__4339),
            .I(N__4333));
    Odrv4 I__900 (
            .O(N__4336),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94));
    LocalMux I__899 (
            .O(N__4333),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94));
    CascadeMux I__898 (
            .O(N__4328),
            .I(N__4325));
    InMux I__897 (
            .O(N__4325),
            .I(N__4322));
    LocalMux I__896 (
            .O(N__4322),
            .I(N__4319));
    Odrv4 I__895 (
            .O(N__4319),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3));
    InMux I__894 (
            .O(N__4316),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__893 (
            .O(N__4313),
            .I(N__4310));
    LocalMux I__892 (
            .O(N__4310),
            .I(N__4307));
    Odrv4 I__891 (
            .O(N__4307),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3));
    CascadeMux I__890 (
            .O(N__4304),
            .I(N__4301));
    InMux I__889 (
            .O(N__4301),
            .I(N__4298));
    LocalMux I__888 (
            .O(N__4298),
            .I(N__4295));
    Odrv4 I__887 (
            .O(N__4295),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_i_7));
    InMux I__886 (
            .O(N__4292),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__885 (
            .O(N__4289),
            .I(N__4286));
    LocalMux I__884 (
            .O(N__4286),
            .I(N__4283));
    Odrv4 I__883 (
            .O(N__4283),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__882 (
            .O(N__4280),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__881 (
            .O(N__4277),
            .I(N__4274));
    LocalMux I__880 (
            .O(N__4274),
            .I(N__4269));
    InMux I__879 (
            .O(N__4273),
            .I(N__4266));
    InMux I__878 (
            .O(N__4272),
            .I(N__4263));
    Span4Mux_s3_h I__877 (
            .O(N__4269),
            .I(N__4258));
    LocalMux I__876 (
            .O(N__4266),
            .I(N__4258));
    LocalMux I__875 (
            .O(N__4263),
            .I(un5_visibley_cry_0_c_RNIJVSBZ0));
    Odrv4 I__874 (
            .O(N__4258),
            .I(un5_visibley_cry_0_c_RNIJVSBZ0));
    CascadeMux I__873 (
            .O(N__4253),
            .I(N_8_cascade_));
    InMux I__872 (
            .O(N__4250),
            .I(N__4247));
    LocalMux I__871 (
            .O(N__4247),
            .I(N__4244));
    Span4Mux_s3_h I__870 (
            .O(N__4244),
            .I(N__4241));
    Odrv4 I__869 (
            .O(N__4241),
            .I(Pixel_0_sqmuxa_i_5));
    InMux I__868 (
            .O(N__4238),
            .I(N__4235));
    LocalMux I__867 (
            .O(N__4235),
            .I(N__4232));
    Odrv4 I__866 (
            .O(N__4232),
            .I(N_94));
    CascadeMux I__865 (
            .O(N__4229),
            .I(N_49_cascade_));
    InMux I__864 (
            .O(N__4226),
            .I(N__4223));
    LocalMux I__863 (
            .O(N__4223),
            .I(N__4220));
    Odrv4 I__862 (
            .O(N__4220),
            .I(N_59));
    IoInMux I__861 (
            .O(N__4217),
            .I(N__4214));
    LocalMux I__860 (
            .O(N__4214),
            .I(N__4210));
    IoInMux I__859 (
            .O(N__4213),
            .I(N__4207));
    Span4Mux_s2_v I__858 (
            .O(N__4210),
            .I(N__4204));
    LocalMux I__857 (
            .O(N__4207),
            .I(N__4201));
    Span4Mux_v I__856 (
            .O(N__4204),
            .I(N__4198));
    IoSpan4Mux I__855 (
            .O(N__4201),
            .I(N__4195));
    Span4Mux_v I__854 (
            .O(N__4198),
            .I(N__4192));
    Span4Mux_s2_v I__853 (
            .O(N__4195),
            .I(N__4189));
    Odrv4 I__852 (
            .O(N__4192),
            .I(Pixel_c));
    Odrv4 I__851 (
            .O(N__4189),
            .I(Pixel_c));
    ClkMux I__850 (
            .O(N__4184),
            .I(N__4160));
    ClkMux I__849 (
            .O(N__4183),
            .I(N__4160));
    ClkMux I__848 (
            .O(N__4182),
            .I(N__4160));
    ClkMux I__847 (
            .O(N__4181),
            .I(N__4160));
    ClkMux I__846 (
            .O(N__4180),
            .I(N__4160));
    ClkMux I__845 (
            .O(N__4179),
            .I(N__4160));
    ClkMux I__844 (
            .O(N__4178),
            .I(N__4160));
    ClkMux I__843 (
            .O(N__4177),
            .I(N__4160));
    GlobalMux I__842 (
            .O(N__4160),
            .I(N__4157));
    gio2CtrlBuf I__841 (
            .O(N__4157),
            .I(PixelClock_g));
    CascadeMux I__840 (
            .O(N__4154),
            .I(N__4151));
    InMux I__839 (
            .O(N__4151),
            .I(N__4146));
    InMux I__838 (
            .O(N__4150),
            .I(N__4143));
    InMux I__837 (
            .O(N__4149),
            .I(N__4140));
    LocalMux I__836 (
            .O(N__4146),
            .I(N__4137));
    LocalMux I__835 (
            .O(N__4143),
            .I(N__4132));
    LocalMux I__834 (
            .O(N__4140),
            .I(N__4132));
    Span4Mux_s3_h I__833 (
            .O(N__4137),
            .I(N__4129));
    Span4Mux_s3_h I__832 (
            .O(N__4132),
            .I(N__4126));
    Odrv4 I__831 (
            .O(N__4129),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum));
    Odrv4 I__830 (
            .O(N__4126),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum));
    InMux I__829 (
            .O(N__4121),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__828 (
            .O(N__4118),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__827 (
            .O(N__4115),
            .I(N__4112));
    LocalMux I__826 (
            .O(N__4112),
            .I(Pixel_1_RNOZ0Z_6));
    InMux I__825 (
            .O(N__4109),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__824 (
            .O(N__4106),
            .I(N__4103));
    InMux I__823 (
            .O(N__4103),
            .I(N__4100));
    LocalMux I__822 (
            .O(N__4100),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0));
    InMux I__821 (
            .O(N__4097),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__820 (
            .O(N__4094),
            .I(N__4091));
    LocalMux I__819 (
            .O(N__4091),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32));
    CascadeMux I__818 (
            .O(N__4088),
            .I(N__4085));
    InMux I__817 (
            .O(N__4085),
            .I(N__4082));
    LocalMux I__816 (
            .O(N__4082),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0));
    InMux I__815 (
            .O(N__4079),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__814 (
            .O(N__4076),
            .I(N__4073));
    LocalMux I__813 (
            .O(N__4073),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0));
    InMux I__812 (
            .O(N__4070),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__811 (
            .O(N__4067),
            .I(N__4064));
    LocalMux I__810 (
            .O(N__4064),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0));
    IoInMux I__809 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__808 (
            .O(N__4058),
            .I(N__4049));
    CascadeMux I__807 (
            .O(N__4057),
            .I(N__4046));
    CascadeMux I__806 (
            .O(N__4056),
            .I(N__4043));
    CascadeMux I__805 (
            .O(N__4055),
            .I(N__4040));
    CascadeMux I__804 (
            .O(N__4054),
            .I(N__4037));
    InMux I__803 (
            .O(N__4053),
            .I(N__4032));
    CascadeMux I__802 (
            .O(N__4052),
            .I(N__4028));
    IoSpan4Mux I__801 (
            .O(N__4049),
            .I(N__4025));
    InMux I__800 (
            .O(N__4046),
            .I(N__4020));
    InMux I__799 (
            .O(N__4043),
            .I(N__4020));
    InMux I__798 (
            .O(N__4040),
            .I(N__4017));
    InMux I__797 (
            .O(N__4037),
            .I(N__4012));
    InMux I__796 (
            .O(N__4036),
            .I(N__4012));
    InMux I__795 (
            .O(N__4035),
            .I(N__4009));
    LocalMux I__794 (
            .O(N__4032),
            .I(N__4006));
    InMux I__793 (
            .O(N__4031),
            .I(N__4003));
    InMux I__792 (
            .O(N__4028),
            .I(N__3997));
    Span4Mux_s0_v I__791 (
            .O(N__4025),
            .I(N__3994));
    LocalMux I__790 (
            .O(N__4020),
            .I(N__3991));
    LocalMux I__789 (
            .O(N__4017),
            .I(N__3986));
    LocalMux I__788 (
            .O(N__4012),
            .I(N__3986));
    LocalMux I__787 (
            .O(N__4009),
            .I(N__3979));
    Span4Mux_v I__786 (
            .O(N__4006),
            .I(N__3979));
    LocalMux I__785 (
            .O(N__4003),
            .I(N__3979));
    InMux I__784 (
            .O(N__4002),
            .I(N__3972));
    InMux I__783 (
            .O(N__4001),
            .I(N__3972));
    InMux I__782 (
            .O(N__4000),
            .I(N__3972));
    LocalMux I__781 (
            .O(N__3997),
            .I(N__3966));
    Span4Mux_v I__780 (
            .O(N__3994),
            .I(N__3957));
    Span4Mux_v I__779 (
            .O(N__3991),
            .I(N__3957));
    Span4Mux_v I__778 (
            .O(N__3986),
            .I(N__3957));
    Span4Mux_v I__777 (
            .O(N__3979),
            .I(N__3957));
    LocalMux I__776 (
            .O(N__3972),
            .I(N__3954));
    InMux I__775 (
            .O(N__3971),
            .I(N__3951));
    InMux I__774 (
            .O(N__3970),
            .I(N__3946));
    InMux I__773 (
            .O(N__3969),
            .I(N__3946));
    Odrv12 I__772 (
            .O(N__3966),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__771 (
            .O(N__3957),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__770 (
            .O(N__3954),
            .I(CONSTANT_ONE_NET));
    LocalMux I__769 (
            .O(N__3951),
            .I(CONSTANT_ONE_NET));
    LocalMux I__768 (
            .O(N__3946),
            .I(CONSTANT_ONE_NET));
    InMux I__767 (
            .O(N__3935),
            .I(N__3932));
    LocalMux I__766 (
            .O(N__3932),
            .I(N__3929));
    Odrv4 I__765 (
            .O(N__3929),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0));
    InMux I__764 (
            .O(N__3926),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__763 (
            .O(N__3923),
            .I(N__3919));
    InMux I__762 (
            .O(N__3922),
            .I(N__3916));
    InMux I__761 (
            .O(N__3919),
            .I(N__3913));
    LocalMux I__760 (
            .O(N__3916),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_axb_6));
    LocalMux I__759 (
            .O(N__3913),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_axb_6));
    InMux I__758 (
            .O(N__3908),
            .I(N__3905));
    LocalMux I__757 (
            .O(N__3905),
            .I(N__3902));
    Odrv4 I__756 (
            .O(N__3902),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__755 (
            .O(N__3899),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__754 (
            .O(N__3896),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_6));
    CascadeMux I__753 (
            .O(N__3893),
            .I(N__3890));
    InMux I__752 (
            .O(N__3890),
            .I(N__3887));
    LocalMux I__751 (
            .O(N__3887),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO));
    InMux I__750 (
            .O(N__3884),
            .I(N__3877));
    InMux I__749 (
            .O(N__3883),
            .I(N__3877));
    InMux I__748 (
            .O(N__3882),
            .I(N__3874));
    LocalMux I__747 (
            .O(N__3877),
            .I(N__3867));
    LocalMux I__746 (
            .O(N__3874),
            .I(N__3867));
    InMux I__745 (
            .O(N__3873),
            .I(N__3862));
    InMux I__744 (
            .O(N__3872),
            .I(N__3862));
    Odrv4 I__743 (
            .O(N__3867),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum));
    LocalMux I__742 (
            .O(N__3862),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum));
    CascadeMux I__741 (
            .O(N__3857),
            .I(N__3854));
    InMux I__740 (
            .O(N__3854),
            .I(N__3851));
    LocalMux I__739 (
            .O(N__3851),
            .I(un5_visibley_cry_8_c_RNI3O5CZ0Z_0));
    InMux I__738 (
            .O(N__3848),
            .I(N__3842));
    InMux I__737 (
            .O(N__3847),
            .I(N__3842));
    LocalMux I__736 (
            .O(N__3842),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum));
    InMux I__735 (
            .O(N__3839),
            .I(N__3836));
    LocalMux I__734 (
            .O(N__3836),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_i_0));
    InMux I__733 (
            .O(N__3833),
            .I(N__3830));
    LocalMux I__732 (
            .O(N__3830),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1));
    InMux I__731 (
            .O(N__3827),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__730 (
            .O(N__3824),
            .I(N__3821));
    InMux I__729 (
            .O(N__3821),
            .I(N__3818));
    LocalMux I__728 (
            .O(N__3818),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1));
    InMux I__727 (
            .O(N__3815),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__726 (
            .O(N__3812),
            .I(N__3809));
    LocalMux I__725 (
            .O(N__3809),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1));
    InMux I__724 (
            .O(N__3806),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__723 (
            .O(N__3803),
            .I(N__3800));
    InMux I__722 (
            .O(N__3800),
            .I(N__3797));
    LocalMux I__721 (
            .O(N__3797),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_i_7));
    InMux I__720 (
            .O(N__3794),
            .I(N__3791));
    LocalMux I__719 (
            .O(N__3791),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_axb_7));
    InMux I__718 (
            .O(N__3788),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5));
    CascadeMux I__717 (
            .O(N__3785),
            .I(N__3780));
    CascadeMux I__716 (
            .O(N__3784),
            .I(N__3777));
    CascadeMux I__715 (
            .O(N__3783),
            .I(N__3773));
    InMux I__714 (
            .O(N__3780),
            .I(N__3764));
    InMux I__713 (
            .O(N__3777),
            .I(N__3764));
    InMux I__712 (
            .O(N__3776),
            .I(N__3764));
    InMux I__711 (
            .O(N__3773),
            .I(N__3764));
    LocalMux I__710 (
            .O(N__3764),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0));
    InMux I__709 (
            .O(N__3761),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__708 (
            .O(N__3758),
            .I(N__3754));
    InMux I__707 (
            .O(N__3757),
            .I(N__3745));
    InMux I__706 (
            .O(N__3754),
            .I(N__3745));
    InMux I__705 (
            .O(N__3753),
            .I(N__3745));
    InMux I__704 (
            .O(N__3752),
            .I(N__3742));
    LocalMux I__703 (
            .O(N__3745),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1));
    LocalMux I__702 (
            .O(N__3742),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1));
    CascadeMux I__701 (
            .O(N__3737),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_));
    CascadeMux I__700 (
            .O(N__3734),
            .I(N__3731));
    InMux I__699 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__698 (
            .O(N__3728),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__697 (
            .O(N__3725),
            .I(N__3719));
    InMux I__696 (
            .O(N__3724),
            .I(N__3719));
    LocalMux I__695 (
            .O(N__3719),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum));
    CascadeMux I__694 (
            .O(N__3716),
            .I(N__3713));
    InMux I__693 (
            .O(N__3713),
            .I(N__3710));
    LocalMux I__692 (
            .O(N__3710),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__691 (
            .O(N__3707),
            .I(N__3700));
    InMux I__690 (
            .O(N__3706),
            .I(N__3700));
    InMux I__689 (
            .O(N__3705),
            .I(N__3697));
    LocalMux I__688 (
            .O(N__3700),
            .I(N_87));
    LocalMux I__687 (
            .O(N__3697),
            .I(N_87));
    CascadeMux I__686 (
            .O(N__3692),
            .I(N_130_cascade_));
    CascadeMux I__685 (
            .O(N__3689),
            .I(N__3683));
    InMux I__684 (
            .O(N__3688),
            .I(N__3680));
    InMux I__683 (
            .O(N__3687),
            .I(N__3677));
    InMux I__682 (
            .O(N__3686),
            .I(N__3674));
    InMux I__681 (
            .O(N__3683),
            .I(N__3671));
    LocalMux I__680 (
            .O(N__3680),
            .I(beamXZ0Z_10));
    LocalMux I__679 (
            .O(N__3677),
            .I(beamXZ0Z_10));
    LocalMux I__678 (
            .O(N__3674),
            .I(beamXZ0Z_10));
    LocalMux I__677 (
            .O(N__3671),
            .I(beamXZ0Z_10));
    IoInMux I__676 (
            .O(N__3662),
            .I(N__3659));
    LocalMux I__675 (
            .O(N__3659),
            .I(N__3656));
    IoSpan4Mux I__674 (
            .O(N__3656),
            .I(N__3653));
    Sp12to4 I__673 (
            .O(N__3653),
            .I(N__3649));
    IoInMux I__672 (
            .O(N__3652),
            .I(N__3646));
    Span12Mux_v I__671 (
            .O(N__3649),
            .I(N__3643));
    LocalMux I__670 (
            .O(N__3646),
            .I(N__3640));
    Odrv12 I__669 (
            .O(N__3643),
            .I(HSync_c));
    Odrv12 I__668 (
            .O(N__3640),
            .I(HSync_c));
    InMux I__667 (
            .O(N__3635),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__666 (
            .O(N__3632),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__665 (
            .O(N__3629),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__664 (
            .O(N__3626),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__663 (
            .O(N__3623),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__662 (
            .O(N__3620),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_));
    InMux I__661 (
            .O(N__3617),
            .I(N__3611));
    InMux I__660 (
            .O(N__3616),
            .I(N__3611));
    LocalMux I__659 (
            .O(N__3611),
            .I(N__3608));
    Odrv4 I__658 (
            .O(N__3608),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum));
    InMux I__657 (
            .O(N__3605),
            .I(N__3602));
    LocalMux I__656 (
            .O(N__3602),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__655 (
            .O(N__3599),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__654 (
            .O(N__3596),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_));
    InMux I__653 (
            .O(N__3593),
            .I(N__3590));
    LocalMux I__652 (
            .O(N__3590),
            .I(Pixel_1_RNOZ0Z_7));
    InMux I__651 (
            .O(N__3587),
            .I(N__3578));
    InMux I__650 (
            .O(N__3586),
            .I(N__3578));
    InMux I__649 (
            .O(N__3585),
            .I(N__3578));
    LocalMux I__648 (
            .O(N__3578),
            .I(un5_visiblex_i));
    InMux I__647 (
            .O(N__3575),
            .I(N__3569));
    InMux I__646 (
            .O(N__3574),
            .I(N__3569));
    LocalMux I__645 (
            .O(N__3569),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0));
    CascadeMux I__644 (
            .O(N__3566),
            .I(un5_visiblex_i_cascade_));
    InMux I__643 (
            .O(N__3563),
            .I(N__3560));
    LocalMux I__642 (
            .O(N__3560),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6));
    InMux I__641 (
            .O(N__3557),
            .I(N__3554));
    LocalMux I__640 (
            .O(N__3554),
            .I(un3_beamx_i_i_a2_4));
    CascadeMux I__639 (
            .O(N__3551),
            .I(un3_beamx_i_i_a2_5_cascade_));
    CEMux I__638 (
            .O(N__3548),
            .I(N__3545));
    LocalMux I__637 (
            .O(N__3545),
            .I(N__3540));
    CEMux I__636 (
            .O(N__3544),
            .I(N__3537));
    CEMux I__635 (
            .O(N__3543),
            .I(N__3533));
    Span4Mux_v I__634 (
            .O(N__3540),
            .I(N__3528));
    LocalMux I__633 (
            .O(N__3537),
            .I(N__3528));
    InMux I__632 (
            .O(N__3536),
            .I(N__3525));
    LocalMux I__631 (
            .O(N__3533),
            .I(N__3520));
    Span4Mux_h I__630 (
            .O(N__3528),
            .I(N__3517));
    LocalMux I__629 (
            .O(N__3525),
            .I(N__3514));
    InMux I__628 (
            .O(N__3524),
            .I(N__3509));
    InMux I__627 (
            .O(N__3523),
            .I(N__3509));
    Span4Mux_v I__626 (
            .O(N__3520),
            .I(N__3504));
    Span4Mux_v I__625 (
            .O(N__3517),
            .I(N__3504));
    Odrv4 I__624 (
            .O(N__3514),
            .I(beamX_RNI5457Z0Z_1));
    LocalMux I__623 (
            .O(N__3509),
            .I(beamX_RNI5457Z0Z_1));
    Odrv4 I__622 (
            .O(N__3504),
            .I(beamX_RNI5457Z0Z_1));
    InMux I__621 (
            .O(N__3497),
            .I(N__3490));
    InMux I__620 (
            .O(N__3496),
            .I(N__3486));
    InMux I__619 (
            .O(N__3495),
            .I(N__3481));
    InMux I__618 (
            .O(N__3494),
            .I(N__3481));
    InMux I__617 (
            .O(N__3493),
            .I(N__3478));
    LocalMux I__616 (
            .O(N__3490),
            .I(N__3475));
    InMux I__615 (
            .O(N__3489),
            .I(N__3472));
    LocalMux I__614 (
            .O(N__3486),
            .I(beamXZ0Z_4));
    LocalMux I__613 (
            .O(N__3481),
            .I(beamXZ0Z_4));
    LocalMux I__612 (
            .O(N__3478),
            .I(beamXZ0Z_4));
    Odrv4 I__611 (
            .O(N__3475),
            .I(beamXZ0Z_4));
    LocalMux I__610 (
            .O(N__3472),
            .I(beamXZ0Z_4));
    CascadeMux I__609 (
            .O(N__3461),
            .I(N__3455));
    InMux I__608 (
            .O(N__3460),
            .I(N__3451));
    InMux I__607 (
            .O(N__3459),
            .I(N__3448));
    InMux I__606 (
            .O(N__3458),
            .I(N__3445));
    InMux I__605 (
            .O(N__3455),
            .I(N__3442));
    InMux I__604 (
            .O(N__3454),
            .I(N__3439));
    LocalMux I__603 (
            .O(N__3451),
            .I(beamXZ0Z_6));
    LocalMux I__602 (
            .O(N__3448),
            .I(beamXZ0Z_6));
    LocalMux I__601 (
            .O(N__3445),
            .I(beamXZ0Z_6));
    LocalMux I__600 (
            .O(N__3442),
            .I(beamXZ0Z_6));
    LocalMux I__599 (
            .O(N__3439),
            .I(beamXZ0Z_6));
    CascadeMux I__598 (
            .O(N__3428),
            .I(N__3424));
    InMux I__597 (
            .O(N__3427),
            .I(N__3418));
    InMux I__596 (
            .O(N__3424),
            .I(N__3413));
    InMux I__595 (
            .O(N__3423),
            .I(N__3413));
    InMux I__594 (
            .O(N__3422),
            .I(N__3410));
    InMux I__593 (
            .O(N__3421),
            .I(N__3407));
    LocalMux I__592 (
            .O(N__3418),
            .I(beamXZ0Z_5));
    LocalMux I__591 (
            .O(N__3413),
            .I(beamXZ0Z_5));
    LocalMux I__590 (
            .O(N__3410),
            .I(beamXZ0Z_5));
    LocalMux I__589 (
            .O(N__3407),
            .I(beamXZ0Z_5));
    InMux I__588 (
            .O(N__3398),
            .I(N__3394));
    CascadeMux I__587 (
            .O(N__3397),
            .I(N__3389));
    LocalMux I__586 (
            .O(N__3394),
            .I(N__3386));
    InMux I__585 (
            .O(N__3393),
            .I(N__3383));
    InMux I__584 (
            .O(N__3392),
            .I(N__3378));
    InMux I__583 (
            .O(N__3389),
            .I(N__3378));
    Odrv4 I__582 (
            .O(N__3386),
            .I(N_97));
    LocalMux I__581 (
            .O(N__3383),
            .I(N_97));
    LocalMux I__580 (
            .O(N__3378),
            .I(N_97));
    InMux I__579 (
            .O(N__3371),
            .I(N__3367));
    InMux I__578 (
            .O(N__3370),
            .I(N__3364));
    LocalMux I__577 (
            .O(N__3367),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1));
    LocalMux I__576 (
            .O(N__3364),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1));
    CascadeMux I__575 (
            .O(N__3359),
            .I(N__3356));
    InMux I__574 (
            .O(N__3356),
            .I(N__3353));
    LocalMux I__573 (
            .O(N__3353),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21));
    InMux I__572 (
            .O(N__3350),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__571 (
            .O(N__3347),
            .I(N__3341));
    InMux I__570 (
            .O(N__3346),
            .I(N__3341));
    LocalMux I__569 (
            .O(N__3341),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__568 (
            .O(N__3338),
            .I(N__3335));
    InMux I__567 (
            .O(N__3335),
            .I(N__3332));
    LocalMux I__566 (
            .O(N__3332),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1));
    InMux I__565 (
            .O(N__3329),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__564 (
            .O(N__3326),
            .I(N__3323));
    LocalMux I__563 (
            .O(N__3323),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__562 (
            .O(N__3320),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__561 (
            .O(N__3317),
            .I(N__3313));
    InMux I__560 (
            .O(N__3316),
            .I(N__3310));
    LocalMux I__559 (
            .O(N__3313),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum));
    LocalMux I__558 (
            .O(N__3310),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum));
    CascadeMux I__557 (
            .O(N__3305),
            .I(N__3302));
    InMux I__556 (
            .O(N__3302),
            .I(N__3299));
    LocalMux I__555 (
            .O(N__3299),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_i));
    InMux I__554 (
            .O(N__3296),
            .I(N__3290));
    InMux I__553 (
            .O(N__3295),
            .I(N__3290));
    LocalMux I__552 (
            .O(N__3290),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum));
    CascadeMux I__551 (
            .O(N__3287),
            .I(N__3284));
    InMux I__550 (
            .O(N__3284),
            .I(N__3281));
    LocalMux I__549 (
            .O(N__3281),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_i));
    InMux I__548 (
            .O(N__3278),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__547 (
            .O(N__3275),
            .I(N__3272));
    LocalMux I__546 (
            .O(N__3272),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1));
    InMux I__545 (
            .O(N__3269),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5));
    CascadeMux I__544 (
            .O(N__3266),
            .I(N__3263));
    InMux I__543 (
            .O(N__3263),
            .I(N__3260));
    LocalMux I__542 (
            .O(N__3260),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2));
    CascadeMux I__541 (
            .O(N__3257),
            .I(N__3253));
    InMux I__540 (
            .O(N__3256),
            .I(N__3249));
    InMux I__539 (
            .O(N__3253),
            .I(N__3244));
    InMux I__538 (
            .O(N__3252),
            .I(N__3244));
    LocalMux I__537 (
            .O(N__3249),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843));
    LocalMux I__536 (
            .O(N__3244),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843));
    InMux I__535 (
            .O(N__3239),
            .I(N__3233));
    InMux I__534 (
            .O(N__3238),
            .I(N__3233));
    LocalMux I__533 (
            .O(N__3233),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__532 (
            .O(N__3230),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__531 (
            .O(N__3227),
            .I(N__3223));
    InMux I__530 (
            .O(N__3226),
            .I(N__3220));
    LocalMux I__529 (
            .O(N__3223),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0));
    LocalMux I__528 (
            .O(N__3220),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0));
    CascadeMux I__527 (
            .O(N__3215),
            .I(N__3212));
    InMux I__526 (
            .O(N__3212),
            .I(N__3209));
    LocalMux I__525 (
            .O(N__3209),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0));
    InMux I__524 (
            .O(N__3206),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__523 (
            .O(N__3203),
            .I(N__3197));
    InMux I__522 (
            .O(N__3202),
            .I(N__3197));
    LocalMux I__521 (
            .O(N__3197),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__520 (
            .O(N__3194),
            .I(N__3191));
    InMux I__519 (
            .O(N__3191),
            .I(N__3188));
    LocalMux I__518 (
            .O(N__3188),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0));
    InMux I__517 (
            .O(N__3185),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__516 (
            .O(N__3182),
            .I(N__3179));
    LocalMux I__515 (
            .O(N__3179),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__514 (
            .O(N__3176),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__513 (
            .O(N__3173),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_));
    CascadeMux I__512 (
            .O(N__3170),
            .I(N__3166));
    InMux I__511 (
            .O(N__3169),
            .I(N__3163));
    InMux I__510 (
            .O(N__3166),
            .I(N__3160));
    LocalMux I__509 (
            .O(N__3163),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum));
    LocalMux I__508 (
            .O(N__3160),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum));
    CascadeMux I__507 (
            .O(N__3155),
            .I(N__3152));
    InMux I__506 (
            .O(N__3152),
            .I(N__3149));
    LocalMux I__505 (
            .O(N__3149),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_i));
    InMux I__504 (
            .O(N__3146),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__503 (
            .O(N__3143),
            .I(N__3134));
    InMux I__502 (
            .O(N__3142),
            .I(N__3134));
    InMux I__501 (
            .O(N__3141),
            .I(N__3134));
    LocalMux I__500 (
            .O(N__3134),
            .I(N__3128));
    InMux I__499 (
            .O(N__3133),
            .I(N__3125));
    CascadeMux I__498 (
            .O(N__3132),
            .I(N__3122));
    InMux I__497 (
            .O(N__3131),
            .I(N__3119));
    Span4Mux_h I__496 (
            .O(N__3128),
            .I(N__3116));
    LocalMux I__495 (
            .O(N__3125),
            .I(N__3113));
    InMux I__494 (
            .O(N__3122),
            .I(N__3110));
    LocalMux I__493 (
            .O(N__3119),
            .I(beamYZ0Z_2));
    Odrv4 I__492 (
            .O(N__3116),
            .I(beamYZ0Z_2));
    Odrv4 I__491 (
            .O(N__3113),
            .I(beamYZ0Z_2));
    LocalMux I__490 (
            .O(N__3110),
            .I(beamYZ0Z_2));
    InMux I__489 (
            .O(N__3101),
            .I(un5_visibley_cry_1));
    CascadeMux I__488 (
            .O(N__3098),
            .I(N__3093));
    CascadeMux I__487 (
            .O(N__3097),
            .I(N__3090));
    InMux I__486 (
            .O(N__3096),
            .I(N__3085));
    InMux I__485 (
            .O(N__3093),
            .I(N__3082));
    InMux I__484 (
            .O(N__3090),
            .I(N__3079));
    CascadeMux I__483 (
            .O(N__3089),
            .I(N__3076));
    InMux I__482 (
            .O(N__3088),
            .I(N__3073));
    LocalMux I__481 (
            .O(N__3085),
            .I(N__3070));
    LocalMux I__480 (
            .O(N__3082),
            .I(N__3065));
    LocalMux I__479 (
            .O(N__3079),
            .I(N__3065));
    InMux I__478 (
            .O(N__3076),
            .I(N__3062));
    LocalMux I__477 (
            .O(N__3073),
            .I(beamYZ0Z_3));
    Odrv4 I__476 (
            .O(N__3070),
            .I(beamYZ0Z_3));
    Odrv4 I__475 (
            .O(N__3065),
            .I(beamYZ0Z_3));
    LocalMux I__474 (
            .O(N__3062),
            .I(beamYZ0Z_3));
    InMux I__473 (
            .O(N__3053),
            .I(un5_visibley_cry_2));
    CascadeMux I__472 (
            .O(N__3050),
            .I(N__3046));
    InMux I__471 (
            .O(N__3049),
            .I(N__3041));
    InMux I__470 (
            .O(N__3046),
            .I(N__3038));
    CascadeMux I__469 (
            .O(N__3045),
            .I(N__3034));
    InMux I__468 (
            .O(N__3044),
            .I(N__3031));
    LocalMux I__467 (
            .O(N__3041),
            .I(N__3028));
    LocalMux I__466 (
            .O(N__3038),
            .I(N__3025));
    InMux I__465 (
            .O(N__3037),
            .I(N__3022));
    InMux I__464 (
            .O(N__3034),
            .I(N__3019));
    LocalMux I__463 (
            .O(N__3031),
            .I(beamYZ0Z_4));
    Odrv4 I__462 (
            .O(N__3028),
            .I(beamYZ0Z_4));
    Odrv4 I__461 (
            .O(N__3025),
            .I(beamYZ0Z_4));
    LocalMux I__460 (
            .O(N__3022),
            .I(beamYZ0Z_4));
    LocalMux I__459 (
            .O(N__3019),
            .I(beamYZ0Z_4));
    InMux I__458 (
            .O(N__3008),
            .I(un5_visibley_cry_3));
    InMux I__457 (
            .O(N__3005),
            .I(N__2999));
    InMux I__456 (
            .O(N__3004),
            .I(N__2996));
    CascadeMux I__455 (
            .O(N__3003),
            .I(N__2992));
    InMux I__454 (
            .O(N__3002),
            .I(N__2989));
    LocalMux I__453 (
            .O(N__2999),
            .I(N__2986));
    LocalMux I__452 (
            .O(N__2996),
            .I(N__2983));
    InMux I__451 (
            .O(N__2995),
            .I(N__2980));
    InMux I__450 (
            .O(N__2992),
            .I(N__2977));
    LocalMux I__449 (
            .O(N__2989),
            .I(beamYZ0Z_5));
    Odrv4 I__448 (
            .O(N__2986),
            .I(beamYZ0Z_5));
    Odrv4 I__447 (
            .O(N__2983),
            .I(beamYZ0Z_5));
    LocalMux I__446 (
            .O(N__2980),
            .I(beamYZ0Z_5));
    LocalMux I__445 (
            .O(N__2977),
            .I(beamYZ0Z_5));
    InMux I__444 (
            .O(N__2966),
            .I(un5_visibley_cry_4));
    InMux I__443 (
            .O(N__2963),
            .I(N__2958));
    InMux I__442 (
            .O(N__2962),
            .I(N__2955));
    InMux I__441 (
            .O(N__2961),
            .I(N__2950));
    LocalMux I__440 (
            .O(N__2958),
            .I(N__2945));
    LocalMux I__439 (
            .O(N__2955),
            .I(N__2945));
    CascadeMux I__438 (
            .O(N__2954),
            .I(N__2942));
    InMux I__437 (
            .O(N__2953),
            .I(N__2939));
    LocalMux I__436 (
            .O(N__2950),
            .I(N__2936));
    Span4Mux_h I__435 (
            .O(N__2945),
            .I(N__2933));
    InMux I__434 (
            .O(N__2942),
            .I(N__2930));
    LocalMux I__433 (
            .O(N__2939),
            .I(beamYZ0Z_6));
    Odrv4 I__432 (
            .O(N__2936),
            .I(beamYZ0Z_6));
    Odrv4 I__431 (
            .O(N__2933),
            .I(beamYZ0Z_6));
    LocalMux I__430 (
            .O(N__2930),
            .I(beamYZ0Z_6));
    InMux I__429 (
            .O(N__2921),
            .I(un5_visibley_cry_5));
    InMux I__428 (
            .O(N__2918),
            .I(N__2912));
    InMux I__427 (
            .O(N__2917),
            .I(N__2909));
    CascadeMux I__426 (
            .O(N__2916),
            .I(N__2906));
    InMux I__425 (
            .O(N__2915),
            .I(N__2903));
    LocalMux I__424 (
            .O(N__2912),
            .I(N__2898));
    LocalMux I__423 (
            .O(N__2909),
            .I(N__2898));
    InMux I__422 (
            .O(N__2906),
            .I(N__2895));
    LocalMux I__421 (
            .O(N__2903),
            .I(beamYZ0Z_7));
    Odrv4 I__420 (
            .O(N__2898),
            .I(beamYZ0Z_7));
    LocalMux I__419 (
            .O(N__2895),
            .I(beamYZ0Z_7));
    InMux I__418 (
            .O(N__2888),
            .I(un5_visibley_cry_6));
    InMux I__417 (
            .O(N__2885),
            .I(N__2878));
    InMux I__416 (
            .O(N__2884),
            .I(N__2873));
    InMux I__415 (
            .O(N__2883),
            .I(N__2873));
    CascadeMux I__414 (
            .O(N__2882),
            .I(N__2870));
    InMux I__413 (
            .O(N__2881),
            .I(N__2867));
    LocalMux I__412 (
            .O(N__2878),
            .I(N__2862));
    LocalMux I__411 (
            .O(N__2873),
            .I(N__2862));
    InMux I__410 (
            .O(N__2870),
            .I(N__2859));
    LocalMux I__409 (
            .O(N__2867),
            .I(beamYZ0Z_8));
    Odrv4 I__408 (
            .O(N__2862),
            .I(beamYZ0Z_8));
    LocalMux I__407 (
            .O(N__2859),
            .I(beamYZ0Z_8));
    InMux I__406 (
            .O(N__2852),
            .I(bfn_8_8_0_));
    InMux I__405 (
            .O(N__2849),
            .I(N__2843));
    InMux I__404 (
            .O(N__2848),
            .I(N__2840));
    InMux I__403 (
            .O(N__2847),
            .I(N__2837));
    InMux I__402 (
            .O(N__2846),
            .I(N__2833));
    LocalMux I__401 (
            .O(N__2843),
            .I(N__2828));
    LocalMux I__400 (
            .O(N__2840),
            .I(N__2828));
    LocalMux I__399 (
            .O(N__2837),
            .I(N__2825));
    InMux I__398 (
            .O(N__2836),
            .I(N__2822));
    LocalMux I__397 (
            .O(N__2833),
            .I(beamYZ0Z_9));
    Odrv4 I__396 (
            .O(N__2828),
            .I(beamYZ0Z_9));
    Odrv4 I__395 (
            .O(N__2825),
            .I(beamYZ0Z_9));
    LocalMux I__394 (
            .O(N__2822),
            .I(beamYZ0Z_9));
    InMux I__393 (
            .O(N__2813),
            .I(un5_visibley_cry_8));
    InMux I__392 (
            .O(N__2810),
            .I(N__2807));
    LocalMux I__391 (
            .O(N__2807),
            .I(un1_beamylto9_0_a2_1));
    CascadeMux I__390 (
            .O(N__2804),
            .I(Pixel_0_sqmuxa_i_4_cascade_));
    InMux I__389 (
            .O(N__2801),
            .I(N__2798));
    LocalMux I__388 (
            .O(N__2798),
            .I(N_99));
    InMux I__387 (
            .O(N__2795),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0));
    InMux I__386 (
            .O(N__2792),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0));
    InMux I__385 (
            .O(N__2789),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0));
    CascadeMux I__384 (
            .O(N__2786),
            .I(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_));
    CascadeMux I__383 (
            .O(N__2783),
            .I(N__2779));
    InMux I__382 (
            .O(N__2782),
            .I(N__2774));
    InMux I__381 (
            .O(N__2779),
            .I(N__2774));
    LocalMux I__380 (
            .O(N__2774),
            .I(N_98));
    CascadeMux I__379 (
            .O(N__2771),
            .I(N__2766));
    CascadeMux I__378 (
            .O(N__2770),
            .I(N__2760));
    InMux I__377 (
            .O(N__2769),
            .I(N__2757));
    InMux I__376 (
            .O(N__2766),
            .I(N__2754));
    InMux I__375 (
            .O(N__2765),
            .I(N__2751));
    InMux I__374 (
            .O(N__2764),
            .I(N__2746));
    InMux I__373 (
            .O(N__2763),
            .I(N__2746));
    InMux I__372 (
            .O(N__2760),
            .I(N__2743));
    LocalMux I__371 (
            .O(N__2757),
            .I(beamYZ0Z_0));
    LocalMux I__370 (
            .O(N__2754),
            .I(beamYZ0Z_0));
    LocalMux I__369 (
            .O(N__2751),
            .I(beamYZ0Z_0));
    LocalMux I__368 (
            .O(N__2746),
            .I(beamYZ0Z_0));
    LocalMux I__367 (
            .O(N__2743),
            .I(beamYZ0Z_0));
    CascadeMux I__366 (
            .O(N__2732),
            .I(N__2724));
    InMux I__365 (
            .O(N__2731),
            .I(N__2721));
    InMux I__364 (
            .O(N__2730),
            .I(N__2718));
    InMux I__363 (
            .O(N__2729),
            .I(N__2713));
    InMux I__362 (
            .O(N__2728),
            .I(N__2713));
    InMux I__361 (
            .O(N__2727),
            .I(N__2710));
    InMux I__360 (
            .O(N__2724),
            .I(N__2707));
    LocalMux I__359 (
            .O(N__2721),
            .I(beamYZ0Z_1));
    LocalMux I__358 (
            .O(N__2718),
            .I(beamYZ0Z_1));
    LocalMux I__357 (
            .O(N__2713),
            .I(beamYZ0Z_1));
    LocalMux I__356 (
            .O(N__2710),
            .I(beamYZ0Z_1));
    LocalMux I__355 (
            .O(N__2707),
            .I(beamYZ0Z_1));
    InMux I__354 (
            .O(N__2696),
            .I(un5_visibley_cry_0));
    InMux I__353 (
            .O(N__2693),
            .I(N__2687));
    InMux I__352 (
            .O(N__2692),
            .I(N__2682));
    InMux I__351 (
            .O(N__2691),
            .I(N__2682));
    InMux I__350 (
            .O(N__2690),
            .I(N__2679));
    LocalMux I__349 (
            .O(N__2687),
            .I(beamXZ0Z_7));
    LocalMux I__348 (
            .O(N__2682),
            .I(beamXZ0Z_7));
    LocalMux I__347 (
            .O(N__2679),
            .I(beamXZ0Z_7));
    InMux I__346 (
            .O(N__2672),
            .I(N__2666));
    InMux I__345 (
            .O(N__2671),
            .I(N__2663));
    InMux I__344 (
            .O(N__2670),
            .I(N__2660));
    InMux I__343 (
            .O(N__2669),
            .I(N__2657));
    LocalMux I__342 (
            .O(N__2666),
            .I(beamXZ0Z_8));
    LocalMux I__341 (
            .O(N__2663),
            .I(beamXZ0Z_8));
    LocalMux I__340 (
            .O(N__2660),
            .I(beamXZ0Z_8));
    LocalMux I__339 (
            .O(N__2657),
            .I(beamXZ0Z_8));
    InMux I__338 (
            .O(N__2648),
            .I(N__2641));
    InMux I__337 (
            .O(N__2647),
            .I(N__2632));
    InMux I__336 (
            .O(N__2646),
            .I(N__2632));
    InMux I__335 (
            .O(N__2645),
            .I(N__2632));
    InMux I__334 (
            .O(N__2644),
            .I(N__2632));
    LocalMux I__333 (
            .O(N__2641),
            .I(N__2629));
    LocalMux I__332 (
            .O(N__2632),
            .I(beamXZ0Z_9));
    Odrv4 I__331 (
            .O(N__2629),
            .I(beamXZ0Z_9));
    CascadeMux I__330 (
            .O(N__2624),
            .I(Pixel_0_sqmuxa_i_2_1_cascade_));
    CascadeMux I__329 (
            .O(N__2621),
            .I(un1_beamylto9_0_a2_1_cascade_));
    IoInMux I__328 (
            .O(N__2618),
            .I(N__2615));
    LocalMux I__327 (
            .O(N__2615),
            .I(N__2612));
    IoSpan4Mux I__326 (
            .O(N__2612),
            .I(N__2609));
    Span4Mux_s1_v I__325 (
            .O(N__2609),
            .I(N__2605));
    IoInMux I__324 (
            .O(N__2608),
            .I(N__2602));
    Sp12to4 I__323 (
            .O(N__2605),
            .I(N__2599));
    LocalMux I__322 (
            .O(N__2602),
            .I(N__2596));
    Odrv12 I__321 (
            .O(N__2599),
            .I(VSync_c));
    Odrv12 I__320 (
            .O(N__2596),
            .I(VSync_c));
    CascadeMux I__319 (
            .O(N__2591),
            .I(N_84_cascade_));
    InMux I__318 (
            .O(N__2588),
            .I(N__2584));
    InMux I__317 (
            .O(N__2587),
            .I(N__2581));
    LocalMux I__316 (
            .O(N__2584),
            .I(N_132));
    LocalMux I__315 (
            .O(N__2581),
            .I(N_132));
    InMux I__314 (
            .O(N__2576),
            .I(N__2573));
    LocalMux I__313 (
            .O(N__2573),
            .I(Pixel_0_sqmuxa_i_2));
    CascadeMux I__312 (
            .O(N__2570),
            .I(N_101_cascade_));
    InMux I__311 (
            .O(N__2567),
            .I(N__2564));
    LocalMux I__310 (
            .O(N__2564),
            .I(Pixel_0_sqmuxa_i_1));
    InMux I__309 (
            .O(N__2561),
            .I(un8_beamx_cry_5));
    InMux I__308 (
            .O(N__2558),
            .I(un8_beamx_cry_6));
    InMux I__307 (
            .O(N__2555),
            .I(un8_beamx_cry_7));
    InMux I__306 (
            .O(N__2552),
            .I(bfn_8_4_0_));
    InMux I__305 (
            .O(N__2549),
            .I(un8_beamx_cry_9));
    CascadeMux I__304 (
            .O(N__2546),
            .I(N__2542));
    InMux I__303 (
            .O(N__2545),
            .I(N__2539));
    InMux I__302 (
            .O(N__2542),
            .I(N__2536));
    LocalMux I__301 (
            .O(N__2539),
            .I(beamXZ0Z_2));
    LocalMux I__300 (
            .O(N__2536),
            .I(beamXZ0Z_2));
    CascadeMux I__299 (
            .O(N__2531),
            .I(N__2528));
    InMux I__298 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__297 (
            .O(N__2525),
            .I(N__2520));
    InMux I__296 (
            .O(N__2524),
            .I(N__2515));
    InMux I__295 (
            .O(N__2523),
            .I(N__2515));
    Odrv4 I__294 (
            .O(N__2520),
            .I(beamXZ0Z_1));
    LocalMux I__293 (
            .O(N__2515),
            .I(beamXZ0Z_1));
    InMux I__292 (
            .O(N__2510),
            .I(N__2504));
    InMux I__291 (
            .O(N__2509),
            .I(N__2497));
    InMux I__290 (
            .O(N__2508),
            .I(N__2497));
    InMux I__289 (
            .O(N__2507),
            .I(N__2497));
    LocalMux I__288 (
            .O(N__2504),
            .I(beamXZ0Z_0));
    LocalMux I__287 (
            .O(N__2497),
            .I(beamXZ0Z_0));
    InMux I__286 (
            .O(N__2492),
            .I(un5_visiblex_cry_5));
    InMux I__285 (
            .O(N__2489),
            .I(un5_visiblex_cry_6));
    InMux I__284 (
            .O(N__2486),
            .I(N__2482));
    InMux I__283 (
            .O(N__2485),
            .I(N__2479));
    LocalMux I__282 (
            .O(N__2482),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum));
    LocalMux I__281 (
            .O(N__2479),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum));
    InMux I__280 (
            .O(N__2474),
            .I(un5_visiblex_cry_7));
    InMux I__279 (
            .O(N__2471),
            .I(un5_visiblex_cry_8));
    InMux I__278 (
            .O(N__2468),
            .I(N__2462));
    InMux I__277 (
            .O(N__2467),
            .I(N__2462));
    LocalMux I__276 (
            .O(N__2462),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum));
    InMux I__275 (
            .O(N__2459),
            .I(un8_beamx_cry_1));
    InMux I__274 (
            .O(N__2456),
            .I(un8_beamx_cry_2));
    InMux I__273 (
            .O(N__2453),
            .I(un8_beamx_cry_3));
    InMux I__272 (
            .O(N__2450),
            .I(un8_beamx_cry_4));
    InMux I__271 (
            .O(N__2447),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__270 (
            .O(N__2444),
            .I(N__2440));
    InMux I__269 (
            .O(N__2443),
            .I(N__2437));
    LocalMux I__268 (
            .O(N__2440),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23));
    LocalMux I__267 (
            .O(N__2437),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23));
    CascadeMux I__266 (
            .O(N__2432),
            .I(N__2429));
    InMux I__265 (
            .O(N__2429),
            .I(N__2426));
    LocalMux I__264 (
            .O(N__2426),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365));
    InMux I__263 (
            .O(N__2423),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__262 (
            .O(N__2420),
            .I(N__2414));
    InMux I__261 (
            .O(N__2419),
            .I(N__2414));
    LocalMux I__260 (
            .O(N__2414),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__259 (
            .O(N__2411),
            .I(N__2408));
    InMux I__258 (
            .O(N__2408),
            .I(N__2405));
    LocalMux I__257 (
            .O(N__2405),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3));
    InMux I__256 (
            .O(N__2402),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__255 (
            .O(N__2399),
            .I(N__2396));
    LocalMux I__254 (
            .O(N__2396),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__253 (
            .O(N__2393),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__252 (
            .O(N__2390),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_));
    CascadeMux I__251 (
            .O(N__2387),
            .I(N__2384));
    InMux I__250 (
            .O(N__2384),
            .I(N__2381));
    LocalMux I__249 (
            .O(N__2381),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_i));
    InMux I__248 (
            .O(N__2378),
            .I(un5_visiblex_cry_4));
    InMux I__247 (
            .O(N__2375),
            .I(un21_beamy_cry_1));
    InMux I__246 (
            .O(N__2372),
            .I(un21_beamy_cry_2));
    InMux I__245 (
            .O(N__2369),
            .I(un21_beamy_cry_3));
    InMux I__244 (
            .O(N__2366),
            .I(un21_beamy_cry_4));
    InMux I__243 (
            .O(N__2363),
            .I(un21_beamy_cry_5));
    InMux I__242 (
            .O(N__2360),
            .I(un21_beamy_cry_6));
    InMux I__241 (
            .O(N__2357),
            .I(un21_beamy_cry_7));
    InMux I__240 (
            .O(N__2354),
            .I(N__2350));
    InMux I__239 (
            .O(N__2353),
            .I(N__2343));
    LocalMux I__238 (
            .O(N__2350),
            .I(N__2340));
    InMux I__237 (
            .O(N__2349),
            .I(N__2335));
    InMux I__236 (
            .O(N__2348),
            .I(N__2335));
    InMux I__235 (
            .O(N__2347),
            .I(N__2330));
    InMux I__234 (
            .O(N__2346),
            .I(N__2330));
    LocalMux I__233 (
            .O(N__2343),
            .I(N__2327));
    Span4Mux_h I__232 (
            .O(N__2340),
            .I(N__2322));
    LocalMux I__231 (
            .O(N__2335),
            .I(N__2322));
    LocalMux I__230 (
            .O(N__2330),
            .I(un5_beamx));
    Odrv4 I__229 (
            .O(N__2327),
            .I(un5_beamx));
    Odrv4 I__228 (
            .O(N__2322),
            .I(un5_beamx));
    InMux I__227 (
            .O(N__2315),
            .I(bfn_7_8_0_));
    CascadeMux I__226 (
            .O(N__2312),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_));
    InMux I__225 (
            .O(N__2309),
            .I(N__2306));
    LocalMux I__224 (
            .O(N__2306),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0));
    InMux I__223 (
            .O(N__2303),
            .I(N__2300));
    LocalMux I__222 (
            .O(N__2300),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_i));
    CascadeMux I__221 (
            .O(N__2297),
            .I(un5_beamx_0_a2_3_cascade_));
    CascadeMux I__220 (
            .O(N__2294),
            .I(un5_beamx_0_a2_5_cascade_));
    InMux I__219 (
            .O(N__2291),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__218 (
            .O(N__2288),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__217 (
            .O(N__2285),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__216 (
            .O(N__2282),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7));
    CascadeMux I__215 (
            .O(N__2279),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_));
    CascadeMux I__214 (
            .O(N__2276),
            .I(N__2273));
    InMux I__213 (
            .O(N__2273),
            .I(N__2270));
    LocalMux I__212 (
            .O(N__2270),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0));
    InMux I__211 (
            .O(N__2267),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__210 (
            .O(N__2264),
            .I(N__2255));
    InMux I__209 (
            .O(N__2263),
            .I(N__2255));
    InMux I__208 (
            .O(N__2262),
            .I(N__2255));
    LocalMux I__207 (
            .O(N__2255),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    IoInMux I__206 (
            .O(N__2252),
            .I(N__2249));
    LocalMux I__205 (
            .O(N__2249),
            .I(N__2246));
    Span4Mux_s1_h I__204 (
            .O(N__2246),
            .I(N__2243));
    Span4Mux_h I__203 (
            .O(N__2243),
            .I(N__2240));
    Sp12to4 I__202 (
            .O(N__2240),
            .I(N__2237));
    Odrv12 I__201 (
            .O(N__2237),
            .I(\Clock50MHz.PixelClock ));
    IoInMux I__200 (
            .O(N__2234),
            .I(N__2231));
    LocalMux I__199 (
            .O(N__2231),
            .I(N__2228));
    IoSpan4Mux I__198 (
            .O(N__2228),
            .I(N__2225));
    Odrv4 I__197 (
            .O(N__2225),
            .I(Clock12MHz_c));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(un5_visibley_cry_7),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_7_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_1_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__2252),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_1_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_1_0 (
            .in0(_gnd_net_),
            .in1(N__2485),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_1_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_7_1_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_7_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_7_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_7_1_1 (
            .in0(_gnd_net_),
            .in1(N__2303),
            .in2(_gnd_net_),
            .in3(N__2291),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPF3_LC_7_1_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPF3_LC_7_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPF3_LC_7_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPF3_LC_7_1_2 (
            .in0(_gnd_net_),
            .in1(N__2309),
            .in2(N__4052),
            .in3(N__2288),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_c_RNIBRH7_LC_7_1_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_c_RNIBRH7_LC_7_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_c_RNIBRH7_LC_7_1_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_c_RNIBRH7_LC_7_1_3 (
            .in0(N__2443),
            .in1(N__2264),
            .in2(N__2276),
            .in3(N__2285),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_7_1_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_7_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_7_1_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_7_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2282),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23),
            .ltout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_7_1_5.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_7_1_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2279),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3U_LC_7_1_7.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3U_LC_7_1_7.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3U_LC_7_1_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3U_LC_7_1_7 (
            .in0(_gnd_net_),
            .in1(N__2262),
            .in2(_gnd_net_),
            .in3(N__2263),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_LC_7_2_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_LC_7_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_LC_7_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(N__2467),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_2_1.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2267),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1F_LC_7_2_2.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1F_LC_7_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1F_LC_7_2_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1F_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2312),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_2_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_2_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_2_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_7_2_7 (
            .in0(N__2468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIS9H2_9_LC_7_5_0.C_ON=1'b0;
    defparam beamY_RNIS9H2_9_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIS9H2_9_LC_7_5_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 beamY_RNIS9H2_9_LC_7_5_0 (
            .in0(N__2847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2917),
            .lcout(N_132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2T15_1_LC_7_5_3.C_ON=1'b0;
    defparam beamY_RNI2T15_1_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI2T15_1_LC_7_5_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 beamY_RNI2T15_1_LC_7_5_3 (
            .in0(N__3096),
            .in1(N__3133),
            .in2(N__3050),
            .in3(N__2730),
            .lcout(),
            .ltout(un5_beamx_0_a2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP1J7_5_LC_7_5_4.C_ON=1'b0;
    defparam beamY_RNIP1J7_5_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIP1J7_5_LC_7_5_4.LUT_INIT=16'b0000000000110000;
    LogicCell40 beamY_RNIP1J7_5_LC_7_5_4 (
            .in0(_gnd_net_),
            .in1(N__2963),
            .in2(N__2297),
            .in3(N__3004),
            .lcout(),
            .ltout(un5_beamx_0_a2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_0_LC_7_5_5.C_ON=1'b0;
    defparam beamY_RNI9DLC_0_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_0_LC_7_5_5.LUT_INIT=16'b0000000001000000;
    LogicCell40 beamY_RNI9DLC_0_LC_7_5_5 (
            .in0(N__2885),
            .in1(N__2588),
            .in2(N__2294),
            .in3(N__2765),
            .lcout(un5_beamx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_5_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_5_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_7_6_3.C_ON=1'b0;
    defparam beamY_1_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_7_6_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_1_LC_7_6_3 (
            .in0(N__2347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4272),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4179),
            .ce(N__3548),
            .sr(_gnd_net_));
    defparam beamY_0_LC_7_6_6.C_ON=1'b0;
    defparam beamY_0_LC_7_6_6.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_7_6_6.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_0_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(N__2346),
            .in2(_gnd_net_),
            .in3(N__2769),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4179),
            .ce(N__3548),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_7_7_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_7_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__2731),
            .in2(N__2771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_7_7_1.C_ON=1'b1;
    defparam beamY_2_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_7_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_2_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__3131),
            .in2(_gnd_net_),
            .in3(N__2375),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_3_LC_7_7_2.C_ON=1'b1;
    defparam beamY_3_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_7_7_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_3_LC_7_7_2 (
            .in0(N__2348),
            .in1(N__3088),
            .in2(_gnd_net_),
            .in3(N__2372),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_4_LC_7_7_3.C_ON=1'b1;
    defparam beamY_4_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_7_7_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_4_LC_7_7_3 (
            .in0(N__2354),
            .in1(N__3044),
            .in2(_gnd_net_),
            .in3(N__2369),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_5_LC_7_7_4.C_ON=1'b1;
    defparam beamY_5_LC_7_7_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_7_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__3002),
            .in2(_gnd_net_),
            .in3(N__2366),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_6_LC_7_7_5.C_ON=1'b1;
    defparam beamY_6_LC_7_7_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_7_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(N__2953),
            .in2(_gnd_net_),
            .in3(N__2363),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_7_LC_7_7_6.C_ON=1'b1;
    defparam beamY_7_LC_7_7_6.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_7_7_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_7_LC_7_7_6 (
            .in0(N__2349),
            .in1(N__2915),
            .in2(_gnd_net_),
            .in3(N__2360),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_8_LC_7_7_7.C_ON=1'b1;
    defparam beamY_8_LC_7_7_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_7_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(N__2881),
            .in2(_gnd_net_),
            .in3(N__2357),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(N__4178),
            .ce(N__3543),
            .sr(_gnd_net_));
    defparam beamY_9_LC_7_8_0.C_ON=1'b0;
    defparam beamY_9_LC_7_8_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_7_8_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_7_8_0 (
            .in0(N__2846),
            .in1(N__2353),
            .in2(_gnd_net_),
            .in3(N__2315),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4177),
            .ce(N__3544),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_1_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3170),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_1_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_1_1 (
            .in0(_gnd_net_),
            .in1(N__2419),
            .in2(N__2387),
            .in3(N__2447),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_1_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_1_2 (
            .in0(_gnd_net_),
            .in1(N__2444),
            .in2(N__2432),
            .in3(N__2423),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI4PN01_LC_8_1_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI4PN01_LC_8_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI4PN01_LC_8_1_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI4PN01_LC_8_1_3 (
            .in0(N__3226),
            .in1(N__2420),
            .in2(N__2411),
            .in3(N__2402),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_LC_8_1_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_LC_8_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_LC_8_1_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_LC_8_1_4 (
            .in0(_gnd_net_),
            .in1(N__2399),
            .in2(_gnd_net_),
            .in3(N__2393),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0),
            .ltout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_0_LC_8_1_5.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_0_LC_8_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_0_LC_8_1_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_0_LC_8_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2390),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_1_6.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_1_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_1_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_8_1_6 (
            .in0(N__2486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_LC_8_2_0.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_LC_8_2_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_LC_8_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_4_c_LC_8_2_0 (
            .in0(_gnd_net_),
            .in1(N__3489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_8_2_1 (
            .in0(_gnd_net_),
            .in1(N__3421),
            .in2(_gnd_net_),
            .in3(N__2378),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_8_2_2 (
            .in0(_gnd_net_),
            .in1(N__3454),
            .in2(N__4056),
            .in3(N__2492),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_8_2_3 (
            .in0(_gnd_net_),
            .in1(N__2690),
            .in2(_gnd_net_),
            .in3(N__2489),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_8_2_4 (
            .in0(_gnd_net_),
            .in1(N__2669),
            .in2(N__4057),
            .in3(N__2474),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_7),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5 (
            .in0(_gnd_net_),
            .in1(N__2648),
            .in2(_gnd_net_),
            .in3(N__2471),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_8_3_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__2510),
            .in2(N__2531),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_8_3_1.C_ON=1'b1;
    defparam beamX_2_LC_8_3_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_8_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(N__2545),
            .in2(_gnd_net_),
            .in3(N__2459),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_8_3_2.C_ON=1'b1;
    defparam beamX_3_LC_8_3_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_8_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(N__3393),
            .in2(_gnd_net_),
            .in3(N__2456),
            .lcout(N_97),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_8_3_3.C_ON=1'b1;
    defparam beamX_4_LC_8_3_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_8_3_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_8_3_3 (
            .in0(N__3536),
            .in1(N__3496),
            .in2(_gnd_net_),
            .in3(N__2453),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_8_3_4.C_ON=1'b1;
    defparam beamX_5_LC_8_3_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_8_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_8_3_4 (
            .in0(_gnd_net_),
            .in1(N__3427),
            .in2(_gnd_net_),
            .in3(N__2450),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_8_3_5.C_ON=1'b1;
    defparam beamX_6_LC_8_3_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_8_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(N__3459),
            .in2(_gnd_net_),
            .in3(N__2561),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_8_3_6.C_ON=1'b1;
    defparam beamX_7_LC_8_3_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_8_3_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(N__2693),
            .in2(_gnd_net_),
            .in3(N__2558),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_8_3_7.C_ON=1'b1;
    defparam beamX_8_LC_8_3_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_8_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_8_3_7 (
            .in0(_gnd_net_),
            .in1(N__2672),
            .in2(_gnd_net_),
            .in3(N__2555),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__4182),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_8_4_0.C_ON=1'b1;
    defparam beamX_9_LC_8_4_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_8_4_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__2647),
            .in2(_gnd_net_),
            .in3(N__2552),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__4181),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_8_4_1.C_ON=1'b0;
    defparam beamX_10_LC_8_4_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_8_4_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_8_4_1 (
            .in0(N__3687),
            .in1(N__3523),
            .in2(_gnd_net_),
            .in3(N__2549),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4181),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNITFL_1_LC_8_4_2.C_ON=1'b0;
    defparam beamX_RNITFL_1_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam beamX_RNITFL_1_LC_8_4_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNITFL_1_LC_8_4_2 (
            .in0(N__2523),
            .in1(N__2507),
            .in2(N__2546),
            .in3(N__3458),
            .lcout(un3_beamx_i_i_a2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_8_4_3.C_ON=1'b0;
    defparam beamX_1_LC_8_4_3.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_8_4_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 beamX_1_LC_8_4_3 (
            .in0(N__2509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2524),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4181),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_8_4_4.C_ON=1'b0;
    defparam beamX_0_LC_8_4_4.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_8_4_4.LUT_INIT=16'b0001000100010001;
    LogicCell40 beamX_0_LC_8_4_4 (
            .in0(N__3524),
            .in1(N__2508),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4181),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNINLG_7_LC_8_4_5.C_ON=1'b0;
    defparam beamX_RNINLG_7_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam beamX_RNINLG_7_LC_8_4_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamX_RNINLG_7_LC_8_4_5 (
            .in0(N__2644),
            .in1(N__2670),
            .in2(_gnd_net_),
            .in3(N__2691),
            .lcout(N_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_15_LC_8_4_6.C_ON=1'b0;
    defparam Pixel_1_RNO_15_LC_8_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_15_LC_8_4_6.LUT_INIT=16'b0111111100000011;
    LogicCell40 Pixel_1_RNO_15_LC_8_4_6 (
            .in0(N__2692),
            .in1(N__2671),
            .in2(N__3461),
            .in3(N__2645),
            .lcout(),
            .ltout(Pixel_0_sqmuxa_i_2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_14_LC_8_4_7.C_ON=1'b0;
    defparam Pixel_1_RNO_14_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_14_LC_8_4_7.LUT_INIT=16'b0001101001011000;
    LogicCell40 Pixel_1_RNO_14_LC_8_4_7 (
            .in0(N__2646),
            .in1(N__3422),
            .in2(N__2624),
            .in3(N__3493),
            .lcout(Pixel_0_sqmuxa_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQUP3_9_LC_8_5_0.C_ON=1'b0;
    defparam beamY_RNIQUP3_9_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIQUP3_9_LC_8_5_0.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_RNIQUP3_9_LC_8_5_0 (
            .in0(N__2849),
            .in1(N__2884),
            .in2(_gnd_net_),
            .in3(N__2918),
            .lcout(un1_beamylto9_0_a2_1),
            .ltout(un1_beamylto9_0_a2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_8_5_1.C_ON=1'b0;
    defparam VSync_1_LC_8_5_1.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_8_5_1.LUT_INIT=16'b1110111110101111;
    LogicCell40 VSync_1_LC_8_5_1 (
            .in0(N__2782),
            .in1(N__3143),
            .in2(N__2621),
            .in3(N__2729),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4180),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_11_LC_8_5_2.C_ON=1'b0;
    defparam Pixel_1_RNO_11_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_11_LC_8_5_2.LUT_INIT=16'b0001111101011111;
    LogicCell40 Pixel_1_RNO_11_LC_8_5_2 (
            .in0(N__3141),
            .in1(N__2727),
            .in2(N__3097),
            .in3(N__2763),
            .lcout(),
            .ltout(N_84_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_8_LC_8_5_3.C_ON=1'b0;
    defparam Pixel_1_RNO_8_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_8_LC_8_5_3.LUT_INIT=16'b0001000101010001;
    LogicCell40 Pixel_1_RNO_8_LC_8_5_3 (
            .in0(N__2962),
            .in1(N__3005),
            .in2(N__2591),
            .in3(N__3049),
            .lcout(N_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_13_LC_8_5_4.C_ON=1'b0;
    defparam Pixel_1_RNO_13_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_13_LC_8_5_4.LUT_INIT=16'b1111110111110101;
    LogicCell40 Pixel_1_RNO_13_LC_8_5_4 (
            .in0(N__3705),
            .in1(N__2848),
            .in2(N__3689),
            .in3(N__2883),
            .lcout(Pixel_0_sqmuxa_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_12_LC_8_5_5.C_ON=1'b0;
    defparam Pixel_1_RNO_12_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_12_LC_8_5_5.LUT_INIT=16'b1111111011111100;
    LogicCell40 Pixel_1_RNO_12_LC_8_5_5 (
            .in0(N__2764),
            .in1(N__3142),
            .in2(N__2783),
            .in3(N__2728),
            .lcout(),
            .ltout(N_101_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_9_LC_8_5_6.C_ON=1'b0;
    defparam Pixel_1_RNO_9_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_9_LC_8_5_6.LUT_INIT=16'b1111111111101100;
    LogicCell40 Pixel_1_RNO_9_LC_8_5_6 (
            .in0(N__2587),
            .in1(N__2576),
            .in2(N__2570),
            .in3(N__2567),
            .lcout(),
            .ltout(Pixel_0_sqmuxa_i_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_3_LC_8_5_7.C_ON=1'b0;
    defparam Pixel_1_RNO_3_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_3_LC_8_5_7.LUT_INIT=16'b1111110011110000;
    LogicCell40 Pixel_1_RNO_3_LC_8_5_7 (
            .in0(_gnd_net_),
            .in1(N__2810),
            .in2(N__2804),
            .in3(N__2801),
            .lcout(Pixel_0_sqmuxa_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_LC_8_6_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__3969),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PP_LC_8_6_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PP_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PP_LC_8_6_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PP_LC_8_6_1 (
            .in0(N__3882),
            .in1(N__3971),
            .in2(_gnd_net_),
            .in3(N__2795),
            .lcout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0),
            .carryout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0_c_RNIR53K_LC_8_6_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0_c_RNIR53K_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0_c_RNIR53K_LC_8_6_2.LUT_INIT=16'b0000000001010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0_c_RNIR53K_LC_8_6_2 (
            .in0(N__3883),
            .in1(N__3970),
            .in2(_gnd_net_),
            .in3(N__2792),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_axb_6),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0),
            .carryout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_LC_8_6_3.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_LC_8_6_3.LUT_INIT=16'b0000111100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_LC_8_6_3 (
            .in0(_gnd_net_),
            .in1(N__3884),
            .in2(N__3893),
            .in3(N__2789),
            .lcout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0),
            .ltout(un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_0_LC_8_6_4.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_0_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_0_LC_8_6_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_0_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2786),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIA525_3_LC_8_6_6.C_ON=1'b0;
    defparam beamY_RNIA525_3_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIA525_3_LC_8_6_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_RNIA525_3_LC_8_6_6 (
            .in0(N__2995),
            .in1(N__3037),
            .in2(N__3098),
            .in3(N__2961),
            .lcout(N_98),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_0_c_LC_8_7_0.C_ON=1'b1;
    defparam un5_visibley_cry_0_c_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_0_c_LC_8_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visibley_cry_0_c_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(un5_visibley_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_8_7_1.C_ON=1'b1;
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_8_7_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_0_c_RNIJVSB_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2732),
            .in3(N__2696),
            .lcout(un5_visibley_cry_0_c_RNIJVSBZ0),
            .ltout(),
            .carryin(un5_visibley_cry_0),
            .carryout(un5_visibley_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_8_7_2.C_ON=1'b1;
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_8_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_1_c_RNIL2UB_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__4000),
            .in2(N__3132),
            .in3(N__3101),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visibley_cry_1),
            .carryout(un5_visibley_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_7_3.C_ON=1'b1;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_7_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_2_c_RNIN5VB_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3089),
            .in3(N__3053),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visibley_cry_2),
            .carryout(un5_visibley_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_7_4.C_ON=1'b1;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_3_c_RNIP80C_LC_8_7_4 (
            .in0(_gnd_net_),
            .in1(N__4001),
            .in2(N__3045),
            .in3(N__3008),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visibley_cry_3),
            .carryout(un5_visibley_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_7_5.C_ON=1'b1;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_7_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_4_c_RNIRB1C_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3003),
            .in3(N__2966),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visibley_cry_4),
            .carryout(un5_visibley_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_7_6.C_ON=1'b1;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_5_c_RNITE2C_LC_8_7_6 (
            .in0(_gnd_net_),
            .in1(N__4002),
            .in2(N__2954),
            .in3(N__2921),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visibley_cry_5),
            .carryout(un5_visibley_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_7_7.C_ON=1'b1;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_6_c_RNIVH3C_LC_8_7_7 (
            .in0(_gnd_net_),
            .in1(N__4031),
            .in2(N__2916),
            .in3(N__2888),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visibley_cry_6),
            .carryout(un5_visibley_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_8_0.C_ON=1'b1;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_7_c_RNI1L4C_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(N__4035),
            .in2(N__2882),
            .in3(N__2852),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(un5_visibley_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_8_1.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_8_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__2836),
            .in2(_gnd_net_),
            .in3(N__2813),
            .lcout(un1_visibley_if_generate_plus_mult1_un26_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_1_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_1_0 (
            .in0(_gnd_net_),
            .in1(N__3316),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FE21_LC_9_1_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FE21_LC_9_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FE21_LC_9_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FE21_LC_9_1_1 (
            .in0(_gnd_net_),
            .in1(N__3202),
            .in2(N__3155),
            .in3(N__3230),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQE1_LC_9_1_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQE1_LC_9_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQE1_LC_9_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQE1_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(N__3227),
            .in2(N__3215),
            .in3(N__3206),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNIAJ623_LC_9_1_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNIAJ623_LC_9_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNIAJ623_LC_9_1_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNIAJ623_LC_9_1_3 (
            .in0(N__3370),
            .in1(N__3203),
            .in2(N__3194),
            .in3(N__3185),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_LC_9_1_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_LC_9_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_LC_9_1_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_LC_9_1_4 (
            .in0(_gnd_net_),
            .in1(N__3182),
            .in2(_gnd_net_),
            .in3(N__3176),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1),
            .ltout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_0_LC_9_1_5.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_0_LC_9_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_0_LC_9_1_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_0_LC_9_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3173),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_1_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_1_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_9_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3169),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_2_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_2_0 (
            .in0(_gnd_net_),
            .in1(N__3295),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BK1_LC_9_2_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BK1_LC_9_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BK1_LC_9_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BK1_LC_9_2_1 (
            .in0(_gnd_net_),
            .in1(N__3346),
            .in2(N__3305),
            .in3(N__3146),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNK2_LC_9_2_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNK2_LC_9_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNK2_LC_9_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNK2_LC_9_2_2 (
            .in0(_gnd_net_),
            .in1(N__3371),
            .in2(N__3359),
            .in3(N__3350),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIQBD56_LC_9_2_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIQBD56_LC_9_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIQBD56_LC_9_2_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIQBD56_LC_9_2_3 (
            .in0(N__3256),
            .in1(N__3347),
            .in2(N__3338),
            .in3(N__3329),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFL843_LC_9_2_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFL843_LC_9_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFL843_LC_9_2_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFL843_LC_9_2_4 (
            .in0(_gnd_net_),
            .in1(N__3326),
            .in2(_gnd_net_),
            .in3(N__3320),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_2_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_2_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_2_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_9_2_6 (
            .in0(N__3317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_9_2_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_9_2_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_9_2_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_9_2_7 (
            .in0(N__3296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_9_3_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_9_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_9_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_9_3_0 (
            .in0(_gnd_net_),
            .in1(N__3585),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_9_3_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_9_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_9_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_9_3_1 (
            .in0(_gnd_net_),
            .in1(N__3238),
            .in2(N__3287),
            .in3(N__3278),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_7_LC_9_3_2.C_ON=1'b1;
    defparam Pixel_1_RNO_7_LC_9_3_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_7_LC_9_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_7_LC_9_3_2 (
            .in0(_gnd_net_),
            .in1(N__3275),
            .in2(N__3257),
            .in3(N__3269),
            .lcout(Pixel_1_RNOZ0Z_7),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_9_3_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_9_3_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_9_3_3 (
            .in0(_gnd_net_),
            .in1(N__3239),
            .in2(N__3266),
            .in3(N__3252),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMD6_LC_9_3_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMD6_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMD6_LC_9_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMD6_LC_9_3_4 (
            .in0(_gnd_net_),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__3599),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6),
            .ltout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_2_LC_9_3_5.C_ON=1'b0;
    defparam Pixel_1_RNO_2_LC_9_3_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_2_LC_9_3_5.LUT_INIT=16'b0100111110110000;
    LogicCell40 Pixel_1_RNO_2_LC_9_3_5 (
            .in0(N__3586),
            .in1(N__3575),
            .in2(N__3596),
            .in3(N__3593),
            .lcout(N_94),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_9_3_6.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_9_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_9_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_9_3_6 (
            .in0(N__4053),
            .in1(N__3587),
            .in2(_gnd_net_),
            .in3(N__3497),
            .lcout(un5_visiblex_i),
            .ltout(un5_visiblex_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_1_LC_9_3_7.C_ON=1'b0;
    defparam Pixel_1_RNO_1_LC_9_3_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_1_LC_9_3_7.LUT_INIT=16'b0011110101110011;
    LogicCell40 Pixel_1_RNO_1_LC_9_3_7 (
            .in0(N__3398),
            .in1(N__3574),
            .in2(N__3566),
            .in3(N__3563),
            .lcout(N_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_10_LC_9_4_1.C_ON=1'b0;
    defparam Pixel_1_RNO_10_LC_9_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_10_LC_9_4_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 Pixel_1_RNO_10_LC_9_4_1 (
            .in0(_gnd_net_),
            .in1(N__4150),
            .in2(_gnd_net_),
            .in3(N__4273),
            .lcout(G_7_0_a4_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIHUU5_10_LC_9_4_3.C_ON=1'b0;
    defparam beamX_RNIHUU5_10_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam beamX_RNIHUU5_10_LC_9_4_3.LUT_INIT=16'b0000001000000000;
    LogicCell40 beamX_RNIHUU5_10_LC_9_4_3 (
            .in0(N__3686),
            .in1(N__3423),
            .in2(N__3397),
            .in3(N__3494),
            .lcout(),
            .ltout(un3_beamx_i_i_a2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_1_LC_9_4_4.C_ON=1'b0;
    defparam beamX_RNI5457_1_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_1_LC_9_4_4.LUT_INIT=16'b0000000011000000;
    LogicCell40 beamX_RNI5457_1_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(N__3557),
            .in2(N__3551),
            .in3(N__3706),
            .lcout(beamX_RNI5457Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_RNO_0_LC_9_4_6.C_ON=1'b0;
    defparam HSync_1_RNO_0_LC_9_4_6.SEQ_MODE=4'b0000;
    defparam HSync_1_RNO_0_LC_9_4_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 HSync_1_RNO_0_LC_9_4_6 (
            .in0(N__3495),
            .in1(N__3460),
            .in2(N__3428),
            .in3(N__3392),
            .lcout(),
            .ltout(N_130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_9_4_7.C_ON=1'b0;
    defparam HSync_1_LC_9_4_7.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_9_4_7.LUT_INIT=16'b1111111111111010;
    LogicCell40 HSync_1_LC_9_4_7 (
            .in0(N__3707),
            .in1(_gnd_net_),
            .in2(N__3692),
            .in3(N__3688),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4183),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_5_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__3616),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJI2_LC_9_5_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJI2_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJI2_LC_9_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJI2_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__3753),
            .in2(N__3716),
            .in3(N__3635),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6P3_LC_9_5_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6P3_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6P3_LC_9_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6P3_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(N__3833),
            .in2(N__3758),
            .in3(N__3632),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QOR3_LC_9_5_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QOR3_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QOR3_LC_9_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QOR3_LC_9_5_3 (
            .in0(_gnd_net_),
            .in1(N__3757),
            .in2(N__3824),
            .in3(N__3629),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNIEFE58_LC_9_5_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNIEFE58_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNIEFE58_LC_9_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNIEFE58_LC_9_5_4 (
            .in0(N__4339),
            .in1(N__3812),
            .in2(N__3734),
            .in3(N__3626),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_LC_9_5_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_LC_9_5_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_LC_9_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(N__3794),
            .in2(_gnd_net_),
            .in3(N__3623),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94),
            .ltout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_0_LC_9_5_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_0_LC_9_5_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_0_LC_9_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_0_LC_9_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3620),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_7 (
            .in0(N__3617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_9_6_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_9_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(N__3724),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVF1_LC_9_6_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVF1_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVF1_LC_9_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVF1_LC_9_6_1 (
            .in0(_gnd_net_),
            .in1(N__3839),
            .in2(N__3783),
            .in3(N__3827),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GI1_LC_9_6_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GI1_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GI1_LC_9_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GI1_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(N__3776),
            .in2(N__4088),
            .in3(N__3815),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6II1_LC_9_6_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6II1_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6II1_LC_9_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6II1_LC_9_6_3 (
            .in0(_gnd_net_),
            .in1(N__4076),
            .in2(N__3784),
            .in3(N__3806),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_c_RNI9GRQ3_LC_9_6_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_c_RNI9GRQ3_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_c_RNI9GRQ3_LC_9_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_c_RNI9GRQ3_LC_9_6_4 (
            .in0(N__3752),
            .in1(N__3935),
            .in2(N__3803),
            .in3(N__3788),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_LC_9_6_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_LC_9_6_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_LC_9_6_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_LC_9_6_5 (
            .in0(N__3922),
            .in1(N__3908),
            .in2(N__3785),
            .in3(N__3761),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1),
            .ltout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_0_LC_9_6_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_0_LC_9_6_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_0_LC_9_6_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_0_LC_9_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3737),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_6_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_6_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_6_7 (
            .in0(N__3725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_9_7_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_9_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_9_7_0 (
            .in0(_gnd_net_),
            .in1(N__3847),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_9_7_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_9_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(N__4036),
            .in2(N__3857),
            .in3(N__4079),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_9_7_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_9_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(N__3873),
            .in2(N__4054),
            .in3(N__4070),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULV_LC_9_7_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULV_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULV_LC_9_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULV_LC_9_7_3 (
            .in0(_gnd_net_),
            .in1(N__4067),
            .in2(N__4055),
            .in3(N__3926),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_9_7_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_9_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3923),
            .in3(N__3899),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_9_7_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_9_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3896),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_9_7_6.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_9_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_0_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3872),
            .lcout(un5_visibley_cry_8_c_RNI3O5CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_sbtinv_LC_9_7_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_sbtinv_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_sbtinv_LC_9_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_sbtinv_LC_9_7_7 (
            .in0(N__3848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_4_LC_11_3_0.C_ON=1'b0;
    defparam Pixel_1_RNO_4_LC_11_3_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_4_LC_11_3_0.LUT_INIT=16'b1110111111111111;
    LogicCell40 Pixel_1_RNO_4_LC_11_3_0 (
            .in0(N__4417),
            .in1(N__4402),
            .in2(N__4154),
            .in3(N__4094),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_0_LC_11_3_1.C_ON=1'b0;
    defparam Pixel_1_RNO_0_LC_11_3_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_0_LC_11_3_1.LUT_INIT=16'b1111111111001011;
    LogicCell40 Pixel_1_RNO_0_LC_11_3_1 (
            .in0(N__4277),
            .in1(N__4115),
            .in2(N__4253),
            .in3(N__4391),
            .lcout(),
            .ltout(N_49_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_11_3_2.C_ON=1'b0;
    defparam Pixel_1_LC_11_3_2.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_11_3_2.LUT_INIT=16'b0001010000000101;
    LogicCell40 Pixel_1_LC_11_3_2 (
            .in0(N__4250),
            .in1(N__4238),
            .in2(N__4229),
            .in3(N__4226),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4184),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_4_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_4_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_4_0 (
            .in0(_gnd_net_),
            .in1(N__4149),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTP21_LC_11_4_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTP21_LC_11_4_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTP21_LC_11_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTP21_LC_11_4_1 (
            .in0(_gnd_net_),
            .in1(N__4385),
            .in2(N__4462),
            .in3(N__4121),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78K1_LC_11_4_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78K1_LC_11_4_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78K1_LC_11_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78K1_LC_11_4_2 (
            .in0(_gnd_net_),
            .in1(N__4457),
            .in2(N__4508),
            .in3(N__4118),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_6_LC_11_4_3.C_ON=1'b1;
    defparam Pixel_1_RNO_6_LC_11_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_6_LC_11_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_6_LC_11_4_3 (
            .in0(_gnd_net_),
            .in1(N__4496),
            .in2(N__4463),
            .in3(N__4109),
            .lcout(Pixel_1_RNOZ0Z_6),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_4_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_4_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_4_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_4_4 (
            .in0(_gnd_net_),
            .in1(N__4487),
            .in2(N__4106),
            .in3(N__4453),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMI32_LC_11_4_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMI32_LC_11_4_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMI32_LC_11_4_5.LUT_INIT=16'b0000111111110000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMI32_LC_11_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4478),
            .in3(N__4097),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32),
            .ltout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_5_LC_11_4_6.C_ON=1'b0;
    defparam Pixel_1_RNO_5_LC_11_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_5_LC_11_4_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_5_LC_11_4_6 (
            .in0(N__4427),
            .in1(N__4418),
            .in2(N__4406),
            .in3(N__4403),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_4_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_4_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4526),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_5_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(N__4540),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TM4_LC_11_5_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TM4_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TM4_LC_11_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TM4_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__4347),
            .in2(N__4379),
            .in3(N__4367),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICA117_LC_11_5_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICA117_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICA117_LC_11_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICA117_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__4364),
            .in2(N__4352),
            .in3(N__4355),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIIL78_LC_11_5_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIIL78_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIIL78_LC_11_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIIL78_LC_11_5_3 (
            .in0(_gnd_net_),
            .in1(N__4351),
            .in2(N__4328),
            .in3(N__4316),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIA6LKG_LC_11_5_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIA6LKG_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIA6LKG_LC_11_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIA6LKG_LC_11_5_4 (
            .in0(N__4643),
            .in1(N__4313),
            .in2(N__4304),
            .in3(N__4292),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_LC_11_5_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_LC_11_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_LC_11_5_5 (
            .in0(_gnd_net_),
            .in1(N__4289),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8),
            .ltout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_0_LC_11_5_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_0_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_0_LC_11_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_0_LC_11_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4544),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_5_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_5_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_5_7 (
            .in0(N__4541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(N__4525),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPH_LC_12_4_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPH_LC_12_4_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPH_LC_12_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPH_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__4572),
            .in2(N__4436),
            .in3(N__4499),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85Q_LC_12_4_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85Q_LC_12_4_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85Q_LC_12_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85Q_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(N__4676),
            .in2(N__4577),
            .in3(N__4490),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPU_LC_12_4_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPU_LC_12_4_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPU_LC_12_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPU_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(N__4576),
            .in2(N__4661),
            .in3(N__4481),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIKSOE32_LC_12_4_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIKSOE32_LC_12_4_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIKSOE32_LC_12_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIKSOE32_LC_12_4_4 (
            .in0(N__4461),
            .in1(N__4619),
            .in2(N__4553),
            .in3(N__4469),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNA21_LC_12_4_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNA21_LC_12_4_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNA21_LC_12_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNA21_LC_12_4_5 (
            .in0(_gnd_net_),
            .in1(N__4595),
            .in2(_gnd_net_),
            .in3(N__4466),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4709),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_5_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_5_0 (
            .in0(_gnd_net_),
            .in1(N__4708),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQN8_LC_12_5_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQN8_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQN8_LC_12_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQN8_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(N__4644),
            .in2(N__4685),
            .in3(N__4670),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCD_LC_12_5_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCD_LC_12_5_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCD_LC_12_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCD_LC_12_5_2 (
            .in0(_gnd_net_),
            .in1(N__4667),
            .in2(N__4649),
            .in3(N__4652),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMF_LC_12_5_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMF_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMF_LC_12_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMF_LC_12_5_3 (
            .in0(_gnd_net_),
            .in1(N__4648),
            .in2(N__4628),
            .in3(N__4613),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGF1T11_LC_12_5_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGF1T11_LC_12_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGF1T11_LC_12_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGF1T11_LC_12_5_4 (
            .in0(N__4571),
            .in1(N__4610),
            .in2(N__4604),
            .in3(N__4589),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_LC_12_5_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_LC_12_5_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_LC_12_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_LC_12_5_5 (
            .in0(_gnd_net_),
            .in1(N__4586),
            .in2(_gnd_net_),
            .in3(N__4580),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0),
            .ltout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_0_LC_12_5_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_0_LC_12_5_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_0_LC_12_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_0_LC_12_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4556),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
