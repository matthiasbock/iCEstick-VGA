PixelClock_inst: PixelClock
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
