-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 16:21:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic;
    Clock12MHz : in std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_1_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_i_0 : std_logic;
signal un13_x_i_i_a2_1 : std_logic;
signal \N_130_cascade_\ : std_logic;
signal \y_RNIA5P7Z0Z_9\ : std_logic;
signal \un13_x_i_i_a2_0_3_cascade_\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \Counter_cry_0\ : std_logic;
signal \Counter_cry_1\ : std_logic;
signal \Counter_cry_2\ : std_logic;
signal \Counter_cry_3\ : std_logic;
signal \Counter_cry_4\ : std_logic;
signal \Counter_cry_5\ : std_logic;
signal \Counter_cry_6\ : std_logic;
signal \Counter_cry_7\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \Counter_cry_8\ : std_logic;
signal \Counter_cry_9\ : std_logic;
signal \Counter_cry_10\ : std_logic;
signal \Counter_cry_11\ : std_logic;
signal \Counter_cry_12\ : std_logic;
signal \ClockVGAZ0\ : std_logic;
signal \Clock12MHz_c_g\ : std_logic;
signal \G_167\ : std_logic;
signal \bfn_2_1_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\ : std_logic;
signal un2_y_if_generate_plus_mult1_un26_sum_cry_5 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_i_7 : std_logic;
signal \N_140\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \yZ0Z_0\ : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \un3_y_cry_1_THRU_CO\ : std_logic;
signal un3_y_cry_1 : std_logic;
signal \yZ0Z_3\ : std_logic;
signal \un3_y_cry_2_THRU_CO\ : std_logic;
signal un3_y_cry_2 : std_logic;
signal \yZ0Z_4\ : std_logic;
signal un3_y_cry_3 : std_logic;
signal \yZ0Z_5\ : std_logic;
signal un3_y_cry_4 : std_logic;
signal \yZ0Z_6\ : std_logic;
signal un3_y_cry_5 : std_logic;
signal \yZ0Z_7\ : std_logic;
signal un3_y_cry_6 : std_logic;
signal \yZ0Z_8\ : std_logic;
signal un3_y_cry_7 : std_logic;
signal un3_y_cry_8 : std_logic;
signal \N_130\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \yZ0Z_9\ : std_logic;
signal \CounterZ0Z_7\ : std_logic;
signal \CounterZ0Z_6\ : std_logic;
signal \CounterZ0Z_8\ : std_logic;
signal \CounterZ0Z_13\ : std_logic;
signal \CounterZ0Z_12\ : std_logic;
signal \un2_counterlt11_cascade_\ : std_logic;
signal un2_counter_0 : std_logic;
signal \CounterZ0Z_4\ : std_logic;
signal \CounterZ0Z_0\ : std_logic;
signal \CounterZ0Z_3\ : std_logic;
signal \CounterZ0Z_2\ : std_logic;
signal \CounterZ0Z_1\ : std_logic;
signal \CounterZ0Z_5\ : std_logic;
signal un2_counterlto4_2 : std_logic;
signal un2_counterlt7 : std_logic;
signal \CounterZ0Z_11\ : std_logic;
signal \CounterZ0Z_9\ : std_logic;
signal \CounterZ0Z_10\ : std_logic;
signal un2_counterlto11_1 : std_logic;
signal \N_83_cascade_\ : std_logic;
signal \N_85\ : std_logic;
signal \un13lto4_i_1_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET_cascade_\ : std_logic;
signal \yZ0Z_2\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_i_0 : std_logic;
signal \bfn_5_1_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO\ : std_logic;
signal un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO\ : std_logic;
signal un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3 : std_logic;
signal \Pixel_RNOZ0Z_4\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1\ : std_logic;
signal \N_49\ : std_logic;
signal un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4 : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \xZ0Z_0\ : std_logic;
signal \xZ0Z_1\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \xZ0Z_2\ : std_logic;
signal un16_x_cry_1 : std_logic;
signal \N_89\ : std_logic;
signal un16_x_cry_2 : std_logic;
signal un16_x_cry_3 : std_logic;
signal un16_x_cry_4 : std_logic;
signal un16_x_cry_5 : std_logic;
signal un16_x_cry_6 : std_logic;
signal un16_x_cry_7 : std_logic;
signal un16_x_cry_8 : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \bfn_6_1_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4 : std_logic;
signal \Pixel_RNOZ0Z_6\ : std_logic;
signal un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5 : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO\ : std_logic;
signal \N_57\ : std_logic;
signal \N_59\ : std_logic;
signal \N_55\ : std_logic;
signal \N_47\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\ : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_i_0 : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_i : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \Pixel_0_sqmuxa_i_1\ : std_logic;
signal \Pixel_0_sqmuxa_i_0\ : std_logic;
signal \HSync_c\ : std_logic;
signal \N_90\ : std_logic;
signal \xZ0Z_5\ : std_logic;
signal \xZ0Z_6\ : std_logic;
signal \xZ0Z_4\ : std_logic;
signal un11_x_0_a2_2_2 : std_logic;
signal \un11_x_0_a2_1_cascade_\ : std_logic;
signal \x_RNID8R22Z0Z_9\ : std_logic;
signal \xZ0Z_9\ : std_logic;
signal un1_xlto9_i_0 : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \xZ0Z_7\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\ : std_logic;
signal \xZ0Z_8\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \y_RNIMA162Z0Z_9\ : std_logic;
signal \VSync_c\ : std_logic;
signal \ClockVGA_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \Clock12MHz_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;

begin
    \Clock12MHz_wire\ <= Clock12MHz;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;

    \Clock12MHz_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__4762\,
            GLOBALBUFFEROUTPUT => \Clock12MHz_c_g\
        );

    \Clock12MHz_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4764\,
            DIN => \N__4763\,
            DOUT => \N__4762\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4764\,
            PADOUT => \N__4763\,
            PADIN => \N__4762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4753\,
            DIN => \N__4752\,
            DOUT => \N__4751\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4753\,
            PADOUT => \N__4752\,
            PADIN => \N__4751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4744\,
            DIN => \N__4743\,
            DOUT => \N__4742\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4744\,
            PADOUT => \N__4743\,
            PADIN => \N__4742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4302\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4735\,
            DIN => \N__4734\,
            DOUT => \N__4733\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4735\,
            PADOUT => \N__4734\,
            PADIN => \N__4733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1021\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4713\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__4710\,
            I => \N__4703\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__4709\,
            I => \N__4700\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__4708\,
            I => \N__4696\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__4707\,
            I => \N__4693\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__4706\,
            I => \N__4690\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4684\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4681\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4676\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4676\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4671\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4671\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4666\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4666\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4663\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4659\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4654\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4654\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4649\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4666\,
            I => \N__4649\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4646\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4643\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__4659\,
            I => \N__4637\
        );

    \I__997\ : Span4Mux_s3_h
    port map (
            O => \N__4654\,
            I => \N__4637\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__4649\,
            I => \N__4632\
        );

    \I__995\ : Span4Mux_v
    port map (
            O => \N__4646\,
            I => \N__4632\
        );

    \I__994\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4627\
        );

    \I__993\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4627\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__4637\,
            I => \CONSTANT_ONE_NET\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__4632\,
            I => \CONSTANT_ONE_NET\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4627\,
            I => \CONSTANT_ONE_NET\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__988\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4614\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\
        );

    \I__986\ : InMux
    port map (
            O => \N__4611\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__985\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4605\,
            I => un2_x_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__983\ : InMux
    port map (
            O => \N__4602\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__982\ : InMux
    port map (
            O => \N__4599\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__981\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4592\
        );

    \I__980\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4592\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4589\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4584\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\
        );

    \I__976\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4575\
        );

    \I__975\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4575\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4575\,
            I => un2_x_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__972\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4560\
        );

    \I__971\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4560\
        );

    \I__970\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4560\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4560\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__968\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4554\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\
        );

    \I__966\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4540\
        );

    \I__965\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4540\
        );

    \I__964\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4535\
        );

    \I__963\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4535\
        );

    \I__962\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4532\
        );

    \I__961\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4529\
        );

    \I__960\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4526\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4521\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4521\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4532\,
            I => \xZ0Z_8\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4529\,
            I => \xZ0Z_8\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4526\,
            I => \xZ0Z_8\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__4521\,
            I => \xZ0Z_8\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__952\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4506\,
            I => un2_x_if_generate_plus_mult1_un47_sum_i
        );

    \I__950\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4499\
        );

    \I__949\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4496\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4491\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4496\,
            I => \N__4491\
        );

    \I__946\ : Odrv12
    port map (
            O => \N__4491\,
            I => \y_RNIMA162Z0Z_9\
        );

    \I__945\ : IoInMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__943\ : Odrv12
    port map (
            O => \N__4482\,
            I => \VSync_c\
        );

    \I__942\ : ClkMux
    port map (
            O => \N__4479\,
            I => \N__4452\
        );

    \I__941\ : ClkMux
    port map (
            O => \N__4478\,
            I => \N__4452\
        );

    \I__940\ : ClkMux
    port map (
            O => \N__4477\,
            I => \N__4452\
        );

    \I__939\ : ClkMux
    port map (
            O => \N__4476\,
            I => \N__4452\
        );

    \I__938\ : ClkMux
    port map (
            O => \N__4475\,
            I => \N__4452\
        );

    \I__937\ : ClkMux
    port map (
            O => \N__4474\,
            I => \N__4452\
        );

    \I__936\ : ClkMux
    port map (
            O => \N__4473\,
            I => \N__4452\
        );

    \I__935\ : ClkMux
    port map (
            O => \N__4472\,
            I => \N__4452\
        );

    \I__934\ : ClkMux
    port map (
            O => \N__4471\,
            I => \N__4452\
        );

    \I__933\ : GlobalMux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__932\ : gio2CtrlBuf
    port map (
            O => \N__4449\,
            I => \ClockVGA_g\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__4446\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\
        );

    \I__930\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4439\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__4442\,
            I => \N__4436\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4439\,
            I => \N__4429\
        );

    \I__927\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4426\
        );

    \I__926\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4423\
        );

    \I__925\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4418\
        );

    \I__924\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4418\
        );

    \I__923\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4415\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__4429\,
            I => \N__4412\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4426\,
            I => \xZ0Z_7\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4423\,
            I => \xZ0Z_7\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4418\,
            I => \xZ0Z_7\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4415\,
            I => \xZ0Z_7\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__4412\,
            I => \xZ0Z_7\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__915\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4395\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\
        );

    \I__913\ : InMux
    port map (
            O => \N__4392\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__911\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4383\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4383\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\
        );

    \I__909\ : InMux
    port map (
            O => \N__4380\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__908\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4374\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4374\,
            I => un2_x_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__906\ : InMux
    port map (
            O => \N__4371\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__905\ : InMux
    port map (
            O => \N__4368\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__904\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4361\
        );

    \I__903\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4358\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4361\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4358\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4353\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\
        );

    \I__899\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4344\
        );

    \I__898\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4344\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4344\,
            I => un2_x_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__896\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4338\,
            I => un2_x_if_generate_plus_mult1_un40_sum_i
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__893\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4329\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\
        );

    \I__891\ : InMux
    port map (
            O => \N__4326\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__4323\,
            I => \N__4320\
        );

    \I__889\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__4314\,
            I => \Pixel_0_sqmuxa_i_1\
        );

    \I__886\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4308\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__4305\,
            I => \Pixel_0_sqmuxa_i_0\
        );

    \I__883\ : IoInMux
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__881\ : IoSpan4Mux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__880\ : Span4Mux_s2_v
    port map (
            O => \N__4293\,
            I => \N__4290\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__4290\,
            I => \HSync_c\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__877\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N_90\
        );

    \I__875\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4270\
        );

    \I__874\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4267\
        );

    \I__873\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4264\
        );

    \I__872\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4257\
        );

    \I__871\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4257\
        );

    \I__870\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4257\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4270\,
            I => \N__4252\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4267\,
            I => \N__4252\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4264\,
            I => \xZ0Z_5\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4257\,
            I => \xZ0Z_5\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4252\,
            I => \xZ0Z_5\
        );

    \I__864\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4237\
        );

    \I__863\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4230\
        );

    \I__862\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4230\
        );

    \I__861\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4230\
        );

    \I__860\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4225\
        );

    \I__859\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4225\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4237\,
            I => \xZ0Z_6\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4230\,
            I => \xZ0Z_6\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4225\,
            I => \xZ0Z_6\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \N__4210\
        );

    \I__854\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4207\
        );

    \I__853\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4202\
        );

    \I__852\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4202\
        );

    \I__851\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4199\
        );

    \I__850\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4194\
        );

    \I__849\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4194\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4191\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4188\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4199\,
            I => \xZ0Z_4\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4194\,
            I => \xZ0Z_4\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4191\,
            I => \xZ0Z_4\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__4188\,
            I => \xZ0Z_4\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__841\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4170\
        );

    \I__840\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4170\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4170\,
            I => un11_x_0_a2_2_2
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4167\,
            I => \un11_x_0_a2_1_cascade_\
        );

    \I__837\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4151\
        );

    \I__836\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4151\
        );

    \I__835\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4144\
        );

    \I__834\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4144\
        );

    \I__833\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4144\
        );

    \I__832\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4135\
        );

    \I__831\ : InMux
    port map (
            O => \N__4158\,
            I => \N__4135\
        );

    \I__830\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4135\
        );

    \I__829\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4135\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4130\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4125\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4125\
        );

    \I__825\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4122\
        );

    \I__824\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4119\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__4130\,
            I => \N__4110\
        );

    \I__822\ : Span4Mux_v
    port map (
            O => \N__4125\,
            I => \N__4110\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4122\,
            I => \N__4110\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4119\,
            I => \N__4107\
        );

    \I__819\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4104\
        );

    \I__818\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4101\
        );

    \I__817\ : Span4Mux_h
    port map (
            O => \N__4110\,
            I => \N__4098\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__4107\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4104\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4101\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__4098\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__812\ : InMux
    port map (
            O => \N__4089\,
            I => \N__4081\
        );

    \I__811\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4072\
        );

    \I__810\ : InMux
    port map (
            O => \N__4087\,
            I => \N__4072\
        );

    \I__809\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4072\
        );

    \I__808\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4072\
        );

    \I__807\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4069\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4081\,
            I => \xZ0Z_9\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4072\,
            I => \xZ0Z_9\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4069\,
            I => \xZ0Z_9\
        );

    \I__803\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4059\,
            I => un1_xlto9_i_0
        );

    \I__801\ : InMux
    port map (
            O => \N__4056\,
            I => un2_x_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__799\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4047\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\
        );

    \I__797\ : InMux
    port map (
            O => \N__4044\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__795\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4035\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\
        );

    \I__793\ : InMux
    port map (
            O => \N__4032\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__792\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4026\,
            I => un2_x_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__790\ : InMux
    port map (
            O => \N__4023\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__789\ : InMux
    port map (
            O => \N__4020\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__788\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4013\
        );

    \I__787\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4010\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4013\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4010\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__4005\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3996\
        );

    \I__782\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3996\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3996\,
            I => un2_x_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__779\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3987\,
            I => un2_x_if_generate_plus_mult1_un61_sum_i
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__776\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3978\,
            I => un2_x_if_generate_plus_mult1_un54_sum_i
        );

    \I__774\ : InMux
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3972\,
            I => \Pixel_RNOZ0Z_6\
        );

    \I__772\ : InMux
    port map (
            O => \N__3969\,
            I => un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__770\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3957\
        );

    \I__769\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3957\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3957\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\
        );

    \I__767\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3948\
        );

    \I__766\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3948\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3948\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__763\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3939\,
            I => \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO\
        );

    \I__761\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3933\,
            I => \N_57\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__758\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3924\,
            I => \N_59\
        );

    \I__756\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3918\,
            I => \N_55\
        );

    \I__754\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3912\,
            I => \N_47\
        );

    \I__752\ : IoInMux
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__750\ : Span4Mux_s0_v
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__3900\,
            I => \Pixel_c\
        );

    \I__748\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3894\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3894\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\
        );

    \I__746\ : InMux
    port map (
            O => \N__3891\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__744\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3882\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3882\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\
        );

    \I__742\ : InMux
    port map (
            O => \N__3879\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__741\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3873\,
            I => un2_x_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__739\ : InMux
    port map (
            O => \N__3870\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__738\ : InMux
    port map (
            O => \N__3867\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__3864\,
            I => \N__3860\
        );

    \I__736\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3856\
        );

    \I__735\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3851\
        );

    \I__734\ : InMux
    port map (
            O => \N__3859\,
            I => \N__3851\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3856\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3851\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\
        );

    \I__731\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3842\
        );

    \I__730\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3839\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3842\,
            I => un2_x_if_generate_plus_mult1_un75_sum_i_0
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3839\,
            I => un2_x_if_generate_plus_mult1_un75_sum_i_0
        );

    \I__727\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3829\
        );

    \I__726\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3826\
        );

    \I__725\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3823\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3829\,
            I => \N__3820\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3826\,
            I => \N_89\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3823\,
            I => \N_89\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__3820\,
            I => \N_89\
        );

    \I__720\ : InMux
    port map (
            O => \N__3813\,
            I => un16_x_cry_2
        );

    \I__719\ : InMux
    port map (
            O => \N__3810\,
            I => un16_x_cry_3
        );

    \I__718\ : InMux
    port map (
            O => \N__3807\,
            I => un16_x_cry_4
        );

    \I__717\ : InMux
    port map (
            O => \N__3804\,
            I => un16_x_cry_5
        );

    \I__716\ : InMux
    port map (
            O => \N__3801\,
            I => un16_x_cry_6
        );

    \I__715\ : InMux
    port map (
            O => \N__3798\,
            I => un16_x_cry_7
        );

    \I__714\ : InMux
    port map (
            O => \N__3795\,
            I => \bfn_5_5_0_\
        );

    \I__713\ : InMux
    port map (
            O => \N__3792\,
            I => un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4
        );

    \I__712\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3783\
        );

    \I__711\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3783\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3783\,
            I => un2_x_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__709\ : InMux
    port map (
            O => \N__3780\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__3777\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__706\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3768\,
            I => un2_x_if_generate_plus_mult1_un68_sum_i
        );

    \I__704\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3759\
        );

    \I__703\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3752\
        );

    \I__702\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3752\
        );

    \I__701\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3752\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3759\,
            I => \xZ0Z_0\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3752\,
            I => \xZ0Z_0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3747\,
            I => \N__3744\
        );

    \I__697\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3739\
        );

    \I__696\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3734\
        );

    \I__695\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3734\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3739\,
            I => \xZ0Z_1\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3734\,
            I => \xZ0Z_1\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3729\,
            I => \N__3725\
        );

    \I__691\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3722\
        );

    \I__690\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3719\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3722\,
            I => \xZ0Z_2\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3719\,
            I => \xZ0Z_2\
        );

    \I__687\ : InMux
    port map (
            O => \N__3714\,
            I => un16_x_cry_1
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3711\,
            I => \CONSTANT_ONE_NET_cascade_\
        );

    \I__685\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3698\
        );

    \I__684\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3698\
        );

    \I__683\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3695\
        );

    \I__682\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3692\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3704\,
            I => \N__3689\
        );

    \I__680\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3685\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3682\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3695\,
            I => \N__3677\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3692\,
            I => \N__3677\
        );

    \I__676\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3674\
        );

    \I__675\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3671\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3685\,
            I => \N__3664\
        );

    \I__673\ : Span4Mux_h
    port map (
            O => \N__3682\,
            I => \N__3664\
        );

    \I__672\ : Span4Mux_s0_v
    port map (
            O => \N__3677\,
            I => \N__3664\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3674\,
            I => \yZ0Z_2\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3671\,
            I => \yZ0Z_2\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__3664\,
            I => \yZ0Z_2\
        );

    \I__668\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3653\
        );

    \I__667\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3650\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3653\,
            I => un2_y_if_generate_plus_mult1_un75_sum_i_0
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3650\,
            I => un2_y_if_generate_plus_mult1_un75_sum_i_0
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3645\,
            I => \N__3641\
        );

    \I__663\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3638\
        );

    \I__662\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3635\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3638\,
            I => \N__3630\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3635\,
            I => \N__3630\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__3630\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0\
        );

    \I__658\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3624\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3624\,
            I => \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO\
        );

    \I__656\ : InMux
    port map (
            O => \N__3621\,
            I => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2
        );

    \I__655\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3615\,
            I => \N__3611\
        );

    \I__653\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3608\
        );

    \I__652\ : Span4Mux_s0_v
    port map (
            O => \N__3611\,
            I => \N__3603\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3608\,
            I => \N__3603\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__3603\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1\
        );

    \I__649\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3597\,
            I => \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO\
        );

    \I__647\ : InMux
    port map (
            O => \N__3594\,
            I => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3
        );

    \I__646\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__3585\,
            I => \Pixel_RNOZ0Z_4\
        );

    \I__643\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3576\
        );

    \I__642\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3569\
        );

    \I__641\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3569\
        );

    \I__640\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3569\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3576\,
            I => \N__3564\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3569\,
            I => \N__3564\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__3564\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__635\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3555\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3555\,
            I => \N_49\
        );

    \I__633\ : InMux
    port map (
            O => \N__3552\,
            I => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4
        );

    \I__632\ : InMux
    port map (
            O => \N__3549\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__631\ : InMux
    port map (
            O => \N__3546\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__630\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3539\
        );

    \I__629\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3536\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3539\,
            I => \CounterZ0Z_13\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3536\,
            I => \CounterZ0Z_13\
        );

    \I__626\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3527\
        );

    \I__625\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3524\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3527\,
            I => \CounterZ0Z_12\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3524\,
            I => \CounterZ0Z_12\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3519\,
            I => \un2_counterlt11_cascade_\
        );

    \I__621\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3495\
        );

    \I__620\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3495\
        );

    \I__619\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3495\
        );

    \I__618\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3486\
        );

    \I__617\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3486\
        );

    \I__616\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3486\
        );

    \I__615\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3486\
        );

    \I__614\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3477\
        );

    \I__613\ : InMux
    port map (
            O => \N__3508\,
            I => \N__3477\
        );

    \I__612\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3477\
        );

    \I__611\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3477\
        );

    \I__610\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3468\
        );

    \I__609\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3468\
        );

    \I__608\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3468\
        );

    \I__607\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3468\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3495\,
            I => un2_counter_0
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3486\,
            I => un2_counter_0
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3477\,
            I => un2_counter_0
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3468\,
            I => un2_counter_0
        );

    \I__602\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3455\
        );

    \I__601\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3452\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3455\,
            I => \CounterZ0Z_4\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3452\,
            I => \CounterZ0Z_4\
        );

    \I__598\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3443\
        );

    \I__597\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3440\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3443\,
            I => \CounterZ0Z_0\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3440\,
            I => \CounterZ0Z_0\
        );

    \I__594\ : InMux
    port map (
            O => \N__3435\,
            I => \N__3431\
        );

    \I__593\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3428\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3431\,
            I => \CounterZ0Z_3\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3428\,
            I => \CounterZ0Z_3\
        );

    \I__590\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3419\
        );

    \I__589\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3416\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3419\,
            I => \CounterZ0Z_2\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3416\,
            I => \CounterZ0Z_2\
        );

    \I__586\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3407\
        );

    \I__585\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3404\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3407\,
            I => \CounterZ0Z_1\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3404\,
            I => \CounterZ0Z_1\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3399\,
            I => \N__3395\
        );

    \I__581\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3392\
        );

    \I__580\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3389\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3392\,
            I => \CounterZ0Z_5\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3389\,
            I => \CounterZ0Z_5\
        );

    \I__577\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3381\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3381\,
            I => un2_counterlto4_2
        );

    \I__575\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3375\,
            I => un2_counterlt7
        );

    \I__573\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3368\
        );

    \I__572\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3365\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3368\,
            I => \CounterZ0Z_11\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3365\,
            I => \CounterZ0Z_11\
        );

    \I__569\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3356\
        );

    \I__568\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3353\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3356\,
            I => \CounterZ0Z_9\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3353\,
            I => \CounterZ0Z_9\
        );

    \I__565\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3344\
        );

    \I__564\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3341\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3344\,
            I => \CounterZ0Z_10\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3341\,
            I => \CounterZ0Z_10\
        );

    \I__561\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3333\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3333\,
            I => un2_counterlto11_1
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3330\,
            I => \N_83_cascade_\
        );

    \I__558\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3324\,
            I => \N__3319\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__3323\,
            I => \N__3315\
        );

    \I__555\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3312\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__3319\,
            I => \N__3309\
        );

    \I__553\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3304\
        );

    \I__552\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3304\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3312\,
            I => \N_85\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__3309\,
            I => \N_85\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3304\,
            I => \N_85\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3297\,
            I => \un13lto4_i_1_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3291\,
            I => \un3_y_cry_1_THRU_CO\
        );

    \I__545\ : InMux
    port map (
            O => \N__3288\,
            I => un3_y_cry_1
        );

    \I__544\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3281\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3284\,
            I => \N__3277\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3281\,
            I => \N__3272\
        );

    \I__541\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3269\
        );

    \I__540\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3266\
        );

    \I__539\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3263\
        );

    \I__538\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3260\
        );

    \I__537\ : Span4Mux_s1_v
    port map (
            O => \N__3272\,
            I => \N__3257\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3254\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3266\,
            I => \yZ0Z_3\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3263\,
            I => \yZ0Z_3\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3260\,
            I => \yZ0Z_3\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__3257\,
            I => \yZ0Z_3\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__3254\,
            I => \yZ0Z_3\
        );

    \I__530\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3240\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3240\,
            I => \un3_y_cry_2_THRU_CO\
        );

    \I__528\ : InMux
    port map (
            O => \N__3237\,
            I => un3_y_cry_2
        );

    \I__527\ : InMux
    port map (
            O => \N__3234\,
            I => \N__3230\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3230\,
            I => \N__3222\
        );

    \I__524\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3219\
        );

    \I__523\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3216\
        );

    \I__522\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3213\
        );

    \I__521\ : Span4Mux_s1_h
    port map (
            O => \N__3222\,
            I => \N__3208\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3219\,
            I => \N__3208\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3216\,
            I => \yZ0Z_4\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3213\,
            I => \yZ0Z_4\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__3208\,
            I => \yZ0Z_4\
        );

    \I__516\ : InMux
    port map (
            O => \N__3201\,
            I => un3_y_cry_3
        );

    \I__515\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3195\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3195\,
            I => \N__3189\
        );

    \I__513\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3186\
        );

    \I__512\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3183\
        );

    \I__511\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3180\
        );

    \I__510\ : Span4Mux_s3_v
    port map (
            O => \N__3189\,
            I => \N__3177\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3186\,
            I => \N__3174\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3183\,
            I => \yZ0Z_5\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3180\,
            I => \yZ0Z_5\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3177\,
            I => \yZ0Z_5\
        );

    \I__505\ : Odrv4
    port map (
            O => \N__3174\,
            I => \yZ0Z_5\
        );

    \I__504\ : InMux
    port map (
            O => \N__3165\,
            I => un3_y_cry_4
        );

    \I__503\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3154\
        );

    \I__502\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3154\
        );

    \I__501\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3151\
        );

    \I__500\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3148\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3154\,
            I => \N__3145\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3151\,
            I => \yZ0Z_6\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3148\,
            I => \yZ0Z_6\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__3145\,
            I => \yZ0Z_6\
        );

    \I__495\ : InMux
    port map (
            O => \N__3138\,
            I => un3_y_cry_5
        );

    \I__494\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3126\
        );

    \I__492\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3123\
        );

    \I__491\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3120\
        );

    \I__490\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3117\
        );

    \I__489\ : Span4Mux_s1_h
    port map (
            O => \N__3126\,
            I => \N__3114\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3123\,
            I => \yZ0Z_7\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3120\,
            I => \yZ0Z_7\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3117\,
            I => \yZ0Z_7\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__3114\,
            I => \yZ0Z_7\
        );

    \I__484\ : InMux
    port map (
            O => \N__3105\,
            I => un3_y_cry_6
        );

    \I__483\ : InMux
    port map (
            O => \N__3102\,
            I => \N__3096\
        );

    \I__482\ : InMux
    port map (
            O => \N__3101\,
            I => \N__3093\
        );

    \I__481\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3088\
        );

    \I__480\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3088\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3096\,
            I => \yZ0Z_8\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3093\,
            I => \yZ0Z_8\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3088\,
            I => \yZ0Z_8\
        );

    \I__476\ : InMux
    port map (
            O => \N__3081\,
            I => un3_y_cry_7
        );

    \I__475\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3073\
        );

    \I__474\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3068\
        );

    \I__473\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3068\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3073\,
            I => \N_130\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3068\,
            I => \N_130\
        );

    \I__470\ : InMux
    port map (
            O => \N__3063\,
            I => \bfn_2_6_0_\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__468\ : InMux
    port map (
            O => \N__3057\,
            I => \N__3052\
        );

    \I__467\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3047\
        );

    \I__466\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3044\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3041\
        );

    \I__464\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3036\
        );

    \I__463\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3036\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3031\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3044\,
            I => \N__3031\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__3041\,
            I => \yZ0Z_9\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3036\,
            I => \yZ0Z_9\
        );

    \I__458\ : Odrv4
    port map (
            O => \N__3031\,
            I => \yZ0Z_9\
        );

    \I__457\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3020\
        );

    \I__456\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3017\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3020\,
            I => \CounterZ0Z_7\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3017\,
            I => \CounterZ0Z_7\
        );

    \I__453\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3008\
        );

    \I__452\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3005\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3008\,
            I => \CounterZ0Z_6\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3005\,
            I => \CounterZ0Z_6\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__3000\,
            I => \N__2996\
        );

    \I__448\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2993\
        );

    \I__447\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2990\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2993\,
            I => \CounterZ0Z_8\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2990\,
            I => \CounterZ0Z_8\
        );

    \I__444\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2982\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0\
        );

    \I__442\ : InMux
    port map (
            O => \N__2979\,
            I => un2_y_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__441\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2973\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2973\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0\
        );

    \I__439\ : InMux
    port map (
            O => \N__2970\,
            I => un2_y_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__438\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2960\
        );

    \I__437\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2960\
        );

    \I__436\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2957\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2960\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2957\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0\
        );

    \I__433\ : InMux
    port map (
            O => \N__2952\,
            I => un2_y_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__432\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2946\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\
        );

    \I__430\ : InMux
    port map (
            O => \N__2943\,
            I => un2_y_if_generate_plus_mult1_un26_sum_cry_5
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__2940\,
            I => \N__2936\
        );

    \I__428\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2927\
        );

    \I__427\ : InMux
    port map (
            O => \N__2936\,
            I => \N__2927\
        );

    \I__426\ : InMux
    port map (
            O => \N__2935\,
            I => \N__2927\
        );

    \I__425\ : InMux
    port map (
            O => \N__2934\,
            I => \N__2924\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2927\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2924\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__2919\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__2916\,
            I => \N__2913\
        );

    \I__420\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2910\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2910\,
            I => un2_y_if_generate_plus_mult1_un33_sum_i_7
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__2907\,
            I => \N__2903\
        );

    \I__417\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2900\
        );

    \I__416\ : InMux
    port map (
            O => \N__2903\,
            I => \N__2897\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2900\,
            I => \N_140\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2897\,
            I => \N_140\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__412\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2886\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2886\,
            I => un2_y_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__2883\,
            I => \N__2877\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__2882\,
            I => \N__2874\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__2881\,
            I => \N__2871\
        );

    \I__407\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2864\
        );

    \I__406\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2864\
        );

    \I__405\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2864\
        );

    \I__404\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2861\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2864\,
            I => \yZ0Z_0\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2861\,
            I => \yZ0Z_0\
        );

    \I__401\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2853\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2\
        );

    \I__399\ : InMux
    port map (
            O => \N__2850\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__398\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2844\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__2841\,
            I => \N__2838\
        );

    \I__395\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2835\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2835\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573\
        );

    \I__393\ : InMux
    port map (
            O => \N__2832\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__2829\,
            I => \N__2825\
        );

    \I__391\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2816\
        );

    \I__390\ : InMux
    port map (
            O => \N__2825\,
            I => \N__2816\
        );

    \I__389\ : InMux
    port map (
            O => \N__2824\,
            I => \N__2816\
        );

    \I__388\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2813\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2816\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2813\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__2808\,
            I => \N__2805\
        );

    \I__384\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2802\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31\
        );

    \I__382\ : InMux
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2796\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3\
        );

    \I__380\ : InMux
    port map (
            O => \N__2793\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__379\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2787\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__376\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2778\,
            I => un2_y_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__374\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2772\,
            I => un2_y_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__372\ : InMux
    port map (
            O => \N__2769\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__371\ : InMux
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2763\,
            I => un2_y_if_generate_plus_mult1_un47_sum_axb_7
        );

    \I__369\ : InMux
    port map (
            O => \N__2760\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__2757\,
            I => \N__2753\
        );

    \I__367\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2744\
        );

    \I__366\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2744\
        );

    \I__365\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2744\
        );

    \I__364\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2741\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2744\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2741\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__2736\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__359\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2727\,
            I => un2_y_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__356\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2718\,
            I => un2_y_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__354\ : InMux
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2712\,
            I => un2_y_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__352\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2706\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2706\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14\
        );

    \I__350\ : InMux
    port map (
            O => \N__2703\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__348\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2694\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2694\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6\
        );

    \I__346\ : InMux
    port map (
            O => \N__2691\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__345\ : InMux
    port map (
            O => \N__2688\,
            I => \N__2685\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2685\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6\
        );

    \I__343\ : InMux
    port map (
            O => \N__2682\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__342\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2676\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2676\,
            I => un2_y_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__340\ : InMux
    port map (
            O => \N__2673\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__339\ : InMux
    port map (
            O => \N__2670\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2667\,
            I => \N__2663\
        );

    \I__337\ : InMux
    port map (
            O => \N__2666\,
            I => \N__2654\
        );

    \I__336\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2654\
        );

    \I__335\ : InMux
    port map (
            O => \N__2662\,
            I => \N__2654\
        );

    \I__334\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2651\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2654\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2651\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__2646\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__2643\,
            I => \N__2640\
        );

    \I__329\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2637\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2637\,
            I => un2_y_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__327\ : InMux
    port map (
            O => \N__2634\,
            I => \Counter_cry_12\
        );

    \I__326\ : IoInMux
    port map (
            O => \N__2631\,
            I => \N__2628\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__324\ : IoSpan4Mux
    port map (
            O => \N__2625\,
            I => \N__2621\
        );

    \I__323\ : InMux
    port map (
            O => \N__2624\,
            I => \N__2618\
        );

    \I__322\ : Odrv4
    port map (
            O => \N__2621\,
            I => \ClockVGAZ0\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2618\,
            I => \ClockVGAZ0\
        );

    \I__320\ : ClkMux
    port map (
            O => \N__2613\,
            I => \N__2607\
        );

    \I__319\ : ClkMux
    port map (
            O => \N__2612\,
            I => \N__2607\
        );

    \I__318\ : GlobalMux
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__317\ : gio2CtrlBuf
    port map (
            O => \N__2604\,
            I => \Clock12MHz_c_g\
        );

    \I__316\ : SRMux
    port map (
            O => \N__2601\,
            I => \N__2597\
        );

    \I__315\ : SRMux
    port map (
            O => \N__2600\,
            I => \N__2594\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2597\,
            I => \N__2589\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2594\,
            I => \N__2586\
        );

    \I__312\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2581\
        );

    \I__311\ : InMux
    port map (
            O => \N__2592\,
            I => \N__2581\
        );

    \I__310\ : Odrv12
    port map (
            O => \N__2589\,
            I => \G_167\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__2586\,
            I => \G_167\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2581\,
            I => \G_167\
        );

    \I__307\ : InMux
    port map (
            O => \N__2574\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2571\,
            I => \N__2568\
        );

    \I__305\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2565\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2565\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0\
        );

    \I__303\ : InMux
    port map (
            O => \N__2562\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__302\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2556\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2556\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0\
        );

    \I__300\ : InMux
    port map (
            O => \N__2553\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__299\ : InMux
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2547\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2544\,
            I => \N__2539\
        );

    \I__296\ : CascadeMux
    port map (
            O => \N__2543\,
            I => \N__2535\
        );

    \I__295\ : InMux
    port map (
            O => \N__2542\,
            I => \N__2531\
        );

    \I__294\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2522\
        );

    \I__293\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2522\
        );

    \I__292\ : InMux
    port map (
            O => \N__2535\,
            I => \N__2522\
        );

    \I__291\ : InMux
    port map (
            O => \N__2534\,
            I => \N__2522\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2531\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2522\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2517\,
            I => \N__2514\
        );

    \I__287\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2511\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2511\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\
        );

    \I__285\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2505\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2505\,
            I => un2_y_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__283\ : InMux
    port map (
            O => \N__2502\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__282\ : InMux
    port map (
            O => \N__2499\,
            I => \Counter_cry_3\
        );

    \I__281\ : InMux
    port map (
            O => \N__2496\,
            I => \Counter_cry_4\
        );

    \I__280\ : InMux
    port map (
            O => \N__2493\,
            I => \Counter_cry_5\
        );

    \I__279\ : InMux
    port map (
            O => \N__2490\,
            I => \Counter_cry_6\
        );

    \I__278\ : InMux
    port map (
            O => \N__2487\,
            I => \bfn_1_7_0_\
        );

    \I__277\ : InMux
    port map (
            O => \N__2484\,
            I => \Counter_cry_8\
        );

    \I__276\ : InMux
    port map (
            O => \N__2481\,
            I => \Counter_cry_9\
        );

    \I__275\ : InMux
    port map (
            O => \N__2478\,
            I => \Counter_cry_10\
        );

    \I__274\ : InMux
    port map (
            O => \N__2475\,
            I => \Counter_cry_11\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2472\,
            I => \un13_x_i_i_a2_0_3_cascade_\
        );

    \I__272\ : InMux
    port map (
            O => \N__2469\,
            I => \bfn_1_6_0_\
        );

    \I__271\ : InMux
    port map (
            O => \N__2466\,
            I => \Counter_cry_0\
        );

    \I__270\ : InMux
    port map (
            O => \N__2463\,
            I => \Counter_cry_1\
        );

    \I__269\ : InMux
    port map (
            O => \N__2460\,
            I => \Counter_cry_2\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__267\ : InMux
    port map (
            O => \N__2454\,
            I => \N__2451\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2451\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\
        );

    \I__265\ : InMux
    port map (
            O => \N__2448\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__264\ : InMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2442\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0\
        );

    \I__262\ : InMux
    port map (
            O => \N__2439\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__261\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2433\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2433\,
            I => un2_y_if_generate_plus_mult1_un40_sum_axb_7
        );

    \I__259\ : InMux
    port map (
            O => \N__2430\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__258\ : InMux
    port map (
            O => \N__2427\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2424\,
            I => \N__2421\
        );

    \I__256\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2418\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2418\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0\
        );

    \I__254\ : CascadeMux
    port map (
            O => \N__2415\,
            I => \N__2412\
        );

    \I__253\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2409\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2409\,
            I => un2_y_if_generate_plus_mult1_un33_sum_i_0
        );

    \I__251\ : InMux
    port map (
            O => \N__2406\,
            I => \N__2403\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2403\,
            I => \N__2400\
        );

    \I__249\ : Odrv12
    port map (
            O => \N__2400\,
            I => un13_x_i_i_a2_1
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2397\,
            I => \N_130_cascade_\
        );

    \I__247\ : InMux
    port map (
            O => \N__2394\,
            I => \N__2391\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2391\,
            I => \y_RNIA5P7Z0Z_9\
        );

    \I__245\ : InMux
    port map (
            O => \N__2388\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__244\ : InMux
    port map (
            O => \N__2385\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__243\ : InMux
    port map (
            O => \N__2382\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__242\ : InMux
    port map (
            O => \N__2379\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__241\ : InMux
    port map (
            O => \N__2376\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__2373\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_\
        );

    \I__239\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2367\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2367\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\
        );

    \I__237\ : InMux
    port map (
            O => \N__2364\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__2361\,
            I => \N__2358\
        );

    \I__235\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2355\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2355\,
            I => un2_y_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__233\ : InMux
    port map (
            O => \N__2352\,
            I => \N__2349\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2349\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7\
        );

    \I__231\ : InMux
    port map (
            O => \N__2346\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__230\ : CascadeMux
    port map (
            O => \N__2343\,
            I => \N__2340\
        );

    \I__229\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2337\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2337\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0\
        );

    \I__227\ : InMux
    port map (
            O => \N__2334\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__226\ : InMux
    port map (
            O => \N__2331\,
            I => \N__2328\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2328\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0\
        );

    \I__224\ : InMux
    port map (
            O => \N__2325\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__223\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2319\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2319\,
            I => un2_y_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__221\ : InMux
    port map (
            O => \N__2316\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__220\ : InMux
    port map (
            O => \N__2313\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__2310\,
            I => \N__2305\
        );

    \I__218\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2301\
        );

    \I__217\ : InMux
    port map (
            O => \N__2308\,
            I => \N__2294\
        );

    \I__216\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2294\
        );

    \I__215\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2294\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2301\,
            I => \N__2291\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2294\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0\
        );

    \I__212\ : Odrv4
    port map (
            O => \N__2291\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0\
        );

    \I__211\ : CascadeMux
    port map (
            O => \N__2286\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_\
        );

    \I__210\ : CascadeMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__209\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__2277\,
            I => un2_y_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__206\ : InMux
    port map (
            O => \N__2271\,
            I => \N__2268\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2268\,
            I => un2_y_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__204\ : InMux
    port map (
            O => \N__2265\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__203\ : InMux
    port map (
            O => \N__2262\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__202\ : InMux
    port map (
            O => \N__2259\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__201\ : InMux
    port map (
            O => \N__2256\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__200\ : InMux
    port map (
            O => \N__2253\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_6
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un3_y_cry_8,
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_1_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_5_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_1_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_6_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_1_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un16_x_cry_8,
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_1_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_1_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Counter_cry_7\,
            carryinitout => \bfn_1_7_0_\
        );

    \ClockVGA_derived_clock_RNIND52\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2631\,
            GLOBALBUFFEROUTPUT => \ClockVGA_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \y_RNI7THF_3_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__3706\,
            in1 => \N__3280\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un13_x_i_i_a2_1,
            ltout => OPEN,
            carryin => \bfn_1_1_0_\,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NF_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2304\,
            in2 => \N__2361\,
            in3 => \N__2265\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3N_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2352\,
            in2 => \N__2310\,
            in3 => \N__2262\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1R_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2308\,
            in2 => \N__2343\,
            in3 => \N__2259\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8LRER1_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2542\,
            in1 => \N__2331\,
            in2 => \N__2283\,
            in3 => \N__2256\,
            lcout => un2_y_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUT_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2322\,
            in2 => \_gnd_net_\,
            in3 => \N__2253\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3234\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3233\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNP7_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2662\,
            in2 => \N__2274\,
            in3 => \N__2346\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONB_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2709\,
            in2 => \N__2667\,
            in3 => \N__2334\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66E_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2666\,
            in2 => \N__2700\,
            in3 => \N__2325\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHL7KT_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2309\,
            in1 => \N__2688\,
            in2 => \N__2643\,
            in3 => \N__2316\,
            lcout => un2_y_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2679\,
            in2 => \_gnd_net_\,
            in3 => \N__2313\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0\,
            ltout => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2286\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3198\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3135\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LP_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2935\,
            in2 => \N__2415\,
            in3 => \N__2388\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QD31_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2370\,
            in2 => \N__2940\,
            in3 => \N__2385\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HA81_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2939\,
            in2 => \N__2457\,
            in3 => \N__2382\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNI5DAA3_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2823\,
            in1 => \N__2445\,
            in2 => \N__2916\,
            in3 => \N__2379\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2436\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12\,
            ltout => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_0_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2373\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3099\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2394\,
            in2 => \N__4706\,
            in3 => \N__2364\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2985\,
            in2 => \N__4709\,
            in3 => \N__2448\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHF_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2976\,
            in2 => \N__4707\,
            in3 => \N__2439\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIM3MO1_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2934\,
            in1 => \N__2967\,
            in2 => \N__2424\,
            in3 => \N__2430\,
            lcout => un2_y_if_generate_plus_mult1_un40_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2427\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBP_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__2965\,
            in1 => \N__2966\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_sbtinv_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un33_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIN6QD2_0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2406\,
            in1 => \N__2906\,
            in2 => \N__2882\,
            in3 => \N__3051\,
            lcout => \N_130\,
            ltout => \N_130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2880\,
            in2 => \N__2397\,
            in3 => \N__4157\,
            lcout => \yZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIA5P7_9_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3050\,
            lcout => \y_RNIA5P7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_2_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011110000"
        )
    port map (
            in0 => \N__3294\,
            in1 => \N__3076\,
            in2 => \N__3704\,
            in3 => \N__4158\,
            lcout => \yZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_1_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__4156\,
            in1 => \_gnd_net_\,
            in2 => \N__2883\,
            in3 => \N__3318\,
            lcout => \N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIO44V_1_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3192\,
            in1 => \N__3159\,
            in2 => \N__3323\,
            in3 => \N__3101\,
            lcout => OPEN,
            ltout => \un13_x_i_i_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNI58ME1_4_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3225\,
            in2 => \N__2472\,
            in3 => \N__3130\,
            lcout => \N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_3_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011110000"
        )
    port map (
            in0 => \N__3243\,
            in1 => \N__3077\,
            in2 => \N__3284\,
            in3 => \N__4159\,
            lcout => \yZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3510\,
            in1 => \N__3447\,
            in2 => \_gnd_net_\,
            in3 => \N__2469\,
            lcout => \CounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \Counter_cry_0\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3502\,
            in1 => \N__3411\,
            in2 => \_gnd_net_\,
            in3 => \N__2466\,
            lcout => \CounterZ0Z_1\,
            ltout => OPEN,
            carryin => \Counter_cry_0\,
            carryout => \Counter_cry_1\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_2_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3511\,
            in1 => \N__3423\,
            in2 => \_gnd_net_\,
            in3 => \N__2463\,
            lcout => \CounterZ0Z_2\,
            ltout => OPEN,
            carryin => \Counter_cry_1\,
            carryout => \Counter_cry_2\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_3_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3503\,
            in1 => \N__3435\,
            in2 => \_gnd_net_\,
            in3 => \N__2460\,
            lcout => \CounterZ0Z_3\,
            ltout => OPEN,
            carryin => \Counter_cry_2\,
            carryout => \Counter_cry_3\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_4_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3512\,
            in1 => \N__3459\,
            in2 => \_gnd_net_\,
            in3 => \N__2499\,
            lcout => \CounterZ0Z_4\,
            ltout => OPEN,
            carryin => \Counter_cry_3\,
            carryout => \Counter_cry_4\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3504\,
            in1 => \N__3398\,
            in2 => \_gnd_net_\,
            in3 => \N__2496\,
            lcout => \CounterZ0Z_5\,
            ltout => OPEN,
            carryin => \Counter_cry_4\,
            carryout => \Counter_cry_5\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3513\,
            in1 => \N__3012\,
            in2 => \_gnd_net_\,
            in3 => \N__2493\,
            lcout => \CounterZ0Z_6\,
            ltout => OPEN,
            carryin => \Counter_cry_5\,
            carryout => \Counter_cry_6\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3505\,
            in1 => \N__3024\,
            in2 => \_gnd_net_\,
            in3 => \N__2490\,
            lcout => \CounterZ0Z_7\,
            ltout => OPEN,
            carryin => \Counter_cry_6\,
            carryout => \Counter_cry_7\,
            clk => \N__2613\,
            ce => 'H',
            sr => \N__2601\
        );

    \Counter_8_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3516\,
            in1 => \N__2999\,
            in2 => \_gnd_net_\,
            in3 => \N__2487\,
            lcout => \CounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \Counter_cry_8\,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Counter_9_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3507\,
            in1 => \N__3360\,
            in2 => \_gnd_net_\,
            in3 => \N__2484\,
            lcout => \CounterZ0Z_9\,
            ltout => OPEN,
            carryin => \Counter_cry_8\,
            carryout => \Counter_cry_9\,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Counter_10_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3514\,
            in1 => \N__3348\,
            in2 => \_gnd_net_\,
            in3 => \N__2481\,
            lcout => \CounterZ0Z_10\,
            ltout => OPEN,
            carryin => \Counter_cry_9\,
            carryout => \Counter_cry_10\,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Counter_11_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3506\,
            in1 => \N__3372\,
            in2 => \_gnd_net_\,
            in3 => \N__2478\,
            lcout => \CounterZ0Z_11\,
            ltout => OPEN,
            carryin => \Counter_cry_10\,
            carryout => \Counter_cry_11\,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Counter_12_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3515\,
            in1 => \N__3531\,
            in2 => \_gnd_net_\,
            in3 => \N__2475\,
            lcout => \CounterZ0Z_12\,
            ltout => OPEN,
            carryin => \Counter_cry_11\,
            carryout => \Counter_cry_12\,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Counter_13_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3508\,
            in1 => \N__3543\,
            in2 => \_gnd_net_\,
            in3 => \N__2634\,
            lcout => \CounterZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \ClockVGA_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2624\,
            in2 => \_gnd_net_\,
            in3 => \N__3509\,
            lcout => \ClockVGAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2612\,
            ce => 'H',
            sr => \N__2600\
        );

    \Reset_latch_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2592\,
            in2 => \_gnd_net_\,
            in3 => \N__2593\,
            lcout => \G_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3705\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_1_0_\,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCU_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2715\,
            in2 => \N__2543\,
            in3 => \N__2574\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1ND1_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2538\,
            in2 => \N__2571\,
            in3 => \N__2562\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_4_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2559\,
            in2 => \N__2544\,
            in3 => \N__2553\,
            lcout => \Pixel_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2550\,
            in2 => \N__2517\,
            in3 => \N__2534\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFR1_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2508\,
            in2 => \_gnd_net_\,
            in3 => \N__2502\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3285\,
            lcout => un2_y_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3194\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2O14_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2752\,
            in2 => \N__2724\,
            in3 => \N__2703\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5G6_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2856\,
            in2 => \N__2757\,
            in3 => \N__2691\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3V6_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2756\,
            in2 => \N__2841\,
            in3 => \N__2682\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNIR1SME_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2661\,
            in1 => \N__2799\,
            in2 => \N__2733\,
            in3 => \N__2673\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2775\,
            in2 => \_gnd_net_\,
            in3 => \N__2670\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7\,
            ltout => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2646\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3161\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8O2_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2824\,
            in2 => \N__2892\,
            in3 => \N__2850\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNION573_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2847\,
            in2 => \N__2829\,
            in3 => \N__2832\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVG3_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2828\,
            in2 => \N__2808\,
            in3 => \N__2793\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI2VUB7_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2751\,
            in1 => \N__2790\,
            in2 => \N__2784\,
            in3 => \N__2769\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2766\,
            in2 => \_gnd_net_\,
            in3 => \N__2760\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3\,
            ltout => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_0_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2736\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3055\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => un2_y_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJC_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4688\,
            in2 => \N__4708\,
            in3 => \N__2979\,
            lcout => \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKC_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4699\,
            in2 => \_gnd_net_\,
            in3 => \N__2970\,
            lcout => \un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLC_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__2952\,
            lcout => \un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un26_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un26_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2949\,
            in2 => \_gnd_net_\,
            in3 => \N__2943\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0\,
            ltout => \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_0_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2919\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un33_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIMA162_9_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3056\,
            in1 => \N__3688\,
            in2 => \N__2907\,
            in3 => \N__3275\,
            lcout => \y_RNIMA162Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => un2_y_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un3_y_cry_1_c_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3322\,
            in2 => \N__2881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => un3_y_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un3_y_cry_1_THRU_LUT4_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3703\,
            in2 => \_gnd_net_\,
            in3 => \N__3288\,
            lcout => \un3_y_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => un3_y_cry_1,
            carryout => un3_y_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un3_y_cry_2_THRU_LUT4_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3276\,
            in2 => \_gnd_net_\,
            in3 => \N__3237\,
            lcout => \un3_y_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => un3_y_cry_2,
            carryout => un3_y_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4160\,
            in1 => \N__3226\,
            in2 => \_gnd_net_\,
            in3 => \N__3201\,
            lcout => \yZ0Z_4\,
            ltout => OPEN,
            carryin => un3_y_cry_3,
            carryout => un3_y_cry_4,
            clk => \N__4473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_5_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4163\,
            in1 => \N__3193\,
            in2 => \_gnd_net_\,
            in3 => \N__3165\,
            lcout => \yZ0Z_5\,
            ltout => OPEN,
            carryin => un3_y_cry_4,
            carryout => un3_y_cry_5,
            clk => \N__4473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_6_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__3160\,
            in2 => \_gnd_net_\,
            in3 => \N__3138\,
            lcout => \yZ0Z_6\,
            ltout => OPEN,
            carryin => un3_y_cry_5,
            carryout => un3_y_cry_6,
            clk => \N__4473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_7_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4164\,
            in1 => \N__3131\,
            in2 => \_gnd_net_\,
            in3 => \N__3105\,
            lcout => \yZ0Z_7\,
            ltout => OPEN,
            carryin => un3_y_cry_6,
            carryout => un3_y_cry_7,
            clk => \N__4473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_8_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4162\,
            in1 => \N__3102\,
            in2 => \_gnd_net_\,
            in3 => \N__3081\,
            lcout => \yZ0Z_8\,
            ltout => OPEN,
            carryin => un3_y_cry_7,
            carryout => un3_y_cry_8,
            clk => \N__4473\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_9_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__3078\,
            in1 => \N__4134\,
            in2 => \N__3060\,
            in3 => \N__3063\,
            lcout => \yZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_RNICJ474_6_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__3023\,
            in1 => \N__3011\,
            in2 => \N__3000\,
            in3 => \N__3378\,
            lcout => OPEN,
            ltout => \un2_counterlt11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_RNI7QMJ6_13_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__3542\,
            in1 => \N__3530\,
            in2 => \N__3519\,
            in3 => \N__3336\,
            lcout => un2_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_RNIVB1D1_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3458\,
            in1 => \N__3446\,
            in2 => \_gnd_net_\,
            in3 => \N__3434\,
            lcout => un2_counterlto4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_RNIVO2Q2_1_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3422\,
            in1 => \N__3410\,
            in2 => \N__3399\,
            in3 => \N__3384\,
            lcout => un2_counterlt7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Counter_RNI4CPD1_9_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3371\,
            in1 => \N__3359\,
            in2 => \_gnd_net_\,
            in3 => \N__3347\,
            lcout => un2_counterlto11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_11_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__3627\,
            in1 => \N__3644\,
            in2 => \_gnd_net_\,
            in3 => \N__3579\,
            lcout => OPEN,
            ltout => \N_83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_9_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110011111"
        )
    port map (
            in0 => \N__3580\,
            in1 => \N__3614\,
            in2 => \N__3330\,
            in3 => \N__3600\,
            lcout => OPEN,
            ltout => \un13lto4_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_5_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111101"
        )
    port map (
            in0 => \N__3327\,
            in1 => \N__3708\,
            in2 => \N__3297\,
            in3 => \N__3581\,
            lcout => \N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => \CONSTANT_ONE_NET_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_inv_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3657\,
            in2 => \N__3711\,
            in3 => \N__3707\,
            lcout => un2_y_if_generate_plus_mult1_un75_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3656\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_1_0_\,
            carryout => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_LUT4_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4642\,
            in2 => \N__3645\,
            in3 => \N__3621\,
            lcout => \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_LUT4_0_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3618\,
            in2 => \N__4662\,
            in3 => \N__3594\,
            lcout => \un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_0_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111101101111"
        )
    port map (
            in0 => \N__3591\,
            in1 => \N__3582\,
            in2 => \N__3561\,
            in3 => \N__3552\,
            lcout => \N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4215\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3788\,
            in2 => \N__3774\,
            in3 => \N__3549\,
            lcout => \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_6_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3897\,
            in2 => \N__3864\,
            in3 => \N__3546\,
            lcout => \Pixel_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3789\,
            in2 => \N__3888\,
            in3 => \N__3859\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__3780\,
            lcout => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\,
            ltout => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_10_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__4216\,
            in1 => \_gnd_net_\,
            in2 => \N__3777\,
            in3 => \N__3834\,
            lcout => \N_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI5UL6_5_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4278\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI6ANQ_1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3742\,
            in1 => \N__3762\,
            in2 => \N__3729\,
            in3 => \N__3832\,
            lcout => un11_x_0_a2_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_0_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3763\,
            lcout => \xZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_1_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3743\,
            lcout => \xZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4476\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un16_x_cry_1_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3765\,
            in2 => \N__3747\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => un16_x_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_2_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3728\,
            in2 => \_gnd_net_\,
            in3 => \N__3714\,
            lcout => \xZ0Z_2\,
            ltout => OPEN,
            carryin => un16_x_cry_1,
            carryout => un16_x_cry_2,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_3_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3833\,
            in2 => \_gnd_net_\,
            in3 => \N__3813\,
            lcout => \N_89\,
            ltout => OPEN,
            carryin => un16_x_cry_2,
            carryout => un16_x_cry_3,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_4_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4214\,
            in2 => \_gnd_net_\,
            in3 => \N__3810\,
            lcout => \xZ0Z_4\,
            ltout => OPEN,
            carryin => un16_x_cry_3,
            carryout => un16_x_cry_4,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_5_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4133\,
            in1 => \N__4276\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \xZ0Z_5\,
            ltout => OPEN,
            carryin => un16_x_cry_4,
            carryout => un16_x_cry_5,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_6_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4245\,
            in2 => \_gnd_net_\,
            in3 => \N__3804\,
            lcout => \xZ0Z_6\,
            ltout => OPEN,
            carryin => un16_x_cry_5,
            carryout => un16_x_cry_6,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_7_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4435\,
            in2 => \_gnd_net_\,
            in3 => \N__3801\,
            lcout => \xZ0Z_7\,
            ltout => OPEN,
            carryin => un16_x_cry_6,
            carryout => un16_x_cry_7,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_8_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__4546\,
            in2 => \_gnd_net_\,
            in3 => \N__3798\,
            lcout => \xZ0Z_8\,
            ltout => OPEN,
            carryin => un16_x_cry_7,
            carryout => un16_x_cry_8,
            clk => \N__4475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_9_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4089\,
            in1 => \N__4118\,
            in2 => \_gnd_net_\,
            in3 => \N__3795\,
            lcout => \xZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3845\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_1_0_\,
            carryout => un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_LUT4_0_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3966\,
            in3 => \N__3792\,
            lcout => \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_1_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101101111"
        )
    port map (
            in0 => \N__3954\,
            in1 => \N__3975\,
            in2 => \N__3930\,
            in3 => \N__3969\,
            lcout => \N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_7_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111111111"
        )
    port map (
            in0 => \N__3962\,
            in1 => \N__3953\,
            in2 => \N__3945\,
            in3 => \N__3936\,
            lcout => \N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__4311\,
            in1 => \N__3921\,
            in2 => \N__4323\,
            in3 => \N__3915\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4277\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4001\,
            in2 => \N__3993\,
            in3 => \N__3891\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4017\,
            in2 => \N__4053\,
            in3 => \N__3879\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3863\,
            in1 => \N__4002\,
            in2 => \N__4041\,
            in3 => \N__3870\,
            lcout => un2_x_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4029\,
            in2 => \_gnd_net_\,
            in3 => \N__3867\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_inv_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__3846\,
            in1 => \N__4687\,
            in2 => \_gnd_net_\,
            in3 => \N__4217\,
            lcout => un2_x_if_generate_plus_mult1_un75_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4240\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4349\,
            in2 => \N__3984\,
            in3 => \N__4044\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4365\,
            in2 => \N__4401\,
            in3 => \N__4032\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4016\,
            in1 => \N__4350\,
            in2 => \N__4389\,
            in3 => \N__4023\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4377\,
            in2 => \_gnd_net_\,
            in3 => \N__4020\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\,
            ltout => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4005\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI6VL6_6_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI70M6_7_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4432\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000010101"
        )
    port map (
            in0 => \N__4087\,
            in1 => \N__4434\,
            in2 => \N__4287\,
            in3 => \N__4547\,
            lcout => \Pixel_0_sqmuxa_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI92M6_9_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4085\,
            lcout => un2_x_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_2_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4502\,
            in1 => \N__4551\,
            in2 => \N__4179\,
            in3 => \N__4088\,
            lcout => \Pixel_0_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSyncZ0_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4275\,
            in1 => \N__4244\,
            in2 => \N__4442\,
            in3 => \N__4062\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_8_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4243\,
            in1 => \N__4213\,
            in2 => \_gnd_net_\,
            in3 => \N__4274\,
            lcout => \N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNIMQNQ_4_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__4242\,
            in2 => \N__4218\,
            in3 => \N__4433\,
            lcout => OPEN,
            ltout => \un11_x_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNID8R22_9_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4175\,
            in1 => \N__4550\,
            in2 => \N__4167\,
            in3 => \N__4086\,
            lcout => \x_RNID8R22Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_RNO_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4084\,
            in2 => \_gnd_net_\,
            in3 => \N__4545\,
            lcout => un1_xlto9_i_0,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => un2_x_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4056\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4446\,
            in3 => \_gnd_net_\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4443\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4580\,
            in2 => \N__4512\,
            in3 => \N__4392\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4596\,
            in2 => \N__4335\,
            in3 => \N__4380\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4364\,
            in1 => \N__4581\,
            in2 => \N__4620\,
            in3 => \N__4371\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4608\,
            in2 => \_gnd_net_\,
            in3 => \N__4368\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\,
            ltout => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4353\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4341\,
            in2 => \_gnd_net_\,
            in3 => \N__4326\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4716\,
            in2 => \N__4710\,
            in3 => \N__4611\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__4557\,
            in2 => \N__4572\,
            in3 => \N__4602\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4599\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\,
            ltout => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4584\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4567\,
            in2 => \_gnd_net_\,
            in3 => \N__4568\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI81M6_8_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSyncZ0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4503\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4478\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
