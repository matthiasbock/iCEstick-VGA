// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 24 2015 16:35:04

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSync,
    SCLK1,
    Pixel,
    HSync,
    nCS2,
    SDATA2,
    SCLK2,
    Clock12MHz,
    nCS1,
    SDATA1);

    output VSync;
    output SCLK1;
    output Pixel;
    output HSync;
    output nCS2;
    output SDATA2;
    output SCLK2;
    input Clock12MHz;
    output nCS1;
    input SDATA1;

    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15791;
    wire N__15790;
    wire N__15789;
    wire N__15782;
    wire N__15781;
    wire N__15780;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15764;
    wire N__15763;
    wire N__15762;
    wire N__15755;
    wire N__15754;
    wire N__15753;
    wire N__15746;
    wire N__15745;
    wire N__15744;
    wire N__15737;
    wire N__15736;
    wire N__15735;
    wire N__15718;
    wire N__15717;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15709;
    wire N__15708;
    wire N__15707;
    wire N__15706;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15672;
    wire N__15667;
    wire N__15662;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15606;
    wire N__15603;
    wire N__15602;
    wire N__15601;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15596;
    wire N__15593;
    wire N__15588;
    wire N__15587;
    wire N__15586;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15551;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15465;
    wire N__15462;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15417;
    wire N__15416;
    wire N__15413;
    wire N__15412;
    wire N__15409;
    wire N__15408;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15378;
    wire N__15377;
    wire N__15374;
    wire N__15369;
    wire N__15364;
    wire N__15363;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15351;
    wire N__15346;
    wire N__15343;
    wire N__15342;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15332;
    wire N__15327;
    wire N__15322;
    wire N__15321;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15294;
    wire N__15293;
    wire N__15292;
    wire N__15291;
    wire N__15290;
    wire N__15289;
    wire N__15286;
    wire N__15281;
    wire N__15280;
    wire N__15275;
    wire N__15274;
    wire N__15273;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15232;
    wire N__15223;
    wire N__15222;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15181;
    wire N__15180;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15155;
    wire N__15148;
    wire N__15145;
    wire N__15140;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15123;
    wire N__15122;
    wire N__15121;
    wire N__15116;
    wire N__15115;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15096;
    wire N__15093;
    wire N__15088;
    wire N__15083;
    wire N__15080;
    wire N__15075;
    wire N__15072;
    wire N__15067;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15059;
    wire N__15058;
    wire N__15057;
    wire N__15056;
    wire N__15053;
    wire N__15052;
    wire N__15049;
    wire N__15044;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15025;
    wire N__15020;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14983;
    wire N__14982;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14967;
    wire N__14966;
    wire N__14959;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14932;
    wire N__14923;
    wire N__14918;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14893;
    wire N__14890;
    wire N__14881;
    wire N__14880;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14873;
    wire N__14868;
    wire N__14861;
    wire N__14858;
    wire N__14851;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14847;
    wire N__14846;
    wire N__14843;
    wire N__14836;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14828;
    wire N__14827;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14800;
    wire N__14791;
    wire N__14790;
    wire N__14789;
    wire N__14788;
    wire N__14787;
    wire N__14786;
    wire N__14785;
    wire N__14784;
    wire N__14783;
    wire N__14782;
    wire N__14777;
    wire N__14770;
    wire N__14769;
    wire N__14766;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14747;
    wire N__14742;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14724;
    wire N__14719;
    wire N__14718;
    wire N__14717;
    wire N__14716;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14705;
    wire N__14704;
    wire N__14703;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14682;
    wire N__14677;
    wire N__14672;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14652;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14646;
    wire N__14643;
    wire N__14642;
    wire N__14633;
    wire N__14628;
    wire N__14625;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14610;
    wire N__14609;
    wire N__14608;
    wire N__14607;
    wire N__14606;
    wire N__14601;
    wire N__14596;
    wire N__14591;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14577;
    wire N__14574;
    wire N__14573;
    wire N__14572;
    wire N__14571;
    wire N__14570;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14556;
    wire N__14551;
    wire N__14542;
    wire N__14541;
    wire N__14540;
    wire N__14539;
    wire N__14538;
    wire N__14537;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14527;
    wire N__14522;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14508;
    wire N__14505;
    wire N__14500;
    wire N__14495;
    wire N__14490;
    wire N__14487;
    wire N__14482;
    wire N__14479;
    wire N__14474;
    wire N__14471;
    wire N__14466;
    wire N__14463;
    wire N__14460;
    wire N__14455;
    wire N__14452;
    wire N__14443;
    wire N__14442;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14434;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14411;
    wire N__14408;
    wire N__14395;
    wire N__14394;
    wire N__14391;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14374;
    wire N__14371;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14359;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14351;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14345;
    wire N__14344;
    wire N__14343;
    wire N__14342;
    wire N__14341;
    wire N__14340;
    wire N__14339;
    wire N__14336;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14280;
    wire N__14279;
    wire N__14278;
    wire N__14277;
    wire N__14276;
    wire N__14275;
    wire N__14274;
    wire N__14269;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14260;
    wire N__14257;
    wire N__14252;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14230;
    wire N__14225;
    wire N__14220;
    wire N__14213;
    wire N__14210;
    wire N__14203;
    wire N__14202;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14142;
    wire N__14137;
    wire N__14134;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14110;
    wire N__14109;
    wire N__14108;
    wire N__14107;
    wire N__14106;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14094;
    wire N__14089;
    wire N__14084;
    wire N__14081;
    wire N__14074;
    wire N__14059;
    wire N__14058;
    wire N__14057;
    wire N__14056;
    wire N__14055;
    wire N__14054;
    wire N__14053;
    wire N__14050;
    wire N__14049;
    wire N__14048;
    wire N__14047;
    wire N__14046;
    wire N__14045;
    wire N__14044;
    wire N__14043;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14035;
    wire N__14032;
    wire N__14025;
    wire N__14022;
    wire N__14017;
    wire N__14010;
    wire N__14003;
    wire N__14000;
    wire N__13995;
    wire N__13978;
    wire N__13975;
    wire N__13974;
    wire N__13973;
    wire N__13970;
    wire N__13965;
    wire N__13960;
    wire N__13957;
    wire N__13956;
    wire N__13955;
    wire N__13954;
    wire N__13951;
    wire N__13950;
    wire N__13949;
    wire N__13948;
    wire N__13945;
    wire N__13940;
    wire N__13937;
    wire N__13930;
    wire N__13921;
    wire N__13918;
    wire N__13917;
    wire N__13916;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13908;
    wire N__13905;
    wire N__13904;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13889;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13855;
    wire N__13852;
    wire N__13851;
    wire N__13850;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13838;
    wire N__13831;
    wire N__13828;
    wire N__13827;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13797;
    wire N__13796;
    wire N__13793;
    wire N__13788;
    wire N__13783;
    wire N__13782;
    wire N__13781;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13762;
    wire N__13759;
    wire N__13758;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13736;
    wire N__13729;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13702;
    wire N__13699;
    wire N__13698;
    wire N__13697;
    wire N__13696;
    wire N__13695;
    wire N__13692;
    wire N__13687;
    wire N__13682;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13635;
    wire N__13632;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13594;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13577;
    wire N__13570;
    wire N__13569;
    wire N__13568;
    wire N__13565;
    wire N__13564;
    wire N__13561;
    wire N__13560;
    wire N__13557;
    wire N__13548;
    wire N__13543;
    wire N__13540;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13530;
    wire N__13529;
    wire N__13526;
    wire N__13521;
    wire N__13520;
    wire N__13519;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13481;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13466;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13452;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13440;
    wire N__13435;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13422;
    wire N__13421;
    wire N__13420;
    wire N__13419;
    wire N__13418;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13392;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13360;
    wire N__13355;
    wire N__13352;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13296;
    wire N__13295;
    wire N__13294;
    wire N__13291;
    wire N__13290;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13284;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13276;
    wire N__13273;
    wire N__13268;
    wire N__13267;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13262;
    wire N__13259;
    wire N__13258;
    wire N__13257;
    wire N__13256;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13248;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13232;
    wire N__13227;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13213;
    wire N__13210;
    wire N__13205;
    wire N__13202;
    wire N__13201;
    wire N__13198;
    wire N__13197;
    wire N__13194;
    wire N__13187;
    wire N__13180;
    wire N__13175;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13152;
    wire N__13147;
    wire N__13140;
    wire N__13135;
    wire N__13132;
    wire N__13127;
    wire N__13114;
    wire N__13113;
    wire N__13110;
    wire N__13109;
    wire N__13108;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13076;
    wire N__13075;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13056;
    wire N__13055;
    wire N__13052;
    wire N__13045;
    wire N__13038;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13006;
    wire N__13003;
    wire N__12998;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12982;
    wire N__12975;
    wire N__12968;
    wire N__12965;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12933;
    wire N__12932;
    wire N__12931;
    wire N__12930;
    wire N__12927;
    wire N__12926;
    wire N__12923;
    wire N__12922;
    wire N__12921;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12917;
    wire N__12914;
    wire N__12913;
    wire N__12912;
    wire N__12911;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12892;
    wire N__12889;
    wire N__12888;
    wire N__12887;
    wire N__12886;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12877;
    wire N__12876;
    wire N__12875;
    wire N__12872;
    wire N__12867;
    wire N__12862;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12858;
    wire N__12857;
    wire N__12856;
    wire N__12853;
    wire N__12848;
    wire N__12839;
    wire N__12838;
    wire N__12835;
    wire N__12830;
    wire N__12825;
    wire N__12822;
    wire N__12815;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12799;
    wire N__12796;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12756;
    wire N__12751;
    wire N__12750;
    wire N__12747;
    wire N__12746;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12725;
    wire N__12718;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12700;
    wire N__12695;
    wire N__12676;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12670;
    wire N__12669;
    wire N__12666;
    wire N__12665;
    wire N__12664;
    wire N__12661;
    wire N__12660;
    wire N__12657;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12642;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12636;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12617;
    wire N__12608;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12589;
    wire N__12588;
    wire N__12587;
    wire N__12586;
    wire N__12585;
    wire N__12582;
    wire N__12575;
    wire N__12572;
    wire N__12563;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12538;
    wire N__12535;
    wire N__12534;
    wire N__12533;
    wire N__12532;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12516;
    wire N__12513;
    wire N__12508;
    wire N__12501;
    wire N__12496;
    wire N__12489;
    wire N__12482;
    wire N__12463;
    wire N__12460;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12452;
    wire N__12447;
    wire N__12442;
    wire N__12441;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12435;
    wire N__12434;
    wire N__12433;
    wire N__12432;
    wire N__12429;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12406;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12398;
    wire N__12395;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12377;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12357;
    wire N__12352;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12310;
    wire N__12309;
    wire N__12308;
    wire N__12307;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12303;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12285;
    wire N__12280;
    wire N__12271;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12192;
    wire N__12175;
    wire N__12172;
    wire N__12171;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12153;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12137;
    wire N__12132;
    wire N__12127;
    wire N__12122;
    wire N__12109;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12099;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12051;
    wire N__12046;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12018;
    wire N__12015;
    wire N__12014;
    wire N__12011;
    wire N__12006;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11985;
    wire N__11984;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11884;
    wire N__11881;
    wire N__11880;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11857;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11684;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11654;
    wire N__11653;
    wire N__11652;
    wire N__11647;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11642;
    wire N__11641;
    wire N__11638;
    wire N__11633;
    wire N__11630;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11590;
    wire N__11589;
    wire N__11586;
    wire N__11581;
    wire N__11576;
    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11526;
    wire N__11525;
    wire N__11522;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11415;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11328;
    wire N__11327;
    wire N__11324;
    wire N__11323;
    wire N__11320;
    wire N__11319;
    wire N__11316;
    wire N__11307;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11238;
    wire N__11235;
    wire N__11230;
    wire N__11229;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11176;
    wire N__11171;
    wire N__11168;
    wire N__11167;
    wire N__11164;
    wire N__11159;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11147;
    wire N__11144;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11119;
    wire N__11116;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11092;
    wire N__11085;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11043;
    wire N__11038;
    wire N__11035;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11023;
    wire N__11020;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11008;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10993;
    wire N__10992;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10974;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10874;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10819;
    wire N__10816;
    wire N__10815;
    wire N__10814;
    wire N__10811;
    wire N__10810;
    wire N__10807;
    wire N__10802;
    wire N__10799;
    wire N__10792;
    wire N__10791;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10701;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10603;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10593;
    wire N__10592;
    wire N__10591;
    wire N__10586;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10556;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10461;
    wire N__10460;
    wire N__10459;
    wire N__10454;
    wire N__10449;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10440;
    wire N__10437;
    wire N__10432;
    wire N__10429;
    wire N__10420;
    wire N__10419;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10371;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10344;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10338;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10330;
    wire N__10327;
    wire N__10326;
    wire N__10323;
    wire N__10318;
    wire N__10315;
    wire N__10308;
    wire N__10305;
    wire N__10300;
    wire N__10297;
    wire N__10292;
    wire N__10289;
    wire N__10284;
    wire N__10279;
    wire N__10278;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10266;
    wire N__10265;
    wire N__10264;
    wire N__10257;
    wire N__10254;
    wire N__10253;
    wire N__10250;
    wire N__10245;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10223;
    wire N__10218;
    wire N__10215;
    wire N__10214;
    wire N__10209;
    wire N__10206;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10185;
    wire N__10182;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10121;
    wire N__10120;
    wire N__10119;
    wire N__10118;
    wire N__10117;
    wire N__10112;
    wire N__10107;
    wire N__10100;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10080;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10005;
    wire N__10004;
    wire N__10003;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9978;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9870;
    wire N__9867;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9846;
    wire N__9843;
    wire N__9842;
    wire N__9841;
    wire N__9840;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9813;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9747;
    wire N__9744;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9732;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9696;
    wire N__9693;
    wire N__9692;
    wire N__9689;
    wire N__9684;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9511;
    wire N__9510;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9488;
    wire N__9483;
    wire N__9480;
    wire N__9473;
    wire N__9468;
    wire N__9467;
    wire N__9464;
    wire N__9459;
    wire N__9458;
    wire N__9455;
    wire N__9446;
    wire N__9443;
    wire N__9438;
    wire N__9435;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9318;
    wire N__9317;
    wire N__9316;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9305;
    wire N__9300;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9278;
    wire N__9275;
    wire N__9270;
    wire N__9265;
    wire N__9262;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9198;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9172;
    wire N__9169;
    wire N__9168;
    wire N__9165;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9145;
    wire N__9144;
    wire N__9139;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9133;
    wire N__9132;
    wire N__9127;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9105;
    wire N__9104;
    wire N__9101;
    wire N__9100;
    wire N__9099;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9074;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9033;
    wire N__9030;
    wire N__9025;
    wire N__9024;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8974;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8961;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8907;
    wire N__8906;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8902;
    wire N__8895;
    wire N__8888;
    wire N__8885;
    wire N__8880;
    wire N__8879;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8723;
    wire N__8718;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8697;
    wire N__8692;
    wire N__8691;
    wire N__8686;
    wire N__8685;
    wire N__8684;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8664;
    wire N__8661;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8541;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8520;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8499;
    wire N__8496;
    wire N__8491;
    wire N__8488;
    wire N__8487;
    wire N__8486;
    wire N__8483;
    wire N__8478;
    wire N__8475;
    wire N__8470;
    wire N__8469;
    wire N__8466;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8440;
    wire N__8439;
    wire N__8436;
    wire N__8435;
    wire N__8434;
    wire N__8431;
    wire N__8430;
    wire N__8429;
    wire N__8424;
    wire N__8421;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8406;
    wire N__8405;
    wire N__8402;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8376;
    wire N__8373;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8327;
    wire N__8326;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8303;
    wire N__8300;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8184;
    wire N__8183;
    wire N__8180;
    wire N__8175;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8142;
    wire N__8141;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8122;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8089;
    wire N__8088;
    wire N__8087;
    wire N__8084;
    wire N__8079;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7961;
    wire N__7960;
    wire N__7957;
    wire N__7952;
    wire N__7949;
    wire N__7948;
    wire N__7945;
    wire N__7940;
    wire N__7939;
    wire N__7934;
    wire N__7931;
    wire N__7930;
    wire N__7927;
    wire N__7922;
    wire N__7919;
    wire N__7914;
    wire N__7913;
    wire N__7910;
    wire N__7903;
    wire N__7900;
    wire N__7899;
    wire N__7896;
    wire N__7895;
    wire N__7894;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7875;
    wire N__7872;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7839;
    wire N__7838;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7826;
    wire N__7825;
    wire N__7824;
    wire N__7823;
    wire N__7822;
    wire N__7821;
    wire N__7816;
    wire N__7815;
    wire N__7814;
    wire N__7813;
    wire N__7812;
    wire N__7809;
    wire N__7808;
    wire N__7805;
    wire N__7800;
    wire N__7795;
    wire N__7792;
    wire N__7783;
    wire N__7780;
    wire N__7775;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7757;
    wire N__7756;
    wire N__7753;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7745;
    wire N__7742;
    wire N__7741;
    wire N__7740;
    wire N__7739;
    wire N__7738;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7724;
    wire N__7721;
    wire N__7714;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7620;
    wire N__7615;
    wire N__7612;
    wire N__7611;
    wire N__7610;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7579;
    wire N__7578;
    wire N__7575;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7542;
    wire N__7539;
    wire N__7528;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7522;
    wire N__7521;
    wire N__7518;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7501;
    wire N__7498;
    wire N__7491;
    wire N__7486;
    wire N__7483;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7458;
    wire N__7457;
    wire N__7456;
    wire N__7453;
    wire N__7448;
    wire N__7445;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7399;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7391;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7362;
    wire N__7355;
    wire N__7352;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7289;
    wire N__7284;
    wire N__7281;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7260;
    wire N__7259;
    wire N__7258;
    wire N__7257;
    wire N__7252;
    wire N__7249;
    wire N__7244;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7221;
    wire N__7216;
    wire N__7213;
    wire N__7212;
    wire N__7211;
    wire N__7210;
    wire N__7209;
    wire N__7204;
    wire N__7201;
    wire N__7200;
    wire N__7195;
    wire N__7190;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7178;
    wire N__7171;
    wire N__7168;
    wire N__7167;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7111;
    wire N__7108;
    wire N__7107;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7041;
    wire N__7040;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7008;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__6999;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6979;
    wire N__6976;
    wire N__6975;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6958;
    wire N__6955;
    wire N__6954;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6935;
    wire N__6932;
    wire N__6925;
    wire N__6920;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6847;
    wire N__6844;
    wire N__6843;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6699;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6672;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6627;
    wire N__6626;
    wire N__6623;
    wire N__6618;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6507;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6449;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire \Clock50MHz.PixelClock ;
    wire GNDG0;
    wire VCCG0;
    wire font_un3_pixel_29_cascade_;
    wire Pixel_RNOZ0Z_18_cascade_;
    wire N_1214_0_cascade_;
    wire g1;
    wire bfn_1_4_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803;
    wire bfn_1_5_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO;
    wire charx_i_24;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3;
    wire charx_i_23;
    wire bfn_1_6_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7;
    wire un18_beamylto9_2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i;
    wire bfn_1_7_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8;
    wire bfn_1_8_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i;
    wire bfn_1_11_0_;
    wire un5_visiblex_cry_0;
    wire un5_visiblex_cry_1;
    wire un5_visiblex_cry_2;
    wire un5_visiblex_cry_3;
    wire un5_visiblex_cry_4;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire bfn_1_12_0_;
    wire un5_visiblex_cry_8;
    wire bfn_1_13_0_;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_1;
    wire charx_if_generate_plus_mult1_un26_sum_axb_3_i;
    wire g1_2_cascade_;
    wire g2_3_0_cascade_;
    wire g2_2_0;
    wire g3_3_cascade_;
    wire g0_0_2_cascade_;
    wire g0_3_cascade_;
    wire N_21_0;
    wire Pixel_RNOZ0Z_37;
    wire font_un126_pixel_m_2_1_1_cascade_;
    wire Pixel_RNOZ0Z_71;
    wire g0_0_1;
    wire font_un3_pixel_29;
    wire font_un126_pixel_m_2_1_cascade_;
    wire g2_2_0_1;
    wire charx_if_generate_plus_mult1_un1_sum_axb1_cascade_;
    wire font_un126_pixel_5_a0_2;
    wire G_19_i_a11_0_1_cascade_;
    wire Pixel_RNOZ0Z_36;
    wire g1_1_0_0_cascade_;
    wire g0_0;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0;
    wire bfn_2_6_0_;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2;
    wire charx_if_generate_plus_mult1_un68_sum_i_5;
    wire charx_if_generate_plus_mult1_un75_sum_cry_3;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1;
    wire charx_if_generate_plus_mult1_un68_sum_i;
    wire un13_beamylt7_0_cascade_;
    wire bfn_2_8_0_;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2;
    wire charx_if_generate_plus_mult1_un75_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_3;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0;
    wire charx_if_generate_plus_mult1_un61_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8;
    wire bfn_2_9_0_;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2;
    wire charx_if_generate_plus_mult1_un68_sum_axb_5;
    wire charx_if_generate_plus_mult1_un61_sum_cry_3;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_;
    wire charx_if_generate_plus_mult1_un61_sum_i_5;
    wire charx_if_generate_plus_mult1_un54_sum_i;
    wire bfn_2_10_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire beamXZ0Z_5;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire beamXZ0Z_8;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire beamXZ0Z_9;
    wire bfn_2_11_0_;
    wire un8_beamx_cry_9;
    wire beamXZ0Z_4;
    wire beamXZ0Z_6;
    wire un3_beamx_5;
    wire un3_beamx_7;
    wire beamXZ0Z_2;
    wire beamXZ0Z_3;
    wire un18_beamylt4;
    wire beamXZ0Z_1;
    wire bfn_2_12_0_;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538;
    wire charx_if_generate_plus_mult1_un33_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4;
    wire un5_visiblex_i_24;
    wire charx_if_generate_plus_mult1_un26_sum_i_5;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5;
    wire bfn_2_13_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7;
    wire g2_1_cascade_;
    wire N_7_cascade_;
    wire g2_1;
    wire g0_1_0_cascade_;
    wire g0_1_3_cascade_;
    wire g3_2_2_cascade_;
    wire N_20;
    wire g0_4_cascade_;
    wire G_21_i_2;
    wire Pixel_c;
    wire g1_1_0;
    wire g0_2_0;
    wire g1_1_cascade_;
    wire g3_1;
    wire g0_5;
    wire g1_0_0;
    wire g0_0_a3_0;
    wire beamXZ0Z_0;
    wire N_35;
    wire N_58_mux;
    wire charx_if_generate_plus_mult1_un1_sum_axb1;
    wire beamY_RNIDQG2Z0Z_0_cascade_;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3;
    wire beamY_RNINKIU27Z0Z_0;
    wire beamY_RNINKIU27Z0Z_0_cascade_;
    wire Pixel_RNOZ0Z_29_cascade_;
    wire N_10;
    wire chessboardpixel_un152_pixel_27;
    wire chessboardpixel_un174_pixellt10;
    wire chessboardpixel_un175_pixel;
    wire g1_2_1;
    wire chessboardpixel_un175_pixel_cascade_;
    wire g2_3_0_0;
    wire un13_beamylt7;
    wire un15_beamy;
    wire un18_beamylt10_0;
    wire un15_beamy_2;
    wire Pixel_RNOZ0Z_44_cascade_;
    wire N_10_0_0;
    wire beamXZ0Z_10;
    wire un1_beamx_2;
    wire beamXZ0Z_7;
    wire un1_beamxlt10_0;
    wire HSync_c;
    wire un4_row;
    wire bfn_4_8_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2;
    wire bfn_4_9_0_;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_axb_3_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum_c5_iZ0;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_2;
    wire if_generate_plus_mult1_un54_sum_axb_4_l_ofx;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum_i_5;
    wire un5_visiblex_i_26;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8;
    wire un4_row_9_2_cascade_;
    wire un4_row_9_5;
    wire un4_row_9_0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i;
    wire column_1_if_generate_plus_mult1_un47_sum_cZ0Z5;
    wire charx_if_generate_plus_mult1_un40_sum;
    wire bfn_4_11_0_;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_3;
    wire charx_if_generate_plus_mult1_un40_sum_axb_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_;
    wire charx_if_generate_plus_mult1_un33_sum;
    wire charx_if_generate_plus_mult1_un33_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum;
    wire bfn_4_12_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0;
    wire charx_if_generate_plus_mult1_un33_sum_i_5;
    wire charx_if_generate_plus_mult1_un26_sum_axb_3;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i;
    wire bfn_4_13_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8;
    wire Pixel_RNOZ0Z_14;
    wire font_un126_pixel_5_a0_1;
    wire N_1740_0;
    wire font_un28_pixel_29_cascade_;
    wire beamY_RNIDA2GGA3Z0Z_0;
    wire g0_1;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1;
    wire beamY_RNIDA2GGA3Z0Z_0_cascade_;
    wire N_19_0_0;
    wire font_un28_pixel_30;
    wire font_un28_pixel_29;
    wire N_15_i;
    wire Pixel_RNOZ0Z_28_cascade_;
    wire Pixel_RNOZ0Z_9;
    wire chary_24;
    wire chary_1_24_cascade_;
    wire N_1737_0;
    wire chary_1_0_24_cascade_;
    wire g2_3_cascade_;
    wire g1_1_1;
    wire un116_pixel_0_0_0;
    wire N_5_1;
    wire g0_0_a3_4;
    wire un8_beamylto9_1_cascade_;
    wire un8_beamy;
    wire N_134_0;
    wire g4_1;
    wire g0_0_a3_5;
    wire m4_rn_1_cascade_;
    wire Pixel_RNOZ0Z_40;
    wire content_content_ram0__RNIR1C2R81Z0Z_0_cascade_;
    wire N_331_i;
    wire un4_row_m7_ns_1_cascade_;
    wire beamY_RNIPAQ91Z0Z_6;
    wire un4_beamy_0;
    wire m4_sn;
    wire content_content_ram0__RNIR1C2R81_0Z0Z_0;
    wire un6_rowlt7_0;
    wire bfn_5_9_0_;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2;
    wire charx_if_generate_plus_mult1_un61_sum_axb_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_3;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7;
    wire charx_if_generate_plus_mult1_un47_sum_i;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6;
    wire charx_if_generate_plus_mult1_un47_sum;
    wire bfn_5_10_0_;
    wire charx_if_generate_plus_mult1_un40_sum_i;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2;
    wire charx_if_generate_plus_mult1_un40_sum_i_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1;
    wire charx_if_generate_plus_mult1_un54_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_3;
    wire charx_if_generate_plus_mult1_un47_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_;
    wire charx_if_generate_plus_mult1_un47_sum_i_5;
    wire bfn_5_11_0_;
    wire un5_visiblex_i_27;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_2;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_4;
    wire if_generate_plus_mult1_un61_sum_s_5_cascade_;
    wire charx_if_generate_plus_mult1_un54_sum;
    wire if_generate_plus_mult1_un54_sum_s_5;
    wire column_1_if_generate_plus_mult1_un54_sum_i_5;
    wire chary_2_24;
    wire beamY_RNI539IG9Z0Z_3;
    wire beamY_RNI539IG9Z0Z_3_cascade_;
    wire g4;
    wire chary_0_24;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_1;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_;
    wire g1_2_0;
    wire beamY_RNIMSO1N7_0Z0Z_2_cascade_;
    wire g4_0;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0;
    wire g2_1_0_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_0_5;
    wire Pixel_RNOZ0Z_66;
    wire un5_visibley_0_28;
    wire g2;
    wire un5_visibley_0_29;
    wire Pixel_RNOZ0Z_67;
    wire un4_beamylt6_cascade_;
    wire un4_beamylt8_0;
    wire GB_BUFFER_Clock12MHz_c_g_THRU_CO;
    wire charx_if_generate_plus_mult1_un75_sum;
    wire bfn_6_9_0_;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_1;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_2;
    wire G_383;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_4;
    wire un6_rowlto0;
    wire column_1_if_generate_plus_mult1_un75_sum_iZ0;
    wire charx_if_generate_plus_mult1_un68_sum;
    wire bfn_6_10_0_;
    wire if_generate_plus_mult1_un75_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_4;
    wire content_column_1_i_2_i_2;
    wire un6_rowlto1;
    wire content_N_25;
    wire bfn_6_11_0_;
    wire column_1_if_generate_plus_mult1_un61_sum_iZ0;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_1;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un61_sum_i_5;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_4;
    wire content_column_1_i_2_2_cascade_;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire if_generate_plus_mult1_un75_sum_axb_4_l_fx;
    wire chessboardpixel_un152_pixel_24;
    wire column_1_if_generate_plus_mult1_un68_sum_iZ0;
    wire content_m7_ns_1_cascade_;
    wire content_N_8;
    wire content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_;
    wire content_content_ram7__RNI6B0NG3Z0Z_0;
    wire content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_2_5;
    wire un5_visibley_2_29;
    wire g2_0_0;
    wire beamY_RNIMSO1N7Z0Z_2;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_1_0_5;
    wire g2_0;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1;
    wire g2_0_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_1_5;
    wire VSync_c;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3;
    wire un5_visibley_3_28;
    wire un5_visibley_3_28_cascade_;
    wire g1_3_cascade_;
    wire g2_0_1;
    wire un1_beamylto9_2;
    wire un5_visibley_1_28;
    wire chessboardpixel_un200_pixellto4_1_cascade_;
    wire chessboardpixel_un200_pixellt10;
    wire un8_beamy_3;
    wire beamY_i_2_cascade_;
    wire beamY_i_2;
    wire bfn_7_8_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0;
    wire chessboardpixel_un178_pixel_26;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0;
    wire row_1_if_generate_plus_mult1_un61_sum_cZ0Z5;
    wire row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3;
    wire if_generate_plus_mult1_un54_sum_axbxc5;
    wire row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0;
    wire content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_;
    wire content_content_ram9__e_0_RNIFBHPN1Z0Z_0;
    wire content_content_ram5__RNIEM2QF3Z0Z_0;
    wire content_ram9_0;
    wire content_ram11_0;
    wire nCS1_c;
    wire un5_visibley_2_28;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0;
    wire beamY_RNIVMI9D5Z0Z_3;
    wire un5_visibley_1_29;
    wire chary_if_generate_plus_mult1_un68_sum_c4;
    wire beamY_RNI8325Z0Z_6_cascade_;
    wire un5_visibley_c5_cascade_;
    wire un1_beamylto9_1;
    wire un5_visibley_c3_cascade_;
    wire un5_beamx_2_0_cascade_;
    wire un5_beamx_3;
    wire un5_visibley_ac0_11_0_1_cascade_;
    wire beamY_RNI8325_0Z0Z_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum;
    wire bfn_8_8_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0;
    wire bfn_8_9_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0;
    wire CO4_1;
    wire row_1_if_generate_plus_mult1_un47_sum_cZ0Z5;
    wire content_ram8_0;
    wire content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_;
    wire content_N_19;
    wire content_column_1_i_2_2;
    wire if_generate_plus_mult1_un61_sum_s_5;
    wire content_content_ram10__e_0_RNIOLNMN1Z0Z_0;
    wire content_ram3_0;
    wire content_awe9;
    wire content_ram0_0;
    wire content_awe8;
    wire content_awe11;
    wire content_ram5_0;
    wire content_ram12_0;
    wire content_awe0_0_a2_0;
    wire content_awe0_0_a2_0_cascade_;
    wire content_ram4_0;
    wire content_N_36;
    wire content_N_36_cascade_;
    wire content_awe7_1_cascade_;
    wire content_ram6_0;
    wire content_awe7_1;
    wire content_ram7_0;
    wire nCS1_0_sqmuxa;
    wire un19_slaveselectlt5_0_cascade_;
    wire un19_slaveselectlt5_0;
    wire counter_RNI4HQB1Z0Z_5_cascade_;
    wire beamY_RNI4FVGVZ0Z_4_cascade_;
    wire chary_if_generate_plus_mult1_un75_sum_c5;
    wire N_596_2;
    wire un5_visibley_4_28_cascade_;
    wire un5_visibley_3_29;
    wire g1_8_1_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_i;
    wire g1_3_0;
    wire un5_visibley_1_0_28;
    wire beamY_RNIJ0H2Z0Z_4_cascade_;
    wire un5_visibley_c5;
    wire un5_visibley_c6_0_0_0;
    wire un5_visibley_c6_0_0_0_cascade_;
    wire un5_visibley_c3;
    wire beamYZ0Z_1;
    wire beamYZ0Z_0;
    wire g2_1_1_0;
    wire bfn_9_7_0_;
    wire beamYZ0Z_2;
    wire un21_beamy_cry_1;
    wire beamYZ0Z_3;
    wire un21_beamy_cry_2;
    wire beamYZ0Z_4;
    wire un21_beamy_cry_3;
    wire beamYZ0Z_5;
    wire un21_beamy_cry_4;
    wire beamYZ0Z_6;
    wire un21_beamy_cry_5;
    wire beamYZ0Z_7;
    wire un21_beamy_cry_6;
    wire beamYZ0Z_8;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire beamY_RNI9DLCZ0Z_1;
    wire bfn_9_8_0_;
    wire beamYZ0Z_9;
    wire PixelClock_g;
    wire beamX_RNI5457Z0Z_5;
    wire bfn_9_9_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0;
    wire bfn_9_10_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0;
    wire content_ram10_0;
    wire content_awe10;
    wire content_N_35_cascade_;
    wire content_awe3_1;
    wire content_awe3_1_cascade_;
    wire content_ram2_0;
    wire content_N_40;
    wire content_N_35;
    wire content_awe1_0_a2_0_cascade_;
    wire content_ram1_0;
    wire un7_slaveselectlt5_cascade_;
    wire N_190_i;
    wire un1_counter_0_1;
    wire un7_slaveselectlt5;
    wire un1_counter_0_1_cascade_;
    wire slaveselect_1lto5_0_cascade_;
    wire slaveselect_1lto5_1;
    wire SCLK1_0_i;
    wire counterZ0Z_1;
    wire counterZ0Z_0;
    wire un7_slaveselectlt2_0;
    wire bfn_9_14_0_;
    wire counterZ0Z_2;
    wire counter_cry_1;
    wire counterZ0Z_3;
    wire counter_cry_2;
    wire counterZ0Z_4;
    wire counter_cry_3;
    wire counter_RNI4HQB1Z0Z_5;
    wire counter_cry_4;
    wire counterZ0Z_5;
    wire SDATA1_c;
    wire slaveselectZ0;
    wire un5_slaveselect;
    wire SDATA2_c;
    wire Clock12MHz_c_g;
    wire chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_;
    wire beamY_RNII78UPZ0Z_4;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_c5;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0;
    wire chary_if_generate_plus_mult1_un61_sum_c5_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_axbxc5_0;
    wire chary_if_generate_plus_mult1_un61_sum_c4;
    wire chary_if_generate_plus_mult1_un47_sum_axb3;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_1;
    wire chary_if_generate_plus_mult1_un54_sum_c5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum;
    wire beamY_RNIFC5HAZ0Z_4;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1;
    wire chary_if_generate_plus_mult1_un47_sum_ac0_8;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_2;
    wire chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_;
    wire chary_if_generate_plus_mult1_un47_sum_axb4;
    wire beamY_RNI65RM4_0Z0Z_9;
    wire beamY_RNIJNLCZ0Z_9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum;
    wire chary_if_generate_plus_mult1_un47_sum_c4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0;
    wire bfn_11_8_0_;
    wire beamY_RNIQ7DB_0Z0Z_9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire chary_if_generate_plus_mult1_un33_sum_axb3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum;
    wire bfn_11_9_0_;
    wire beamY_RNITSR8_0Z0Z_8;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0;
    wire CONSTANT_ONE_NET;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__10363),
            .RESETB(N__15601),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF Clock12MHz_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__15818),
            .GLOBALBUFFEROUTPUT(Clock12MHz_c_g));
    defparam Clock12MHz_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_gb_io_iopad (
            .OE(N__15820),
            .DIN(N__15819),
            .DOUT(N__15818),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_gb_io_preio (
            .PADOEN(N__15820),
            .PADOUT(N__15819),
            .PADIN(N__15818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__15809),
            .DIN(N__15808),
            .DOUT(N__15807),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__15809),
            .PADOUT(N__15808),
            .PADIN(N__15807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10753),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__15800),
            .DIN(N__15799),
            .DOUT(N__15798),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__15800),
            .PADOUT(N__15799),
            .PADIN(N__15798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8353),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SDATA2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SDATA2_obuf_iopad (
            .OE(N__15791),
            .DIN(N__15790),
            .DOUT(N__15789),
            .PACKAGEPIN(SDATA2));
    defparam SDATA2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SDATA2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SDATA2_obuf_preio (
            .PADOEN(N__15791),
            .PADOUT(N__15790),
            .PADIN(N__15789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14374),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS1_obuf_iopad (
            .OE(N__15782),
            .DIN(N__15781),
            .DOUT(N__15780),
            .PACKAGEPIN(nCS1));
    defparam nCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS1_obuf_preio (
            .PADOEN(N__15782),
            .PADOUT(N__15781),
            .PADIN(N__15780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__15773),
            .DIN(N__15772),
            .DOUT(N__15771),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__15773),
            .PADOUT(N__15772),
            .PADIN(N__15771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8035),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK1_obuf_iopad (
            .OE(N__15764),
            .DIN(N__15763),
            .DOUT(N__15762),
            .PACKAGEPIN(SCLK1));
    defparam SCLK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCLK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCLK1_obuf_preio (
            .PADOEN(N__15764),
            .PADOUT(N__15763),
            .PADIN(N__15762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK2_obuf_iopad (
            .OE(N__15755),
            .DIN(N__15754),
            .DOUT(N__15753),
            .PACKAGEPIN(SCLK2));
    defparam SCLK2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCLK2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCLK2_obuf_preio (
            .PADOEN(N__15755),
            .PADOUT(N__15754),
            .PADIN(N__15753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14133),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS2_obuf_iopad (
            .OE(N__15746),
            .DIN(N__15745),
            .DOUT(N__15744),
            .PACKAGEPIN(nCS2));
    defparam nCS2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS2_obuf_preio (
            .PADOEN(N__15746),
            .PADOUT(N__15745),
            .PADIN(N__15744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SDATA1_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SDATA1_ibuf_iopad (
            .OE(N__15737),
            .DIN(N__15736),
            .DOUT(N__15735),
            .PACKAGEPIN(SDATA1));
    defparam SDATA1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SDATA1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SDATA1_ibuf_preio (
            .PADOEN(N__15737),
            .PADOUT(N__15736),
            .PADIN(N__15735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SDATA1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3653 (
            .O(N__15718),
            .I(N__15713));
    InMux I__3652 (
            .O(N__15717),
            .I(N__15710));
    InMux I__3651 (
            .O(N__15716),
            .I(N__15701));
    LocalMux I__3650 (
            .O(N__15713),
            .I(N__15696));
    LocalMux I__3649 (
            .O(N__15710),
            .I(N__15696));
    InMux I__3648 (
            .O(N__15709),
            .I(N__15693));
    InMux I__3647 (
            .O(N__15708),
            .I(N__15690));
    InMux I__3646 (
            .O(N__15707),
            .I(N__15683));
    InMux I__3645 (
            .O(N__15706),
            .I(N__15683));
    InMux I__3644 (
            .O(N__15705),
            .I(N__15683));
    InMux I__3643 (
            .O(N__15704),
            .I(N__15680));
    LocalMux I__3642 (
            .O(N__15701),
            .I(N__15677));
    Span4Mux_v I__3641 (
            .O(N__15696),
            .I(N__15672));
    LocalMux I__3640 (
            .O(N__15693),
            .I(N__15672));
    LocalMux I__3639 (
            .O(N__15690),
            .I(N__15667));
    LocalMux I__3638 (
            .O(N__15683),
            .I(N__15667));
    LocalMux I__3637 (
            .O(N__15680),
            .I(N__15662));
    Span4Mux_s3_h I__3636 (
            .O(N__15677),
            .I(N__15662));
    Odrv4 I__3635 (
            .O(N__15672),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3634 (
            .O(N__15667),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3633 (
            .O(N__15662),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    InMux I__3632 (
            .O(N__15655),
            .I(N__15652));
    LocalMux I__3631 (
            .O(N__15652),
            .I(beamY_RNITSR8_0Z0Z_8));
    CascadeMux I__3630 (
            .O(N__15649),
            .I(N__15646));
    InMux I__3629 (
            .O(N__15646),
            .I(N__15643));
    LocalMux I__3628 (
            .O(N__15643),
            .I(N__15640));
    Odrv4 I__3627 (
            .O(N__15640),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0));
    InMux I__3626 (
            .O(N__15637),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__3625 (
            .O(N__15634),
            .I(N__15631));
    InMux I__3624 (
            .O(N__15631),
            .I(N__15628));
    LocalMux I__3623 (
            .O(N__15628),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0));
    InMux I__3622 (
            .O(N__15625),
            .I(N__15622));
    LocalMux I__3621 (
            .O(N__15622),
            .I(N__15619));
    Odrv12 I__3620 (
            .O(N__15619),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0));
    InMux I__3619 (
            .O(N__15616),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__3618 (
            .O(N__15613),
            .I(N__15610));
    LocalMux I__3617 (
            .O(N__15610),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0));
    CascadeMux I__3616 (
            .O(N__15607),
            .I(N__15603));
    InMux I__3615 (
            .O(N__15606),
            .I(N__15593));
    InMux I__3614 (
            .O(N__15603),
            .I(N__15588));
    InMux I__3613 (
            .O(N__15602),
            .I(N__15588));
    IoInMux I__3612 (
            .O(N__15601),
            .I(N__15582));
    InMux I__3611 (
            .O(N__15600),
            .I(N__15579));
    CascadeMux I__3610 (
            .O(N__15599),
            .I(N__15576));
    CascadeMux I__3609 (
            .O(N__15598),
            .I(N__15572));
    CascadeMux I__3608 (
            .O(N__15597),
            .I(N__15569));
    CascadeMux I__3607 (
            .O(N__15596),
            .I(N__15566));
    LocalMux I__3606 (
            .O(N__15593),
            .I(N__15561));
    LocalMux I__3605 (
            .O(N__15588),
            .I(N__15561));
    CascadeMux I__3604 (
            .O(N__15587),
            .I(N__15558));
    CascadeMux I__3603 (
            .O(N__15586),
            .I(N__15555));
    CascadeMux I__3602 (
            .O(N__15585),
            .I(N__15552));
    LocalMux I__3601 (
            .O(N__15582),
            .I(N__15547));
    LocalMux I__3600 (
            .O(N__15579),
            .I(N__15544));
    InMux I__3599 (
            .O(N__15576),
            .I(N__15537));
    InMux I__3598 (
            .O(N__15575),
            .I(N__15537));
    InMux I__3597 (
            .O(N__15572),
            .I(N__15537));
    InMux I__3596 (
            .O(N__15569),
            .I(N__15534));
    InMux I__3595 (
            .O(N__15566),
            .I(N__15531));
    Span4Mux_h I__3594 (
            .O(N__15561),
            .I(N__15528));
    InMux I__3593 (
            .O(N__15558),
            .I(N__15525));
    InMux I__3592 (
            .O(N__15555),
            .I(N__15522));
    InMux I__3591 (
            .O(N__15552),
            .I(N__15519));
    CascadeMux I__3590 (
            .O(N__15551),
            .I(N__15516));
    CascadeMux I__3589 (
            .O(N__15550),
            .I(N__15513));
    Span4Mux_s3_v I__3588 (
            .O(N__15547),
            .I(N__15510));
    Span4Mux_v I__3587 (
            .O(N__15544),
            .I(N__15507));
    LocalMux I__3586 (
            .O(N__15537),
            .I(N__15504));
    LocalMux I__3585 (
            .O(N__15534),
            .I(N__15493));
    LocalMux I__3584 (
            .O(N__15531),
            .I(N__15493));
    Sp12to4 I__3583 (
            .O(N__15528),
            .I(N__15493));
    LocalMux I__3582 (
            .O(N__15525),
            .I(N__15493));
    LocalMux I__3581 (
            .O(N__15522),
            .I(N__15493));
    LocalMux I__3580 (
            .O(N__15519),
            .I(N__15490));
    InMux I__3579 (
            .O(N__15516),
            .I(N__15487));
    InMux I__3578 (
            .O(N__15513),
            .I(N__15484));
    Span4Mux_h I__3577 (
            .O(N__15510),
            .I(N__15480));
    Span4Mux_v I__3576 (
            .O(N__15507),
            .I(N__15477));
    Span12Mux_s6_h I__3575 (
            .O(N__15504),
            .I(N__15474));
    Span12Mux_s8_v I__3574 (
            .O(N__15493),
            .I(N__15465));
    Span12Mux_s7_v I__3573 (
            .O(N__15490),
            .I(N__15465));
    LocalMux I__3572 (
            .O(N__15487),
            .I(N__15465));
    LocalMux I__3571 (
            .O(N__15484),
            .I(N__15465));
    InMux I__3570 (
            .O(N__15483),
            .I(N__15462));
    Odrv4 I__3569 (
            .O(N__15480),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3568 (
            .O(N__15477),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3567 (
            .O(N__15474),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3566 (
            .O(N__15465),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3565 (
            .O(N__15462),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__3564 (
            .O(N__15451),
            .I(N__15448));
    InMux I__3563 (
            .O(N__15448),
            .I(N__15445));
    LocalMux I__3562 (
            .O(N__15445),
            .I(N__15442));
    Odrv4 I__3561 (
            .O(N__15442),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0));
    InMux I__3560 (
            .O(N__15439),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__3559 (
            .O(N__15436),
            .I(N__15433));
    InMux I__3558 (
            .O(N__15433),
            .I(N__15430));
    LocalMux I__3557 (
            .O(N__15430),
            .I(N__15427));
    Odrv4 I__3556 (
            .O(N__15427),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__3555 (
            .O(N__15424),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__3554 (
            .O(N__15421),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__3553 (
            .O(N__15418),
            .I(N__15413));
    CascadeMux I__3552 (
            .O(N__15417),
            .I(N__15409));
    InMux I__3551 (
            .O(N__15416),
            .I(N__15397));
    InMux I__3550 (
            .O(N__15413),
            .I(N__15397));
    InMux I__3549 (
            .O(N__15412),
            .I(N__15397));
    InMux I__3548 (
            .O(N__15409),
            .I(N__15397));
    InMux I__3547 (
            .O(N__15408),
            .I(N__15397));
    LocalMux I__3546 (
            .O(N__15397),
            .I(N__15394));
    Odrv4 I__3545 (
            .O(N__15394),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9));
    InMux I__3544 (
            .O(N__15391),
            .I(N__15385));
    InMux I__3543 (
            .O(N__15390),
            .I(N__15385));
    LocalMux I__3542 (
            .O(N__15385),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__3541 (
            .O(N__15382),
            .I(N__15379));
    LocalMux I__3540 (
            .O(N__15379),
            .I(N__15374));
    InMux I__3539 (
            .O(N__15378),
            .I(N__15369));
    InMux I__3538 (
            .O(N__15377),
            .I(N__15369));
    Odrv4 I__3537 (
            .O(N__15374),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__3536 (
            .O(N__15369),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    InMux I__3535 (
            .O(N__15364),
            .I(N__15358));
    InMux I__3534 (
            .O(N__15363),
            .I(N__15358));
    LocalMux I__3533 (
            .O(N__15358),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_2));
    CascadeMux I__3532 (
            .O(N__15355),
            .I(chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_));
    InMux I__3531 (
            .O(N__15352),
            .I(N__15346));
    InMux I__3530 (
            .O(N__15351),
            .I(N__15346));
    LocalMux I__3529 (
            .O(N__15346),
            .I(chary_if_generate_plus_mult1_un47_sum_axb4));
    InMux I__3528 (
            .O(N__15343),
            .I(N__15337));
    InMux I__3527 (
            .O(N__15342),
            .I(N__15337));
    LocalMux I__3526 (
            .O(N__15337),
            .I(N__15332));
    InMux I__3525 (
            .O(N__15336),
            .I(N__15327));
    InMux I__3524 (
            .O(N__15335),
            .I(N__15327));
    Odrv4 I__3523 (
            .O(N__15332),
            .I(beamY_RNI65RM4_0Z0Z_9));
    LocalMux I__3522 (
            .O(N__15327),
            .I(beamY_RNI65RM4_0Z0Z_9));
    CascadeMux I__3521 (
            .O(N__15322),
            .I(N__15316));
    CascadeMux I__3520 (
            .O(N__15321),
            .I(N__15313));
    InMux I__3519 (
            .O(N__15320),
            .I(N__15304));
    InMux I__3518 (
            .O(N__15319),
            .I(N__15304));
    InMux I__3517 (
            .O(N__15316),
            .I(N__15304));
    InMux I__3516 (
            .O(N__15313),
            .I(N__15304));
    LocalMux I__3515 (
            .O(N__15304),
            .I(N__15301));
    Span4Mux_s3_h I__3514 (
            .O(N__15301),
            .I(N__15298));
    Odrv4 I__3513 (
            .O(N__15298),
            .I(beamY_RNIJNLCZ0Z_9));
    CascadeMux I__3512 (
            .O(N__15295),
            .I(N__15286));
    InMux I__3511 (
            .O(N__15294),
            .I(N__15281));
    InMux I__3510 (
            .O(N__15293),
            .I(N__15281));
    InMux I__3509 (
            .O(N__15292),
            .I(N__15275));
    InMux I__3508 (
            .O(N__15291),
            .I(N__15275));
    InMux I__3507 (
            .O(N__15290),
            .I(N__15268));
    InMux I__3506 (
            .O(N__15289),
            .I(N__15268));
    InMux I__3505 (
            .O(N__15286),
            .I(N__15265));
    LocalMux I__3504 (
            .O(N__15281),
            .I(N__15262));
    InMux I__3503 (
            .O(N__15280),
            .I(N__15259));
    LocalMux I__3502 (
            .O(N__15275),
            .I(N__15256));
    InMux I__3501 (
            .O(N__15274),
            .I(N__15253));
    InMux I__3500 (
            .O(N__15273),
            .I(N__15250));
    LocalMux I__3499 (
            .O(N__15268),
            .I(N__15245));
    LocalMux I__3498 (
            .O(N__15265),
            .I(N__15245));
    Span4Mux_s3_h I__3497 (
            .O(N__15262),
            .I(N__15242));
    LocalMux I__3496 (
            .O(N__15259),
            .I(N__15239));
    Span4Mux_s3_h I__3495 (
            .O(N__15256),
            .I(N__15232));
    LocalMux I__3494 (
            .O(N__15253),
            .I(N__15232));
    LocalMux I__3493 (
            .O(N__15250),
            .I(N__15232));
    Odrv4 I__3492 (
            .O(N__15245),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3491 (
            .O(N__15242),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv12 I__3490 (
            .O(N__15239),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3489 (
            .O(N__15232),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    InMux I__3488 (
            .O(N__15223),
            .I(N__15217));
    InMux I__3487 (
            .O(N__15222),
            .I(N__15217));
    LocalMux I__3486 (
            .O(N__15217),
            .I(chary_if_generate_plus_mult1_un47_sum_c4));
    InMux I__3485 (
            .O(N__15214),
            .I(N__15211));
    LocalMux I__3484 (
            .O(N__15211),
            .I(N__15208));
    Span4Mux_s2_h I__3483 (
            .O(N__15208),
            .I(N__15205));
    Odrv4 I__3482 (
            .O(N__15205),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0));
    InMux I__3481 (
            .O(N__15202),
            .I(N__15199));
    LocalMux I__3480 (
            .O(N__15199),
            .I(beamY_RNIQ7DB_0Z0Z_9));
    InMux I__3479 (
            .O(N__15196),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__3478 (
            .O(N__15193),
            .I(N__15185));
    CascadeMux I__3477 (
            .O(N__15192),
            .I(N__15182));
    InMux I__3476 (
            .O(N__15191),
            .I(N__15176));
    InMux I__3475 (
            .O(N__15190),
            .I(N__15173));
    InMux I__3474 (
            .O(N__15189),
            .I(N__15168));
    InMux I__3473 (
            .O(N__15188),
            .I(N__15168));
    LocalMux I__3472 (
            .O(N__15185),
            .I(N__15165));
    InMux I__3471 (
            .O(N__15182),
            .I(N__15162));
    InMux I__3470 (
            .O(N__15181),
            .I(N__15155));
    InMux I__3469 (
            .O(N__15180),
            .I(N__15155));
    InMux I__3468 (
            .O(N__15179),
            .I(N__15155));
    LocalMux I__3467 (
            .O(N__15176),
            .I(N__15148));
    LocalMux I__3466 (
            .O(N__15173),
            .I(N__15148));
    LocalMux I__3465 (
            .O(N__15168),
            .I(N__15148));
    Span4Mux_s3_h I__3464 (
            .O(N__15165),
            .I(N__15145));
    LocalMux I__3463 (
            .O(N__15162),
            .I(N__15140));
    LocalMux I__3462 (
            .O(N__15155),
            .I(N__15140));
    Odrv4 I__3461 (
            .O(N__15148),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__3460 (
            .O(N__15145),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv12 I__3459 (
            .O(N__15140),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    InMux I__3458 (
            .O(N__15133),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__3457 (
            .O(N__15130),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5));
    CascadeMux I__3456 (
            .O(N__15127),
            .I(N__15124));
    InMux I__3455 (
            .O(N__15124),
            .I(N__15116));
    InMux I__3454 (
            .O(N__15123),
            .I(N__15116));
    InMux I__3453 (
            .O(N__15122),
            .I(N__15109));
    InMux I__3452 (
            .O(N__15121),
            .I(N__15106));
    LocalMux I__3451 (
            .O(N__15116),
            .I(N__15103));
    InMux I__3450 (
            .O(N__15115),
            .I(N__15096));
    InMux I__3449 (
            .O(N__15114),
            .I(N__15096));
    InMux I__3448 (
            .O(N__15113),
            .I(N__15096));
    InMux I__3447 (
            .O(N__15112),
            .I(N__15093));
    LocalMux I__3446 (
            .O(N__15109),
            .I(N__15088));
    LocalMux I__3445 (
            .O(N__15106),
            .I(N__15088));
    Span4Mux_h I__3444 (
            .O(N__15103),
            .I(N__15083));
    LocalMux I__3443 (
            .O(N__15096),
            .I(N__15083));
    LocalMux I__3442 (
            .O(N__15093),
            .I(N__15080));
    Span4Mux_v I__3441 (
            .O(N__15088),
            .I(N__15075));
    Span4Mux_v I__3440 (
            .O(N__15083),
            .I(N__15075));
    Span4Mux_s2_h I__3439 (
            .O(N__15080),
            .I(N__15072));
    Odrv4 I__3438 (
            .O(N__15075),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__3437 (
            .O(N__15072),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    InMux I__3436 (
            .O(N__15067),
            .I(N__15064));
    LocalMux I__3435 (
            .O(N__15064),
            .I(N__15060));
    InMux I__3434 (
            .O(N__15063),
            .I(N__15053));
    Span4Mux_h I__3433 (
            .O(N__15060),
            .I(N__15049));
    InMux I__3432 (
            .O(N__15059),
            .I(N__15044));
    InMux I__3431 (
            .O(N__15058),
            .I(N__15044));
    InMux I__3430 (
            .O(N__15057),
            .I(N__15039));
    InMux I__3429 (
            .O(N__15056),
            .I(N__15039));
    LocalMux I__3428 (
            .O(N__15053),
            .I(N__15036));
    InMux I__3427 (
            .O(N__15052),
            .I(N__15033));
    Span4Mux_h I__3426 (
            .O(N__15049),
            .I(N__15030));
    LocalMux I__3425 (
            .O(N__15044),
            .I(N__15025));
    LocalMux I__3424 (
            .O(N__15039),
            .I(N__15025));
    Span4Mux_v I__3423 (
            .O(N__15036),
            .I(N__15020));
    LocalMux I__3422 (
            .O(N__15033),
            .I(N__15020));
    Odrv4 I__3421 (
            .O(N__15030),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv12 I__3420 (
            .O(N__15025),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    Odrv4 I__3419 (
            .O(N__15020),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    InMux I__3418 (
            .O(N__15013),
            .I(N__15010));
    LocalMux I__3417 (
            .O(N__15010),
            .I(chary_if_generate_plus_mult1_un61_sum_c4));
    CascadeMux I__3416 (
            .O(N__15007),
            .I(N__15003));
    CascadeMux I__3415 (
            .O(N__15006),
            .I(N__15000));
    InMux I__3414 (
            .O(N__15003),
            .I(N__14995));
    InMux I__3413 (
            .O(N__15000),
            .I(N__14995));
    LocalMux I__3412 (
            .O(N__14995),
            .I(N__14992));
    Odrv4 I__3411 (
            .O(N__14992),
            .I(chary_if_generate_plus_mult1_un47_sum_axb3));
    CascadeMux I__3410 (
            .O(N__14989),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_));
    CascadeMux I__3409 (
            .O(N__14986),
            .I(N__14978));
    CascadeMux I__3408 (
            .O(N__14985),
            .I(N__14975));
    CascadeMux I__3407 (
            .O(N__14984),
            .I(N__14971));
    CascadeMux I__3406 (
            .O(N__14983),
            .I(N__14968));
    InMux I__3405 (
            .O(N__14982),
            .I(N__14959));
    InMux I__3404 (
            .O(N__14981),
            .I(N__14959));
    InMux I__3403 (
            .O(N__14978),
            .I(N__14959));
    InMux I__3402 (
            .O(N__14975),
            .I(N__14954));
    InMux I__3401 (
            .O(N__14974),
            .I(N__14954));
    InMux I__3400 (
            .O(N__14971),
            .I(N__14943));
    InMux I__3399 (
            .O(N__14968),
            .I(N__14943));
    InMux I__3398 (
            .O(N__14967),
            .I(N__14940));
    InMux I__3397 (
            .O(N__14966),
            .I(N__14937));
    LocalMux I__3396 (
            .O(N__14959),
            .I(N__14932));
    LocalMux I__3395 (
            .O(N__14954),
            .I(N__14932));
    InMux I__3394 (
            .O(N__14953),
            .I(N__14923));
    InMux I__3393 (
            .O(N__14952),
            .I(N__14923));
    InMux I__3392 (
            .O(N__14951),
            .I(N__14923));
    InMux I__3391 (
            .O(N__14950),
            .I(N__14923));
    InMux I__3390 (
            .O(N__14949),
            .I(N__14918));
    InMux I__3389 (
            .O(N__14948),
            .I(N__14918));
    LocalMux I__3388 (
            .O(N__14943),
            .I(N__14914));
    LocalMux I__3387 (
            .O(N__14940),
            .I(N__14911));
    LocalMux I__3386 (
            .O(N__14937),
            .I(N__14904));
    Span4Mux_h I__3385 (
            .O(N__14932),
            .I(N__14904));
    LocalMux I__3384 (
            .O(N__14923),
            .I(N__14904));
    LocalMux I__3383 (
            .O(N__14918),
            .I(N__14901));
    InMux I__3382 (
            .O(N__14917),
            .I(N__14898));
    Span4Mux_h I__3381 (
            .O(N__14914),
            .I(N__14893));
    Span4Mux_h I__3380 (
            .O(N__14911),
            .I(N__14893));
    Span4Mux_h I__3379 (
            .O(N__14904),
            .I(N__14890));
    Odrv12 I__3378 (
            .O(N__14901),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    LocalMux I__3377 (
            .O(N__14898),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    Odrv4 I__3376 (
            .O(N__14893),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    Odrv4 I__3375 (
            .O(N__14890),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    CascadeMux I__3374 (
            .O(N__14881),
            .I(N__14876));
    InMux I__3373 (
            .O(N__14880),
            .I(N__14868));
    InMux I__3372 (
            .O(N__14879),
            .I(N__14868));
    InMux I__3371 (
            .O(N__14876),
            .I(N__14861));
    InMux I__3370 (
            .O(N__14875),
            .I(N__14861));
    InMux I__3369 (
            .O(N__14874),
            .I(N__14861));
    InMux I__3368 (
            .O(N__14873),
            .I(N__14858));
    LocalMux I__3367 (
            .O(N__14868),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__3366 (
            .O(N__14861),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__3365 (
            .O(N__14858),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    InMux I__3364 (
            .O(N__14851),
            .I(N__14843));
    InMux I__3363 (
            .O(N__14850),
            .I(N__14836));
    InMux I__3362 (
            .O(N__14849),
            .I(N__14836));
    InMux I__3361 (
            .O(N__14848),
            .I(N__14836));
    InMux I__3360 (
            .O(N__14847),
            .I(N__14832));
    CascadeMux I__3359 (
            .O(N__14846),
            .I(N__14829));
    LocalMux I__3358 (
            .O(N__14843),
            .I(N__14822));
    LocalMux I__3357 (
            .O(N__14836),
            .I(N__14822));
    InMux I__3356 (
            .O(N__14835),
            .I(N__14819));
    LocalMux I__3355 (
            .O(N__14832),
            .I(N__14816));
    InMux I__3354 (
            .O(N__14829),
            .I(N__14811));
    InMux I__3353 (
            .O(N__14828),
            .I(N__14811));
    InMux I__3352 (
            .O(N__14827),
            .I(N__14808));
    Span4Mux_v I__3351 (
            .O(N__14822),
            .I(N__14805));
    LocalMux I__3350 (
            .O(N__14819),
            .I(N__14800));
    Span4Mux_v I__3349 (
            .O(N__14816),
            .I(N__14800));
    LocalMux I__3348 (
            .O(N__14811),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    LocalMux I__3347 (
            .O(N__14808),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__3346 (
            .O(N__14805),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__3345 (
            .O(N__14800),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    InMux I__3344 (
            .O(N__14791),
            .I(N__14777));
    InMux I__3343 (
            .O(N__14790),
            .I(N__14777));
    InMux I__3342 (
            .O(N__14789),
            .I(N__14770));
    InMux I__3341 (
            .O(N__14788),
            .I(N__14770));
    InMux I__3340 (
            .O(N__14787),
            .I(N__14770));
    InMux I__3339 (
            .O(N__14786),
            .I(N__14766));
    InMux I__3338 (
            .O(N__14785),
            .I(N__14757));
    InMux I__3337 (
            .O(N__14784),
            .I(N__14757));
    InMux I__3336 (
            .O(N__14783),
            .I(N__14757));
    InMux I__3335 (
            .O(N__14782),
            .I(N__14757));
    LocalMux I__3334 (
            .O(N__14777),
            .I(N__14754));
    LocalMux I__3333 (
            .O(N__14770),
            .I(N__14751));
    InMux I__3332 (
            .O(N__14769),
            .I(N__14748));
    LocalMux I__3331 (
            .O(N__14766),
            .I(N__14742));
    LocalMux I__3330 (
            .O(N__14757),
            .I(N__14742));
    Span4Mux_h I__3329 (
            .O(N__14754),
            .I(N__14735));
    Span4Mux_s3_h I__3328 (
            .O(N__14751),
            .I(N__14735));
    LocalMux I__3327 (
            .O(N__14748),
            .I(N__14735));
    InMux I__3326 (
            .O(N__14747),
            .I(N__14732));
    Span4Mux_s2_h I__3325 (
            .O(N__14742),
            .I(N__14729));
    Sp12to4 I__3324 (
            .O(N__14735),
            .I(N__14724));
    LocalMux I__3323 (
            .O(N__14732),
            .I(N__14724));
    Odrv4 I__3322 (
            .O(N__14729),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__3321 (
            .O(N__14724),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    InMux I__3320 (
            .O(N__14719),
            .I(N__14712));
    InMux I__3319 (
            .O(N__14718),
            .I(N__14709));
    InMux I__3318 (
            .O(N__14717),
            .I(N__14706));
    CascadeMux I__3317 (
            .O(N__14716),
            .I(N__14699));
    CascadeMux I__3316 (
            .O(N__14715),
            .I(N__14696));
    LocalMux I__3315 (
            .O(N__14712),
            .I(N__14693));
    LocalMux I__3314 (
            .O(N__14709),
            .I(N__14690));
    LocalMux I__3313 (
            .O(N__14706),
            .I(N__14687));
    InMux I__3312 (
            .O(N__14705),
            .I(N__14682));
    InMux I__3311 (
            .O(N__14704),
            .I(N__14682));
    InMux I__3310 (
            .O(N__14703),
            .I(N__14677));
    InMux I__3309 (
            .O(N__14702),
            .I(N__14677));
    InMux I__3308 (
            .O(N__14699),
            .I(N__14672));
    InMux I__3307 (
            .O(N__14696),
            .I(N__14672));
    Span4Mux_v I__3306 (
            .O(N__14693),
            .I(N__14659));
    Span4Mux_h I__3305 (
            .O(N__14690),
            .I(N__14659));
    Span4Mux_v I__3304 (
            .O(N__14687),
            .I(N__14659));
    LocalMux I__3303 (
            .O(N__14682),
            .I(N__14659));
    LocalMux I__3302 (
            .O(N__14677),
            .I(N__14659));
    LocalMux I__3301 (
            .O(N__14672),
            .I(N__14659));
    Span4Mux_h I__3300 (
            .O(N__14659),
            .I(N__14656));
    Odrv4 I__3299 (
            .O(N__14656),
            .I(beamY_RNIFC5HAZ0Z_4));
    CascadeMux I__3298 (
            .O(N__14653),
            .I(N__14647));
    CascadeMux I__3297 (
            .O(N__14652),
            .I(N__14643));
    InMux I__3296 (
            .O(N__14651),
            .I(N__14633));
    InMux I__3295 (
            .O(N__14650),
            .I(N__14633));
    InMux I__3294 (
            .O(N__14647),
            .I(N__14633));
    InMux I__3293 (
            .O(N__14646),
            .I(N__14633));
    InMux I__3292 (
            .O(N__14643),
            .I(N__14628));
    InMux I__3291 (
            .O(N__14642),
            .I(N__14628));
    LocalMux I__3290 (
            .O(N__14633),
            .I(N__14625));
    LocalMux I__3289 (
            .O(N__14628),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    Odrv4 I__3288 (
            .O(N__14625),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    CascadeMux I__3287 (
            .O(N__14620),
            .I(N__14617));
    InMux I__3286 (
            .O(N__14617),
            .I(N__14614));
    LocalMux I__3285 (
            .O(N__14614),
            .I(chary_if_generate_plus_mult1_un47_sum_ac0_8));
    InMux I__3284 (
            .O(N__14611),
            .I(N__14601));
    InMux I__3283 (
            .O(N__14610),
            .I(N__14601));
    InMux I__3282 (
            .O(N__14609),
            .I(N__14596));
    InMux I__3281 (
            .O(N__14608),
            .I(N__14596));
    InMux I__3280 (
            .O(N__14607),
            .I(N__14591));
    InMux I__3279 (
            .O(N__14606),
            .I(N__14591));
    LocalMux I__3278 (
            .O(N__14601),
            .I(counter_RNI4HQB1Z0Z_5));
    LocalMux I__3277 (
            .O(N__14596),
            .I(counter_RNI4HQB1Z0Z_5));
    LocalMux I__3276 (
            .O(N__14591),
            .I(counter_RNI4HQB1Z0Z_5));
    InMux I__3275 (
            .O(N__14584),
            .I(counter_cry_4));
    CascadeMux I__3274 (
            .O(N__14581),
            .I(N__14578));
    InMux I__3273 (
            .O(N__14578),
            .I(N__14574));
    InMux I__3272 (
            .O(N__14577),
            .I(N__14566));
    LocalMux I__3271 (
            .O(N__14574),
            .I(N__14563));
    InMux I__3270 (
            .O(N__14573),
            .I(N__14556));
    InMux I__3269 (
            .O(N__14572),
            .I(N__14556));
    InMux I__3268 (
            .O(N__14571),
            .I(N__14556));
    InMux I__3267 (
            .O(N__14570),
            .I(N__14551));
    InMux I__3266 (
            .O(N__14569),
            .I(N__14551));
    LocalMux I__3265 (
            .O(N__14566),
            .I(counterZ0Z_5));
    Odrv4 I__3264 (
            .O(N__14563),
            .I(counterZ0Z_5));
    LocalMux I__3263 (
            .O(N__14556),
            .I(counterZ0Z_5));
    LocalMux I__3262 (
            .O(N__14551),
            .I(counterZ0Z_5));
    InMux I__3261 (
            .O(N__14542),
            .I(N__14527));
    InMux I__3260 (
            .O(N__14541),
            .I(N__14522));
    InMux I__3259 (
            .O(N__14540),
            .I(N__14522));
    InMux I__3258 (
            .O(N__14539),
            .I(N__14518));
    InMux I__3257 (
            .O(N__14538),
            .I(N__14515));
    InMux I__3256 (
            .O(N__14537),
            .I(N__14508));
    InMux I__3255 (
            .O(N__14536),
            .I(N__14508));
    InMux I__3254 (
            .O(N__14535),
            .I(N__14508));
    InMux I__3253 (
            .O(N__14534),
            .I(N__14505));
    InMux I__3252 (
            .O(N__14533),
            .I(N__14500));
    InMux I__3251 (
            .O(N__14532),
            .I(N__14500));
    InMux I__3250 (
            .O(N__14531),
            .I(N__14495));
    InMux I__3249 (
            .O(N__14530),
            .I(N__14495));
    LocalMux I__3248 (
            .O(N__14527),
            .I(N__14490));
    LocalMux I__3247 (
            .O(N__14522),
            .I(N__14490));
    InMux I__3246 (
            .O(N__14521),
            .I(N__14487));
    LocalMux I__3245 (
            .O(N__14518),
            .I(N__14482));
    LocalMux I__3244 (
            .O(N__14515),
            .I(N__14482));
    LocalMux I__3243 (
            .O(N__14508),
            .I(N__14479));
    LocalMux I__3242 (
            .O(N__14505),
            .I(N__14474));
    LocalMux I__3241 (
            .O(N__14500),
            .I(N__14474));
    LocalMux I__3240 (
            .O(N__14495),
            .I(N__14471));
    Span4Mux_h I__3239 (
            .O(N__14490),
            .I(N__14466));
    LocalMux I__3238 (
            .O(N__14487),
            .I(N__14466));
    Span12Mux_s9_h I__3237 (
            .O(N__14482),
            .I(N__14463));
    Span4Mux_h I__3236 (
            .O(N__14479),
            .I(N__14460));
    Span4Mux_v I__3235 (
            .O(N__14474),
            .I(N__14455));
    Span4Mux_h I__3234 (
            .O(N__14471),
            .I(N__14455));
    Span4Mux_v I__3233 (
            .O(N__14466),
            .I(N__14452));
    Odrv12 I__3232 (
            .O(N__14463),
            .I(SDATA1_c));
    Odrv4 I__3231 (
            .O(N__14460),
            .I(SDATA1_c));
    Odrv4 I__3230 (
            .O(N__14455),
            .I(SDATA1_c));
    Odrv4 I__3229 (
            .O(N__14452),
            .I(SDATA1_c));
    CascadeMux I__3228 (
            .O(N__14443),
            .I(N__14437));
    InMux I__3227 (
            .O(N__14442),
            .I(N__14430));
    InMux I__3226 (
            .O(N__14441),
            .I(N__14427));
    InMux I__3225 (
            .O(N__14440),
            .I(N__14424));
    InMux I__3224 (
            .O(N__14437),
            .I(N__14421));
    InMux I__3223 (
            .O(N__14436),
            .I(N__14418));
    InMux I__3222 (
            .O(N__14435),
            .I(N__14411));
    InMux I__3221 (
            .O(N__14434),
            .I(N__14411));
    InMux I__3220 (
            .O(N__14433),
            .I(N__14411));
    LocalMux I__3219 (
            .O(N__14430),
            .I(N__14408));
    LocalMux I__3218 (
            .O(N__14427),
            .I(slaveselectZ0));
    LocalMux I__3217 (
            .O(N__14424),
            .I(slaveselectZ0));
    LocalMux I__3216 (
            .O(N__14421),
            .I(slaveselectZ0));
    LocalMux I__3215 (
            .O(N__14418),
            .I(slaveselectZ0));
    LocalMux I__3214 (
            .O(N__14411),
            .I(slaveselectZ0));
    Odrv4 I__3213 (
            .O(N__14408),
            .I(slaveselectZ0));
    CascadeMux I__3212 (
            .O(N__14395),
            .I(N__14391));
    InMux I__3211 (
            .O(N__14394),
            .I(N__14387));
    InMux I__3210 (
            .O(N__14391),
            .I(N__14384));
    InMux I__3209 (
            .O(N__14390),
            .I(N__14381));
    LocalMux I__3208 (
            .O(N__14387),
            .I(un5_slaveselect));
    LocalMux I__3207 (
            .O(N__14384),
            .I(un5_slaveselect));
    LocalMux I__3206 (
            .O(N__14381),
            .I(un5_slaveselect));
    IoInMux I__3205 (
            .O(N__14374),
            .I(N__14371));
    LocalMux I__3204 (
            .O(N__14371),
            .I(N__14367));
    InMux I__3203 (
            .O(N__14370),
            .I(N__14364));
    Odrv4 I__3202 (
            .O(N__14367),
            .I(SDATA2_c));
    LocalMux I__3201 (
            .O(N__14364),
            .I(SDATA2_c));
    InMux I__3200 (
            .O(N__14359),
            .I(N__14355));
    InMux I__3199 (
            .O(N__14358),
            .I(N__14352));
    LocalMux I__3198 (
            .O(N__14355),
            .I(N__14348));
    LocalMux I__3197 (
            .O(N__14352),
            .I(N__14336));
    ClkMux I__3196 (
            .O(N__14351),
            .I(N__14311));
    Glb2LocalMux I__3195 (
            .O(N__14348),
            .I(N__14311));
    ClkMux I__3194 (
            .O(N__14347),
            .I(N__14311));
    ClkMux I__3193 (
            .O(N__14346),
            .I(N__14311));
    ClkMux I__3192 (
            .O(N__14345),
            .I(N__14311));
    ClkMux I__3191 (
            .O(N__14344),
            .I(N__14311));
    ClkMux I__3190 (
            .O(N__14343),
            .I(N__14311));
    ClkMux I__3189 (
            .O(N__14342),
            .I(N__14311));
    ClkMux I__3188 (
            .O(N__14341),
            .I(N__14311));
    ClkMux I__3187 (
            .O(N__14340),
            .I(N__14311));
    ClkMux I__3186 (
            .O(N__14339),
            .I(N__14311));
    Glb2LocalMux I__3185 (
            .O(N__14336),
            .I(N__14311));
    GlobalMux I__3184 (
            .O(N__14311),
            .I(N__14308));
    gio2CtrlBuf I__3183 (
            .O(N__14308),
            .I(Clock12MHz_c_g));
    CascadeMux I__3182 (
            .O(N__14305),
            .I(chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_));
    InMux I__3181 (
            .O(N__14302),
            .I(N__14299));
    LocalMux I__3180 (
            .O(N__14299),
            .I(N__14296));
    Span4Mux_v I__3179 (
            .O(N__14296),
            .I(N__14293));
    Odrv4 I__3178 (
            .O(N__14293),
            .I(beamY_RNII78UPZ0Z_4));
    CascadeMux I__3177 (
            .O(N__14290),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_));
    CascadeMux I__3176 (
            .O(N__14287),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_));
    InMux I__3175 (
            .O(N__14284),
            .I(N__14269));
    InMux I__3174 (
            .O(N__14283),
            .I(N__14269));
    InMux I__3173 (
            .O(N__14282),
            .I(N__14260));
    InMux I__3172 (
            .O(N__14281),
            .I(N__14260));
    InMux I__3171 (
            .O(N__14280),
            .I(N__14257));
    InMux I__3170 (
            .O(N__14279),
            .I(N__14252));
    InMux I__3169 (
            .O(N__14278),
            .I(N__14252));
    InMux I__3168 (
            .O(N__14277),
            .I(N__14245));
    InMux I__3167 (
            .O(N__14276),
            .I(N__14245));
    InMux I__3166 (
            .O(N__14275),
            .I(N__14245));
    InMux I__3165 (
            .O(N__14274),
            .I(N__14242));
    LocalMux I__3164 (
            .O(N__14269),
            .I(N__14239));
    InMux I__3163 (
            .O(N__14268),
            .I(N__14230));
    InMux I__3162 (
            .O(N__14267),
            .I(N__14230));
    InMux I__3161 (
            .O(N__14266),
            .I(N__14230));
    InMux I__3160 (
            .O(N__14265),
            .I(N__14230));
    LocalMux I__3159 (
            .O(N__14260),
            .I(N__14225));
    LocalMux I__3158 (
            .O(N__14257),
            .I(N__14225));
    LocalMux I__3157 (
            .O(N__14252),
            .I(N__14220));
    LocalMux I__3156 (
            .O(N__14245),
            .I(N__14220));
    LocalMux I__3155 (
            .O(N__14242),
            .I(N__14213));
    Span4Mux_v I__3154 (
            .O(N__14239),
            .I(N__14213));
    LocalMux I__3153 (
            .O(N__14230),
            .I(N__14213));
    Span4Mux_h I__3152 (
            .O(N__14225),
            .I(N__14210));
    Odrv12 I__3151 (
            .O(N__14220),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    Odrv4 I__3150 (
            .O(N__14213),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    Odrv4 I__3149 (
            .O(N__14210),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    InMux I__3148 (
            .O(N__14203),
            .I(N__14197));
    InMux I__3147 (
            .O(N__14202),
            .I(N__14197));
    LocalMux I__3146 (
            .O(N__14197),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0));
    CascadeMux I__3145 (
            .O(N__14194),
            .I(chary_if_generate_plus_mult1_un61_sum_c5_cascade_));
    InMux I__3144 (
            .O(N__14191),
            .I(N__14188));
    LocalMux I__3143 (
            .O(N__14188),
            .I(N__14185));
    Span4Mux_s3_v I__3142 (
            .O(N__14185),
            .I(N__14181));
    InMux I__3141 (
            .O(N__14184),
            .I(N__14178));
    Odrv4 I__3140 (
            .O(N__14181),
            .I(un1_counter_0_1));
    LocalMux I__3139 (
            .O(N__14178),
            .I(un1_counter_0_1));
    InMux I__3138 (
            .O(N__14173),
            .I(N__14167));
    InMux I__3137 (
            .O(N__14172),
            .I(N__14164));
    InMux I__3136 (
            .O(N__14171),
            .I(N__14161));
    InMux I__3135 (
            .O(N__14170),
            .I(N__14158));
    LocalMux I__3134 (
            .O(N__14167),
            .I(un7_slaveselectlt5));
    LocalMux I__3133 (
            .O(N__14164),
            .I(un7_slaveselectlt5));
    LocalMux I__3132 (
            .O(N__14161),
            .I(un7_slaveselectlt5));
    LocalMux I__3131 (
            .O(N__14158),
            .I(un7_slaveselectlt5));
    CascadeMux I__3130 (
            .O(N__14149),
            .I(un1_counter_0_1_cascade_));
    CascadeMux I__3129 (
            .O(N__14146),
            .I(slaveselect_1lto5_0_cascade_));
    InMux I__3128 (
            .O(N__14143),
            .I(N__14137));
    InMux I__3127 (
            .O(N__14142),
            .I(N__14137));
    LocalMux I__3126 (
            .O(N__14137),
            .I(slaveselect_1lto5_1));
    IoInMux I__3125 (
            .O(N__14134),
            .I(N__14130));
    IoInMux I__3124 (
            .O(N__14133),
            .I(N__14127));
    LocalMux I__3123 (
            .O(N__14130),
            .I(N__14122));
    LocalMux I__3122 (
            .O(N__14127),
            .I(N__14122));
    Span4Mux_s3_v I__3121 (
            .O(N__14122),
            .I(N__14119));
    Odrv4 I__3120 (
            .O(N__14119),
            .I(SCLK1_0_i));
    InMux I__3119 (
            .O(N__14116),
            .I(N__14102));
    InMux I__3118 (
            .O(N__14115),
            .I(N__14099));
    InMux I__3117 (
            .O(N__14114),
            .I(N__14094));
    InMux I__3116 (
            .O(N__14113),
            .I(N__14094));
    InMux I__3115 (
            .O(N__14112),
            .I(N__14089));
    InMux I__3114 (
            .O(N__14111),
            .I(N__14089));
    InMux I__3113 (
            .O(N__14110),
            .I(N__14084));
    InMux I__3112 (
            .O(N__14109),
            .I(N__14084));
    InMux I__3111 (
            .O(N__14108),
            .I(N__14081));
    InMux I__3110 (
            .O(N__14107),
            .I(N__14074));
    InMux I__3109 (
            .O(N__14106),
            .I(N__14074));
    InMux I__3108 (
            .O(N__14105),
            .I(N__14074));
    LocalMux I__3107 (
            .O(N__14102),
            .I(counterZ0Z_1));
    LocalMux I__3106 (
            .O(N__14099),
            .I(counterZ0Z_1));
    LocalMux I__3105 (
            .O(N__14094),
            .I(counterZ0Z_1));
    LocalMux I__3104 (
            .O(N__14089),
            .I(counterZ0Z_1));
    LocalMux I__3103 (
            .O(N__14084),
            .I(counterZ0Z_1));
    LocalMux I__3102 (
            .O(N__14081),
            .I(counterZ0Z_1));
    LocalMux I__3101 (
            .O(N__14074),
            .I(counterZ0Z_1));
    CascadeMux I__3100 (
            .O(N__14059),
            .I(N__14050));
    CascadeMux I__3099 (
            .O(N__14058),
            .I(N__14039));
    CascadeMux I__3098 (
            .O(N__14057),
            .I(N__14036));
    InMux I__3097 (
            .O(N__14056),
            .I(N__14032));
    InMux I__3096 (
            .O(N__14055),
            .I(N__14025));
    InMux I__3095 (
            .O(N__14054),
            .I(N__14025));
    InMux I__3094 (
            .O(N__14053),
            .I(N__14025));
    InMux I__3093 (
            .O(N__14050),
            .I(N__14022));
    InMux I__3092 (
            .O(N__14049),
            .I(N__14017));
    InMux I__3091 (
            .O(N__14048),
            .I(N__14017));
    InMux I__3090 (
            .O(N__14047),
            .I(N__14010));
    InMux I__3089 (
            .O(N__14046),
            .I(N__14010));
    InMux I__3088 (
            .O(N__14045),
            .I(N__14010));
    InMux I__3087 (
            .O(N__14044),
            .I(N__14003));
    InMux I__3086 (
            .O(N__14043),
            .I(N__14003));
    InMux I__3085 (
            .O(N__14042),
            .I(N__14003));
    InMux I__3084 (
            .O(N__14039),
            .I(N__14000));
    InMux I__3083 (
            .O(N__14036),
            .I(N__13995));
    InMux I__3082 (
            .O(N__14035),
            .I(N__13995));
    LocalMux I__3081 (
            .O(N__14032),
            .I(counterZ0Z_0));
    LocalMux I__3080 (
            .O(N__14025),
            .I(counterZ0Z_0));
    LocalMux I__3079 (
            .O(N__14022),
            .I(counterZ0Z_0));
    LocalMux I__3078 (
            .O(N__14017),
            .I(counterZ0Z_0));
    LocalMux I__3077 (
            .O(N__14010),
            .I(counterZ0Z_0));
    LocalMux I__3076 (
            .O(N__14003),
            .I(counterZ0Z_0));
    LocalMux I__3075 (
            .O(N__14000),
            .I(counterZ0Z_0));
    LocalMux I__3074 (
            .O(N__13995),
            .I(counterZ0Z_0));
    InMux I__3073 (
            .O(N__13978),
            .I(N__13975));
    LocalMux I__3072 (
            .O(N__13975),
            .I(N__13970));
    InMux I__3071 (
            .O(N__13974),
            .I(N__13965));
    InMux I__3070 (
            .O(N__13973),
            .I(N__13965));
    Odrv4 I__3069 (
            .O(N__13970),
            .I(un7_slaveselectlt2_0));
    LocalMux I__3068 (
            .O(N__13965),
            .I(un7_slaveselectlt2_0));
    CascadeMux I__3067 (
            .O(N__13960),
            .I(N__13957));
    InMux I__3066 (
            .O(N__13957),
            .I(N__13951));
    InMux I__3065 (
            .O(N__13956),
            .I(N__13945));
    InMux I__3064 (
            .O(N__13955),
            .I(N__13940));
    InMux I__3063 (
            .O(N__13954),
            .I(N__13940));
    LocalMux I__3062 (
            .O(N__13951),
            .I(N__13937));
    InMux I__3061 (
            .O(N__13950),
            .I(N__13930));
    InMux I__3060 (
            .O(N__13949),
            .I(N__13930));
    InMux I__3059 (
            .O(N__13948),
            .I(N__13930));
    LocalMux I__3058 (
            .O(N__13945),
            .I(counterZ0Z_2));
    LocalMux I__3057 (
            .O(N__13940),
            .I(counterZ0Z_2));
    Odrv4 I__3056 (
            .O(N__13937),
            .I(counterZ0Z_2));
    LocalMux I__3055 (
            .O(N__13930),
            .I(counterZ0Z_2));
    InMux I__3054 (
            .O(N__13921),
            .I(counter_cry_1));
    CascadeMux I__3053 (
            .O(N__13918),
            .I(N__13912));
    CascadeMux I__3052 (
            .O(N__13917),
            .I(N__13909));
    CascadeMux I__3051 (
            .O(N__13916),
            .I(N__13905));
    InMux I__3050 (
            .O(N__13915),
            .I(N__13900));
    InMux I__3049 (
            .O(N__13912),
            .I(N__13897));
    InMux I__3048 (
            .O(N__13909),
            .I(N__13894));
    InMux I__3047 (
            .O(N__13908),
            .I(N__13889));
    InMux I__3046 (
            .O(N__13905),
            .I(N__13889));
    InMux I__3045 (
            .O(N__13904),
            .I(N__13885));
    InMux I__3044 (
            .O(N__13903),
            .I(N__13882));
    LocalMux I__3043 (
            .O(N__13900),
            .I(N__13877));
    LocalMux I__3042 (
            .O(N__13897),
            .I(N__13877));
    LocalMux I__3041 (
            .O(N__13894),
            .I(N__13874));
    LocalMux I__3040 (
            .O(N__13889),
            .I(N__13871));
    InMux I__3039 (
            .O(N__13888),
            .I(N__13868));
    LocalMux I__3038 (
            .O(N__13885),
            .I(counterZ0Z_3));
    LocalMux I__3037 (
            .O(N__13882),
            .I(counterZ0Z_3));
    Odrv4 I__3036 (
            .O(N__13877),
            .I(counterZ0Z_3));
    Odrv4 I__3035 (
            .O(N__13874),
            .I(counterZ0Z_3));
    Odrv4 I__3034 (
            .O(N__13871),
            .I(counterZ0Z_3));
    LocalMux I__3033 (
            .O(N__13868),
            .I(counterZ0Z_3));
    InMux I__3032 (
            .O(N__13855),
            .I(counter_cry_2));
    InMux I__3031 (
            .O(N__13852),
            .I(N__13846));
    InMux I__3030 (
            .O(N__13851),
            .I(N__13843));
    InMux I__3029 (
            .O(N__13850),
            .I(N__13838));
    InMux I__3028 (
            .O(N__13849),
            .I(N__13838));
    LocalMux I__3027 (
            .O(N__13846),
            .I(counterZ0Z_4));
    LocalMux I__3026 (
            .O(N__13843),
            .I(counterZ0Z_4));
    LocalMux I__3025 (
            .O(N__13838),
            .I(counterZ0Z_4));
    InMux I__3024 (
            .O(N__13831),
            .I(counter_cry_3));
    InMux I__3023 (
            .O(N__13828),
            .I(N__13822));
    InMux I__3022 (
            .O(N__13827),
            .I(N__13822));
    LocalMux I__3021 (
            .O(N__13822),
            .I(content_ram10_0));
    CEMux I__3020 (
            .O(N__13819),
            .I(N__13816));
    LocalMux I__3019 (
            .O(N__13816),
            .I(N__13813));
    Odrv12 I__3018 (
            .O(N__13813),
            .I(content_awe10));
    CascadeMux I__3017 (
            .O(N__13810),
            .I(content_N_35_cascade_));
    InMux I__3016 (
            .O(N__13807),
            .I(N__13804));
    LocalMux I__3015 (
            .O(N__13804),
            .I(content_awe3_1));
    CascadeMux I__3014 (
            .O(N__13801),
            .I(content_awe3_1_cascade_));
    InMux I__3013 (
            .O(N__13798),
            .I(N__13793));
    InMux I__3012 (
            .O(N__13797),
            .I(N__13788));
    InMux I__3011 (
            .O(N__13796),
            .I(N__13788));
    LocalMux I__3010 (
            .O(N__13793),
            .I(content_ram2_0));
    LocalMux I__3009 (
            .O(N__13788),
            .I(content_ram2_0));
    InMux I__3008 (
            .O(N__13783),
            .I(N__13778));
    InMux I__3007 (
            .O(N__13782),
            .I(N__13775));
    InMux I__3006 (
            .O(N__13781),
            .I(N__13772));
    LocalMux I__3005 (
            .O(N__13778),
            .I(content_N_40));
    LocalMux I__3004 (
            .O(N__13775),
            .I(content_N_40));
    LocalMux I__3003 (
            .O(N__13772),
            .I(content_N_40));
    CascadeMux I__3002 (
            .O(N__13765),
            .I(N__13759));
    CascadeMux I__3001 (
            .O(N__13764),
            .I(N__13754));
    CascadeMux I__3000 (
            .O(N__13763),
            .I(N__13751));
    InMux I__2999 (
            .O(N__13762),
            .I(N__13748));
    InMux I__2998 (
            .O(N__13759),
            .I(N__13745));
    InMux I__2997 (
            .O(N__13758),
            .I(N__13736));
    InMux I__2996 (
            .O(N__13757),
            .I(N__13736));
    InMux I__2995 (
            .O(N__13754),
            .I(N__13736));
    InMux I__2994 (
            .O(N__13751),
            .I(N__13736));
    LocalMux I__2993 (
            .O(N__13748),
            .I(content_N_35));
    LocalMux I__2992 (
            .O(N__13745),
            .I(content_N_35));
    LocalMux I__2991 (
            .O(N__13736),
            .I(content_N_35));
    CascadeMux I__2990 (
            .O(N__13729),
            .I(content_awe1_0_a2_0_cascade_));
    CascadeMux I__2989 (
            .O(N__13726),
            .I(N__13722));
    InMux I__2988 (
            .O(N__13725),
            .I(N__13717));
    InMux I__2987 (
            .O(N__13722),
            .I(N__13717));
    LocalMux I__2986 (
            .O(N__13717),
            .I(N__13713));
    InMux I__2985 (
            .O(N__13716),
            .I(N__13710));
    Span4Mux_h I__2984 (
            .O(N__13713),
            .I(N__13707));
    LocalMux I__2983 (
            .O(N__13710),
            .I(content_ram1_0));
    Odrv4 I__2982 (
            .O(N__13707),
            .I(content_ram1_0));
    CascadeMux I__2981 (
            .O(N__13702),
            .I(un7_slaveselectlt5_cascade_));
    InMux I__2980 (
            .O(N__13699),
            .I(N__13692));
    InMux I__2979 (
            .O(N__13698),
            .I(N__13687));
    InMux I__2978 (
            .O(N__13697),
            .I(N__13687));
    InMux I__2977 (
            .O(N__13696),
            .I(N__13682));
    InMux I__2976 (
            .O(N__13695),
            .I(N__13682));
    LocalMux I__2975 (
            .O(N__13692),
            .I(N_190_i));
    LocalMux I__2974 (
            .O(N__13687),
            .I(N_190_i));
    LocalMux I__2973 (
            .O(N__13682),
            .I(N_190_i));
    CascadeMux I__2972 (
            .O(N__13675),
            .I(N__13672));
    InMux I__2971 (
            .O(N__13672),
            .I(N__13669));
    LocalMux I__2970 (
            .O(N__13669),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0));
    InMux I__2969 (
            .O(N__13666),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__2968 (
            .O(N__13663),
            .I(N__13660));
    InMux I__2967 (
            .O(N__13660),
            .I(N__13657));
    LocalMux I__2966 (
            .O(N__13657),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0));
    CascadeMux I__2965 (
            .O(N__13654),
            .I(N__13651));
    InMux I__2964 (
            .O(N__13651),
            .I(N__13648));
    LocalMux I__2963 (
            .O(N__13648),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1));
    InMux I__2962 (
            .O(N__13645),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2961 (
            .O(N__13642),
            .I(N__13639));
    LocalMux I__2960 (
            .O(N__13639),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41));
    CascadeMux I__2959 (
            .O(N__13636),
            .I(N__13632));
    InMux I__2958 (
            .O(N__13635),
            .I(N__13627));
    InMux I__2957 (
            .O(N__13632),
            .I(N__13627));
    LocalMux I__2956 (
            .O(N__13627),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02));
    InMux I__2955 (
            .O(N__13624),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__2954 (
            .O(N__13621),
            .I(N__13618));
    InMux I__2953 (
            .O(N__13618),
            .I(N__13615));
    LocalMux I__2952 (
            .O(N__13615),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81));
    InMux I__2951 (
            .O(N__13612),
            .I(N__13609));
    LocalMux I__2950 (
            .O(N__13609),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__2949 (
            .O(N__13606),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__2948 (
            .O(N__13603),
            .I(N__13600));
    LocalMux I__2947 (
            .O(N__13600),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__2946 (
            .O(N__13597),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__2945 (
            .O(N__13594),
            .I(N__13587));
    InMux I__2944 (
            .O(N__13593),
            .I(N__13584));
    InMux I__2943 (
            .O(N__13592),
            .I(N__13577));
    InMux I__2942 (
            .O(N__13591),
            .I(N__13577));
    InMux I__2941 (
            .O(N__13590),
            .I(N__13577));
    LocalMux I__2940 (
            .O(N__13587),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42));
    LocalMux I__2939 (
            .O(N__13584),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42));
    LocalMux I__2938 (
            .O(N__13577),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42));
    CascadeMux I__2937 (
            .O(N__13570),
            .I(N__13565));
    CascadeMux I__2936 (
            .O(N__13569),
            .I(N__13561));
    InMux I__2935 (
            .O(N__13568),
            .I(N__13557));
    InMux I__2934 (
            .O(N__13565),
            .I(N__13548));
    InMux I__2933 (
            .O(N__13564),
            .I(N__13548));
    InMux I__2932 (
            .O(N__13561),
            .I(N__13548));
    InMux I__2931 (
            .O(N__13560),
            .I(N__13548));
    LocalMux I__2930 (
            .O(N__13557),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0));
    LocalMux I__2929 (
            .O(N__13548),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0));
    InMux I__2928 (
            .O(N__13543),
            .I(N__13540));
    LocalMux I__2927 (
            .O(N__13540),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7));
    InMux I__2926 (
            .O(N__13537),
            .I(N__13534));
    LocalMux I__2925 (
            .O(N__13534),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__2924 (
            .O(N__13531),
            .I(N__13526));
    InMux I__2923 (
            .O(N__13530),
            .I(N__13521));
    InMux I__2922 (
            .O(N__13529),
            .I(N__13521));
    LocalMux I__2921 (
            .O(N__13526),
            .I(N__13515));
    LocalMux I__2920 (
            .O(N__13521),
            .I(N__13512));
    InMux I__2919 (
            .O(N__13520),
            .I(N__13509));
    InMux I__2918 (
            .O(N__13519),
            .I(N__13506));
    InMux I__2917 (
            .O(N__13518),
            .I(N__13503));
    Span4Mux_h I__2916 (
            .O(N__13515),
            .I(N__13500));
    Odrv4 I__2915 (
            .O(N__13512),
            .I(beamY_RNI9DLCZ0Z_1));
    LocalMux I__2914 (
            .O(N__13509),
            .I(beamY_RNI9DLCZ0Z_1));
    LocalMux I__2913 (
            .O(N__13506),
            .I(beamY_RNI9DLCZ0Z_1));
    LocalMux I__2912 (
            .O(N__13503),
            .I(beamY_RNI9DLCZ0Z_1));
    Odrv4 I__2911 (
            .O(N__13500),
            .I(beamY_RNI9DLCZ0Z_1));
    InMux I__2910 (
            .O(N__13489),
            .I(bfn_9_8_0_));
    InMux I__2909 (
            .O(N__13486),
            .I(N__13482));
    InMux I__2908 (
            .O(N__13485),
            .I(N__13477));
    LocalMux I__2907 (
            .O(N__13482),
            .I(N__13474));
    InMux I__2906 (
            .O(N__13481),
            .I(N__13469));
    InMux I__2905 (
            .O(N__13480),
            .I(N__13469));
    LocalMux I__2904 (
            .O(N__13477),
            .I(N__13459));
    Span4Mux_v I__2903 (
            .O(N__13474),
            .I(N__13459));
    LocalMux I__2902 (
            .O(N__13469),
            .I(N__13459));
    InMux I__2901 (
            .O(N__13468),
            .I(N__13456));
    InMux I__2900 (
            .O(N__13467),
            .I(N__13453));
    InMux I__2899 (
            .O(N__13466),
            .I(N__13448));
    Span4Mux_h I__2898 (
            .O(N__13459),
            .I(N__13445));
    LocalMux I__2897 (
            .O(N__13456),
            .I(N__13440));
    LocalMux I__2896 (
            .O(N__13453),
            .I(N__13440));
    InMux I__2895 (
            .O(N__13452),
            .I(N__13435));
    InMux I__2894 (
            .O(N__13451),
            .I(N__13435));
    LocalMux I__2893 (
            .O(N__13448),
            .I(beamYZ0Z_9));
    Odrv4 I__2892 (
            .O(N__13445),
            .I(beamYZ0Z_9));
    Odrv4 I__2891 (
            .O(N__13440),
            .I(beamYZ0Z_9));
    LocalMux I__2890 (
            .O(N__13435),
            .I(beamYZ0Z_9));
    ClkMux I__2889 (
            .O(N__13426),
            .I(N__13399));
    ClkMux I__2888 (
            .O(N__13425),
            .I(N__13399));
    ClkMux I__2887 (
            .O(N__13424),
            .I(N__13399));
    ClkMux I__2886 (
            .O(N__13423),
            .I(N__13399));
    ClkMux I__2885 (
            .O(N__13422),
            .I(N__13399));
    ClkMux I__2884 (
            .O(N__13421),
            .I(N__13399));
    ClkMux I__2883 (
            .O(N__13420),
            .I(N__13399));
    ClkMux I__2882 (
            .O(N__13419),
            .I(N__13399));
    ClkMux I__2881 (
            .O(N__13418),
            .I(N__13399));
    GlobalMux I__2880 (
            .O(N__13399),
            .I(N__13396));
    gio2CtrlBuf I__2879 (
            .O(N__13396),
            .I(PixelClock_g));
    CEMux I__2878 (
            .O(N__13393),
            .I(N__13388));
    CEMux I__2877 (
            .O(N__13392),
            .I(N__13385));
    InMux I__2876 (
            .O(N__13391),
            .I(N__13381));
    LocalMux I__2875 (
            .O(N__13388),
            .I(N__13378));
    LocalMux I__2874 (
            .O(N__13385),
            .I(N__13375));
    InMux I__2873 (
            .O(N__13384),
            .I(N__13370));
    LocalMux I__2872 (
            .O(N__13381),
            .I(N__13367));
    Span4Mux_v I__2871 (
            .O(N__13378),
            .I(N__13364));
    Span4Mux_v I__2870 (
            .O(N__13375),
            .I(N__13361));
    InMux I__2869 (
            .O(N__13374),
            .I(N__13355));
    InMux I__2868 (
            .O(N__13373),
            .I(N__13355));
    LocalMux I__2867 (
            .O(N__13370),
            .I(N__13352));
    Span4Mux_v I__2866 (
            .O(N__13367),
            .I(N__13345));
    Span4Mux_h I__2865 (
            .O(N__13364),
            .I(N__13345));
    Span4Mux_h I__2864 (
            .O(N__13361),
            .I(N__13345));
    InMux I__2863 (
            .O(N__13360),
            .I(N__13342));
    LocalMux I__2862 (
            .O(N__13355),
            .I(N__13339));
    Span12Mux_s8_v I__2861 (
            .O(N__13352),
            .I(N__13336));
    Span4Mux_h I__2860 (
            .O(N__13345),
            .I(N__13333));
    LocalMux I__2859 (
            .O(N__13342),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__2858 (
            .O(N__13339),
            .I(beamX_RNI5457Z0Z_5));
    Odrv12 I__2857 (
            .O(N__13336),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__2856 (
            .O(N__13333),
            .I(beamX_RNI5457Z0Z_5));
    InMux I__2855 (
            .O(N__13324),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__2854 (
            .O(N__13321),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__2853 (
            .O(N__13318),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__2852 (
            .O(N__13315),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__2851 (
            .O(N__13312),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__2850 (
            .O(N__13309),
            .I(N__13306));
    LocalMux I__2849 (
            .O(N__13306),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__2848 (
            .O(N__13303),
            .I(N__13300));
    LocalMux I__2847 (
            .O(N__13300),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__2846 (
            .O(N__13297),
            .I(N__13291));
    CascadeMux I__2845 (
            .O(N__13296),
            .I(N__13284));
    CascadeMux I__2844 (
            .O(N__13295),
            .I(N__13280));
    CascadeMux I__2843 (
            .O(N__13294),
            .I(N__13277));
    LocalMux I__2842 (
            .O(N__13291),
            .I(N__13273));
    InMux I__2841 (
            .O(N__13290),
            .I(N__13268));
    InMux I__2840 (
            .O(N__13289),
            .I(N__13268));
    CascadeMux I__2839 (
            .O(N__13288),
            .I(N__13259));
    InMux I__2838 (
            .O(N__13287),
            .I(N__13253));
    InMux I__2837 (
            .O(N__13284),
            .I(N__13248));
    InMux I__2836 (
            .O(N__13283),
            .I(N__13243));
    InMux I__2835 (
            .O(N__13280),
            .I(N__13243));
    InMux I__2834 (
            .O(N__13277),
            .I(N__13240));
    InMux I__2833 (
            .O(N__13276),
            .I(N__13237));
    Span4Mux_v I__2832 (
            .O(N__13273),
            .I(N__13232));
    LocalMux I__2831 (
            .O(N__13268),
            .I(N__13232));
    InMux I__2830 (
            .O(N__13267),
            .I(N__13227));
    InMux I__2829 (
            .O(N__13266),
            .I(N__13227));
    CascadeMux I__2828 (
            .O(N__13265),
            .I(N__13223));
    InMux I__2827 (
            .O(N__13264),
            .I(N__13220));
    InMux I__2826 (
            .O(N__13263),
            .I(N__13213));
    InMux I__2825 (
            .O(N__13262),
            .I(N__13213));
    InMux I__2824 (
            .O(N__13259),
            .I(N__13213));
    InMux I__2823 (
            .O(N__13258),
            .I(N__13210));
    InMux I__2822 (
            .O(N__13257),
            .I(N__13205));
    InMux I__2821 (
            .O(N__13256),
            .I(N__13205));
    LocalMux I__2820 (
            .O(N__13253),
            .I(N__13202));
    InMux I__2819 (
            .O(N__13252),
            .I(N__13198));
    InMux I__2818 (
            .O(N__13251),
            .I(N__13194));
    LocalMux I__2817 (
            .O(N__13248),
            .I(N__13187));
    LocalMux I__2816 (
            .O(N__13243),
            .I(N__13187));
    LocalMux I__2815 (
            .O(N__13240),
            .I(N__13187));
    LocalMux I__2814 (
            .O(N__13237),
            .I(N__13180));
    Span4Mux_s2_v I__2813 (
            .O(N__13232),
            .I(N__13180));
    LocalMux I__2812 (
            .O(N__13227),
            .I(N__13180));
    InMux I__2811 (
            .O(N__13226),
            .I(N__13175));
    InMux I__2810 (
            .O(N__13223),
            .I(N__13175));
    LocalMux I__2809 (
            .O(N__13220),
            .I(N__13166));
    LocalMux I__2808 (
            .O(N__13213),
            .I(N__13166));
    LocalMux I__2807 (
            .O(N__13210),
            .I(N__13166));
    LocalMux I__2806 (
            .O(N__13205),
            .I(N__13166));
    Span4Mux_v I__2805 (
            .O(N__13202),
            .I(N__13163));
    InMux I__2804 (
            .O(N__13201),
            .I(N__13160));
    LocalMux I__2803 (
            .O(N__13198),
            .I(N__13157));
    InMux I__2802 (
            .O(N__13197),
            .I(N__13152));
    LocalMux I__2801 (
            .O(N__13194),
            .I(N__13147));
    Span12Mux_s6_h I__2800 (
            .O(N__13187),
            .I(N__13147));
    Span4Mux_v I__2799 (
            .O(N__13180),
            .I(N__13140));
    LocalMux I__2798 (
            .O(N__13175),
            .I(N__13140));
    Span4Mux_v I__2797 (
            .O(N__13166),
            .I(N__13140));
    Span4Mux_h I__2796 (
            .O(N__13163),
            .I(N__13135));
    LocalMux I__2795 (
            .O(N__13160),
            .I(N__13135));
    Span4Mux_h I__2794 (
            .O(N__13157),
            .I(N__13132));
    InMux I__2793 (
            .O(N__13156),
            .I(N__13127));
    InMux I__2792 (
            .O(N__13155),
            .I(N__13127));
    LocalMux I__2791 (
            .O(N__13152),
            .I(beamYZ0Z_1));
    Odrv12 I__2790 (
            .O(N__13147),
            .I(beamYZ0Z_1));
    Odrv4 I__2789 (
            .O(N__13140),
            .I(beamYZ0Z_1));
    Odrv4 I__2788 (
            .O(N__13135),
            .I(beamYZ0Z_1));
    Odrv4 I__2787 (
            .O(N__13132),
            .I(beamYZ0Z_1));
    LocalMux I__2786 (
            .O(N__13127),
            .I(beamYZ0Z_1));
    CascadeMux I__2785 (
            .O(N__13114),
            .I(N__13110));
    InMux I__2784 (
            .O(N__13113),
            .I(N__13102));
    InMux I__2783 (
            .O(N__13110),
            .I(N__13094));
    InMux I__2782 (
            .O(N__13109),
            .I(N__13094));
    InMux I__2781 (
            .O(N__13108),
            .I(N__13086));
    InMux I__2780 (
            .O(N__13107),
            .I(N__13083));
    InMux I__2779 (
            .O(N__13106),
            .I(N__13080));
    CascadeMux I__2778 (
            .O(N__13105),
            .I(N__13077));
    LocalMux I__2777 (
            .O(N__13102),
            .I(N__13071));
    InMux I__2776 (
            .O(N__13101),
            .I(N__13068));
    InMux I__2775 (
            .O(N__13100),
            .I(N__13063));
    InMux I__2774 (
            .O(N__13099),
            .I(N__13063));
    LocalMux I__2773 (
            .O(N__13094),
            .I(N__13060));
    InMux I__2772 (
            .O(N__13093),
            .I(N__13057));
    InMux I__2771 (
            .O(N__13092),
            .I(N__13052));
    InMux I__2770 (
            .O(N__13091),
            .I(N__13045));
    InMux I__2769 (
            .O(N__13090),
            .I(N__13045));
    InMux I__2768 (
            .O(N__13089),
            .I(N__13045));
    LocalMux I__2767 (
            .O(N__13086),
            .I(N__13038));
    LocalMux I__2766 (
            .O(N__13083),
            .I(N__13038));
    LocalMux I__2765 (
            .O(N__13080),
            .I(N__13038));
    InMux I__2764 (
            .O(N__13077),
            .I(N__13033));
    InMux I__2763 (
            .O(N__13076),
            .I(N__13033));
    InMux I__2762 (
            .O(N__13075),
            .I(N__13030));
    CascadeMux I__2761 (
            .O(N__13074),
            .I(N__13027));
    Span4Mux_h I__2760 (
            .O(N__13071),
            .I(N__13023));
    LocalMux I__2759 (
            .O(N__13068),
            .I(N__13020));
    LocalMux I__2758 (
            .O(N__13063),
            .I(N__13017));
    Span4Mux_h I__2757 (
            .O(N__13060),
            .I(N__13014));
    LocalMux I__2756 (
            .O(N__13057),
            .I(N__13011));
    InMux I__2755 (
            .O(N__13056),
            .I(N__13006));
    InMux I__2754 (
            .O(N__13055),
            .I(N__13006));
    LocalMux I__2753 (
            .O(N__13052),
            .I(N__13003));
    LocalMux I__2752 (
            .O(N__13045),
            .I(N__12998));
    Span4Mux_s3_v I__2751 (
            .O(N__13038),
            .I(N__12998));
    LocalMux I__2750 (
            .O(N__13033),
            .I(N__12993));
    LocalMux I__2749 (
            .O(N__13030),
            .I(N__12993));
    InMux I__2748 (
            .O(N__13027),
            .I(N__12990));
    InMux I__2747 (
            .O(N__13026),
            .I(N__12987));
    Span4Mux_v I__2746 (
            .O(N__13023),
            .I(N__12982));
    Span4Mux_h I__2745 (
            .O(N__13020),
            .I(N__12982));
    Span4Mux_v I__2744 (
            .O(N__13017),
            .I(N__12975));
    Span4Mux_v I__2743 (
            .O(N__13014),
            .I(N__12975));
    Span4Mux_h I__2742 (
            .O(N__13011),
            .I(N__12975));
    LocalMux I__2741 (
            .O(N__13006),
            .I(N__12968));
    Span4Mux_s3_v I__2740 (
            .O(N__13003),
            .I(N__12968));
    Span4Mux_h I__2739 (
            .O(N__12998),
            .I(N__12968));
    Span4Mux_v I__2738 (
            .O(N__12993),
            .I(N__12965));
    LocalMux I__2737 (
            .O(N__12990),
            .I(beamYZ0Z_0));
    LocalMux I__2736 (
            .O(N__12987),
            .I(beamYZ0Z_0));
    Odrv4 I__2735 (
            .O(N__12982),
            .I(beamYZ0Z_0));
    Odrv4 I__2734 (
            .O(N__12975),
            .I(beamYZ0Z_0));
    Odrv4 I__2733 (
            .O(N__12968),
            .I(beamYZ0Z_0));
    Odrv4 I__2732 (
            .O(N__12965),
            .I(beamYZ0Z_0));
    CascadeMux I__2731 (
            .O(N__12952),
            .I(N__12949));
    InMux I__2730 (
            .O(N__12949),
            .I(N__12946));
    LocalMux I__2729 (
            .O(N__12946),
            .I(N__12943));
    Span4Mux_h I__2728 (
            .O(N__12943),
            .I(N__12940));
    Span4Mux_h I__2727 (
            .O(N__12940),
            .I(N__12937));
    Odrv4 I__2726 (
            .O(N__12937),
            .I(g2_1_1_0));
    CascadeMux I__2725 (
            .O(N__12934),
            .I(N__12927));
    CascadeMux I__2724 (
            .O(N__12933),
            .I(N__12923));
    CascadeMux I__2723 (
            .O(N__12932),
            .I(N__12914));
    CascadeMux I__2722 (
            .O(N__12931),
            .I(N__12907));
    InMux I__2721 (
            .O(N__12930),
            .I(N__12904));
    InMux I__2720 (
            .O(N__12927),
            .I(N__12901));
    InMux I__2719 (
            .O(N__12926),
            .I(N__12892));
    InMux I__2718 (
            .O(N__12923),
            .I(N__12892));
    InMux I__2717 (
            .O(N__12922),
            .I(N__12892));
    InMux I__2716 (
            .O(N__12921),
            .I(N__12892));
    InMux I__2715 (
            .O(N__12920),
            .I(N__12889));
    CascadeMux I__2714 (
            .O(N__12919),
            .I(N__12883));
    InMux I__2713 (
            .O(N__12918),
            .I(N__12872));
    InMux I__2712 (
            .O(N__12917),
            .I(N__12867));
    InMux I__2711 (
            .O(N__12914),
            .I(N__12867));
    InMux I__2710 (
            .O(N__12913),
            .I(N__12862));
    InMux I__2709 (
            .O(N__12912),
            .I(N__12862));
    InMux I__2708 (
            .O(N__12911),
            .I(N__12853));
    InMux I__2707 (
            .O(N__12910),
            .I(N__12848));
    InMux I__2706 (
            .O(N__12907),
            .I(N__12848));
    LocalMux I__2705 (
            .O(N__12904),
            .I(N__12839));
    LocalMux I__2704 (
            .O(N__12901),
            .I(N__12839));
    LocalMux I__2703 (
            .O(N__12892),
            .I(N__12839));
    LocalMux I__2702 (
            .O(N__12889),
            .I(N__12839));
    InMux I__2701 (
            .O(N__12888),
            .I(N__12835));
    InMux I__2700 (
            .O(N__12887),
            .I(N__12830));
    InMux I__2699 (
            .O(N__12886),
            .I(N__12830));
    InMux I__2698 (
            .O(N__12883),
            .I(N__12825));
    InMux I__2697 (
            .O(N__12882),
            .I(N__12825));
    InMux I__2696 (
            .O(N__12881),
            .I(N__12822));
    InMux I__2695 (
            .O(N__12880),
            .I(N__12815));
    InMux I__2694 (
            .O(N__12879),
            .I(N__12815));
    InMux I__2693 (
            .O(N__12878),
            .I(N__12815));
    InMux I__2692 (
            .O(N__12877),
            .I(N__12808));
    InMux I__2691 (
            .O(N__12876),
            .I(N__12808));
    InMux I__2690 (
            .O(N__12875),
            .I(N__12808));
    LocalMux I__2689 (
            .O(N__12872),
            .I(N__12799));
    LocalMux I__2688 (
            .O(N__12867),
            .I(N__12799));
    LocalMux I__2687 (
            .O(N__12862),
            .I(N__12796));
    InMux I__2686 (
            .O(N__12861),
            .I(N__12789));
    InMux I__2685 (
            .O(N__12860),
            .I(N__12789));
    InMux I__2684 (
            .O(N__12859),
            .I(N__12789));
    InMux I__2683 (
            .O(N__12858),
            .I(N__12786));
    InMux I__2682 (
            .O(N__12857),
            .I(N__12783));
    InMux I__2681 (
            .O(N__12856),
            .I(N__12780));
    LocalMux I__2680 (
            .O(N__12853),
            .I(N__12775));
    LocalMux I__2679 (
            .O(N__12848),
            .I(N__12775));
    Span4Mux_v I__2678 (
            .O(N__12839),
            .I(N__12772));
    InMux I__2677 (
            .O(N__12838),
            .I(N__12769));
    LocalMux I__2676 (
            .O(N__12835),
            .I(N__12756));
    LocalMux I__2675 (
            .O(N__12830),
            .I(N__12756));
    LocalMux I__2674 (
            .O(N__12825),
            .I(N__12756));
    LocalMux I__2673 (
            .O(N__12822),
            .I(N__12756));
    LocalMux I__2672 (
            .O(N__12815),
            .I(N__12756));
    LocalMux I__2671 (
            .O(N__12808),
            .I(N__12756));
    InMux I__2670 (
            .O(N__12807),
            .I(N__12751));
    InMux I__2669 (
            .O(N__12806),
            .I(N__12751));
    CascadeMux I__2668 (
            .O(N__12805),
            .I(N__12747));
    InMux I__2667 (
            .O(N__12804),
            .I(N__12739));
    Span4Mux_h I__2666 (
            .O(N__12799),
            .I(N__12736));
    Span4Mux_h I__2665 (
            .O(N__12796),
            .I(N__12725));
    LocalMux I__2664 (
            .O(N__12789),
            .I(N__12725));
    LocalMux I__2663 (
            .O(N__12786),
            .I(N__12725));
    LocalMux I__2662 (
            .O(N__12783),
            .I(N__12725));
    LocalMux I__2661 (
            .O(N__12780),
            .I(N__12725));
    Span12Mux_s6_v I__2660 (
            .O(N__12775),
            .I(N__12718));
    Sp12to4 I__2659 (
            .O(N__12772),
            .I(N__12718));
    LocalMux I__2658 (
            .O(N__12769),
            .I(N__12718));
    Span4Mux_v I__2657 (
            .O(N__12756),
            .I(N__12713));
    LocalMux I__2656 (
            .O(N__12751),
            .I(N__12713));
    InMux I__2655 (
            .O(N__12750),
            .I(N__12710));
    InMux I__2654 (
            .O(N__12747),
            .I(N__12707));
    InMux I__2653 (
            .O(N__12746),
            .I(N__12700));
    InMux I__2652 (
            .O(N__12745),
            .I(N__12700));
    InMux I__2651 (
            .O(N__12744),
            .I(N__12700));
    InMux I__2650 (
            .O(N__12743),
            .I(N__12695));
    InMux I__2649 (
            .O(N__12742),
            .I(N__12695));
    LocalMux I__2648 (
            .O(N__12739),
            .I(beamYZ0Z_2));
    Odrv4 I__2647 (
            .O(N__12736),
            .I(beamYZ0Z_2));
    Odrv4 I__2646 (
            .O(N__12725),
            .I(beamYZ0Z_2));
    Odrv12 I__2645 (
            .O(N__12718),
            .I(beamYZ0Z_2));
    Odrv4 I__2644 (
            .O(N__12713),
            .I(beamYZ0Z_2));
    LocalMux I__2643 (
            .O(N__12710),
            .I(beamYZ0Z_2));
    LocalMux I__2642 (
            .O(N__12707),
            .I(beamYZ0Z_2));
    LocalMux I__2641 (
            .O(N__12700),
            .I(beamYZ0Z_2));
    LocalMux I__2640 (
            .O(N__12695),
            .I(beamYZ0Z_2));
    InMux I__2639 (
            .O(N__12676),
            .I(un21_beamy_cry_1));
    CascadeMux I__2638 (
            .O(N__12673),
            .I(N__12666));
    CascadeMux I__2637 (
            .O(N__12672),
            .I(N__12661));
    CascadeMux I__2636 (
            .O(N__12671),
            .I(N__12657));
    CascadeMux I__2635 (
            .O(N__12670),
            .I(N__12645));
    CascadeMux I__2634 (
            .O(N__12669),
            .I(N__12639));
    InMux I__2633 (
            .O(N__12666),
            .I(N__12631));
    InMux I__2632 (
            .O(N__12665),
            .I(N__12631));
    InMux I__2631 (
            .O(N__12664),
            .I(N__12628));
    InMux I__2630 (
            .O(N__12661),
            .I(N__12625));
    InMux I__2629 (
            .O(N__12660),
            .I(N__12622));
    InMux I__2628 (
            .O(N__12657),
            .I(N__12617));
    InMux I__2627 (
            .O(N__12656),
            .I(N__12617));
    InMux I__2626 (
            .O(N__12655),
            .I(N__12608));
    InMux I__2625 (
            .O(N__12654),
            .I(N__12608));
    InMux I__2624 (
            .O(N__12653),
            .I(N__12608));
    InMux I__2623 (
            .O(N__12652),
            .I(N__12608));
    InMux I__2622 (
            .O(N__12651),
            .I(N__12601));
    InMux I__2621 (
            .O(N__12650),
            .I(N__12601));
    InMux I__2620 (
            .O(N__12649),
            .I(N__12601));
    InMux I__2619 (
            .O(N__12648),
            .I(N__12596));
    InMux I__2618 (
            .O(N__12645),
            .I(N__12589));
    InMux I__2617 (
            .O(N__12644),
            .I(N__12589));
    InMux I__2616 (
            .O(N__12643),
            .I(N__12589));
    InMux I__2615 (
            .O(N__12642),
            .I(N__12582));
    InMux I__2614 (
            .O(N__12639),
            .I(N__12575));
    InMux I__2613 (
            .O(N__12638),
            .I(N__12575));
    InMux I__2612 (
            .O(N__12637),
            .I(N__12575));
    InMux I__2611 (
            .O(N__12636),
            .I(N__12572));
    LocalMux I__2610 (
            .O(N__12631),
            .I(N__12563));
    LocalMux I__2609 (
            .O(N__12628),
            .I(N__12563));
    LocalMux I__2608 (
            .O(N__12625),
            .I(N__12563));
    LocalMux I__2607 (
            .O(N__12622),
            .I(N__12563));
    LocalMux I__2606 (
            .O(N__12617),
            .I(N__12556));
    LocalMux I__2605 (
            .O(N__12608),
            .I(N__12556));
    LocalMux I__2604 (
            .O(N__12601),
            .I(N__12556));
    InMux I__2603 (
            .O(N__12600),
            .I(N__12553));
    InMux I__2602 (
            .O(N__12599),
            .I(N__12550));
    LocalMux I__2601 (
            .O(N__12596),
            .I(N__12545));
    LocalMux I__2600 (
            .O(N__12589),
            .I(N__12545));
    InMux I__2599 (
            .O(N__12588),
            .I(N__12542));
    InMux I__2598 (
            .O(N__12587),
            .I(N__12539));
    CascadeMux I__2597 (
            .O(N__12586),
            .I(N__12535));
    InMux I__2596 (
            .O(N__12585),
            .I(N__12526));
    LocalMux I__2595 (
            .O(N__12582),
            .I(N__12523));
    LocalMux I__2594 (
            .O(N__12575),
            .I(N__12516));
    LocalMux I__2593 (
            .O(N__12572),
            .I(N__12516));
    Span4Mux_h I__2592 (
            .O(N__12563),
            .I(N__12516));
    Span4Mux_h I__2591 (
            .O(N__12556),
            .I(N__12513));
    LocalMux I__2590 (
            .O(N__12553),
            .I(N__12508));
    LocalMux I__2589 (
            .O(N__12550),
            .I(N__12508));
    Span4Mux_v I__2588 (
            .O(N__12545),
            .I(N__12501));
    LocalMux I__2587 (
            .O(N__12542),
            .I(N__12501));
    LocalMux I__2586 (
            .O(N__12539),
            .I(N__12501));
    InMux I__2585 (
            .O(N__12538),
            .I(N__12496));
    InMux I__2584 (
            .O(N__12535),
            .I(N__12496));
    InMux I__2583 (
            .O(N__12534),
            .I(N__12489));
    InMux I__2582 (
            .O(N__12533),
            .I(N__12489));
    InMux I__2581 (
            .O(N__12532),
            .I(N__12489));
    InMux I__2580 (
            .O(N__12531),
            .I(N__12482));
    InMux I__2579 (
            .O(N__12530),
            .I(N__12482));
    InMux I__2578 (
            .O(N__12529),
            .I(N__12482));
    LocalMux I__2577 (
            .O(N__12526),
            .I(beamYZ0Z_3));
    Odrv12 I__2576 (
            .O(N__12523),
            .I(beamYZ0Z_3));
    Odrv4 I__2575 (
            .O(N__12516),
            .I(beamYZ0Z_3));
    Odrv4 I__2574 (
            .O(N__12513),
            .I(beamYZ0Z_3));
    Odrv4 I__2573 (
            .O(N__12508),
            .I(beamYZ0Z_3));
    Odrv4 I__2572 (
            .O(N__12501),
            .I(beamYZ0Z_3));
    LocalMux I__2571 (
            .O(N__12496),
            .I(beamYZ0Z_3));
    LocalMux I__2570 (
            .O(N__12489),
            .I(beamYZ0Z_3));
    LocalMux I__2569 (
            .O(N__12482),
            .I(beamYZ0Z_3));
    InMux I__2568 (
            .O(N__12463),
            .I(un21_beamy_cry_2));
    InMux I__2567 (
            .O(N__12460),
            .I(N__12452));
    InMux I__2566 (
            .O(N__12459),
            .I(N__12447));
    InMux I__2565 (
            .O(N__12458),
            .I(N__12447));
    InMux I__2564 (
            .O(N__12457),
            .I(N__12442));
    InMux I__2563 (
            .O(N__12456),
            .I(N__12442));
    InMux I__2562 (
            .O(N__12455),
            .I(N__12429));
    LocalMux I__2561 (
            .O(N__12452),
            .I(N__12424));
    LocalMux I__2560 (
            .O(N__12447),
            .I(N__12424));
    LocalMux I__2559 (
            .O(N__12442),
            .I(N__12421));
    InMux I__2558 (
            .O(N__12441),
            .I(N__12418));
    InMux I__2557 (
            .O(N__12440),
            .I(N__12413));
    InMux I__2556 (
            .O(N__12439),
            .I(N__12413));
    InMux I__2555 (
            .O(N__12438),
            .I(N__12410));
    InMux I__2554 (
            .O(N__12437),
            .I(N__12407));
    CascadeMux I__2553 (
            .O(N__12436),
            .I(N__12402));
    CascadeMux I__2552 (
            .O(N__12435),
            .I(N__12399));
    CascadeMux I__2551 (
            .O(N__12434),
            .I(N__12395));
    InMux I__2550 (
            .O(N__12433),
            .I(N__12391));
    InMux I__2549 (
            .O(N__12432),
            .I(N__12388));
    LocalMux I__2548 (
            .O(N__12429),
            .I(N__12385));
    Span4Mux_h I__2547 (
            .O(N__12424),
            .I(N__12382));
    Span4Mux_v I__2546 (
            .O(N__12421),
            .I(N__12377));
    LocalMux I__2545 (
            .O(N__12418),
            .I(N__12377));
    LocalMux I__2544 (
            .O(N__12413),
            .I(N__12370));
    LocalMux I__2543 (
            .O(N__12410),
            .I(N__12370));
    LocalMux I__2542 (
            .O(N__12407),
            .I(N__12370));
    InMux I__2541 (
            .O(N__12406),
            .I(N__12367));
    InMux I__2540 (
            .O(N__12405),
            .I(N__12364));
    InMux I__2539 (
            .O(N__12402),
            .I(N__12357));
    InMux I__2538 (
            .O(N__12399),
            .I(N__12357));
    InMux I__2537 (
            .O(N__12398),
            .I(N__12357));
    InMux I__2536 (
            .O(N__12395),
            .I(N__12352));
    InMux I__2535 (
            .O(N__12394),
            .I(N__12352));
    LocalMux I__2534 (
            .O(N__12391),
            .I(beamYZ0Z_4));
    LocalMux I__2533 (
            .O(N__12388),
            .I(beamYZ0Z_4));
    Odrv12 I__2532 (
            .O(N__12385),
            .I(beamYZ0Z_4));
    Odrv4 I__2531 (
            .O(N__12382),
            .I(beamYZ0Z_4));
    Odrv4 I__2530 (
            .O(N__12377),
            .I(beamYZ0Z_4));
    Odrv4 I__2529 (
            .O(N__12370),
            .I(beamYZ0Z_4));
    LocalMux I__2528 (
            .O(N__12367),
            .I(beamYZ0Z_4));
    LocalMux I__2527 (
            .O(N__12364),
            .I(beamYZ0Z_4));
    LocalMux I__2526 (
            .O(N__12357),
            .I(beamYZ0Z_4));
    LocalMux I__2525 (
            .O(N__12352),
            .I(beamYZ0Z_4));
    InMux I__2524 (
            .O(N__12331),
            .I(un21_beamy_cry_3));
    InMux I__2523 (
            .O(N__12328),
            .I(N__12325));
    LocalMux I__2522 (
            .O(N__12325),
            .I(N__12318));
    InMux I__2521 (
            .O(N__12324),
            .I(N__12315));
    InMux I__2520 (
            .O(N__12323),
            .I(N__12310));
    InMux I__2519 (
            .O(N__12322),
            .I(N__12310));
    InMux I__2518 (
            .O(N__12321),
            .I(N__12299));
    Span4Mux_h I__2517 (
            .O(N__12318),
            .I(N__12296));
    LocalMux I__2516 (
            .O(N__12315),
            .I(N__12293));
    LocalMux I__2515 (
            .O(N__12310),
            .I(N__12290));
    InMux I__2514 (
            .O(N__12309),
            .I(N__12285));
    InMux I__2513 (
            .O(N__12308),
            .I(N__12285));
    InMux I__2512 (
            .O(N__12307),
            .I(N__12280));
    InMux I__2511 (
            .O(N__12306),
            .I(N__12280));
    InMux I__2510 (
            .O(N__12305),
            .I(N__12271));
    InMux I__2509 (
            .O(N__12304),
            .I(N__12271));
    InMux I__2508 (
            .O(N__12303),
            .I(N__12271));
    InMux I__2507 (
            .O(N__12302),
            .I(N__12271));
    LocalMux I__2506 (
            .O(N__12299),
            .I(beamYZ0Z_5));
    Odrv4 I__2505 (
            .O(N__12296),
            .I(beamYZ0Z_5));
    Odrv12 I__2504 (
            .O(N__12293),
            .I(beamYZ0Z_5));
    Odrv4 I__2503 (
            .O(N__12290),
            .I(beamYZ0Z_5));
    LocalMux I__2502 (
            .O(N__12285),
            .I(beamYZ0Z_5));
    LocalMux I__2501 (
            .O(N__12280),
            .I(beamYZ0Z_5));
    LocalMux I__2500 (
            .O(N__12271),
            .I(beamYZ0Z_5));
    InMux I__2499 (
            .O(N__12256),
            .I(un21_beamy_cry_4));
    CascadeMux I__2498 (
            .O(N__12253),
            .I(N__12250));
    InMux I__2497 (
            .O(N__12250),
            .I(N__12247));
    LocalMux I__2496 (
            .O(N__12247),
            .I(N__12244));
    Span4Mux_h I__2495 (
            .O(N__12244),
            .I(N__12237));
    InMux I__2494 (
            .O(N__12243),
            .I(N__12234));
    InMux I__2493 (
            .O(N__12242),
            .I(N__12229));
    InMux I__2492 (
            .O(N__12241),
            .I(N__12229));
    InMux I__2491 (
            .O(N__12240),
            .I(N__12219));
    Span4Mux_s3_h I__2490 (
            .O(N__12237),
            .I(N__12216));
    LocalMux I__2489 (
            .O(N__12234),
            .I(N__12213));
    LocalMux I__2488 (
            .O(N__12229),
            .I(N__12210));
    InMux I__2487 (
            .O(N__12228),
            .I(N__12205));
    InMux I__2486 (
            .O(N__12227),
            .I(N__12205));
    InMux I__2485 (
            .O(N__12226),
            .I(N__12202));
    InMux I__2484 (
            .O(N__12225),
            .I(N__12199));
    InMux I__2483 (
            .O(N__12224),
            .I(N__12192));
    InMux I__2482 (
            .O(N__12223),
            .I(N__12192));
    InMux I__2481 (
            .O(N__12222),
            .I(N__12192));
    LocalMux I__2480 (
            .O(N__12219),
            .I(beamYZ0Z_6));
    Odrv4 I__2479 (
            .O(N__12216),
            .I(beamYZ0Z_6));
    Odrv12 I__2478 (
            .O(N__12213),
            .I(beamYZ0Z_6));
    Odrv4 I__2477 (
            .O(N__12210),
            .I(beamYZ0Z_6));
    LocalMux I__2476 (
            .O(N__12205),
            .I(beamYZ0Z_6));
    LocalMux I__2475 (
            .O(N__12202),
            .I(beamYZ0Z_6));
    LocalMux I__2474 (
            .O(N__12199),
            .I(beamYZ0Z_6));
    LocalMux I__2473 (
            .O(N__12192),
            .I(beamYZ0Z_6));
    InMux I__2472 (
            .O(N__12175),
            .I(un21_beamy_cry_5));
    InMux I__2471 (
            .O(N__12172),
            .I(N__12166));
    InMux I__2470 (
            .O(N__12171),
            .I(N__12166));
    LocalMux I__2469 (
            .O(N__12166),
            .I(N__12160));
    InMux I__2468 (
            .O(N__12165),
            .I(N__12157));
    InMux I__2467 (
            .O(N__12164),
            .I(N__12154));
    InMux I__2466 (
            .O(N__12163),
            .I(N__12145));
    Span4Mux_h I__2465 (
            .O(N__12160),
            .I(N__12142));
    LocalMux I__2464 (
            .O(N__12157),
            .I(N__12137));
    LocalMux I__2463 (
            .O(N__12154),
            .I(N__12137));
    InMux I__2462 (
            .O(N__12153),
            .I(N__12132));
    InMux I__2461 (
            .O(N__12152),
            .I(N__12132));
    InMux I__2460 (
            .O(N__12151),
            .I(N__12127));
    InMux I__2459 (
            .O(N__12150),
            .I(N__12127));
    InMux I__2458 (
            .O(N__12149),
            .I(N__12122));
    InMux I__2457 (
            .O(N__12148),
            .I(N__12122));
    LocalMux I__2456 (
            .O(N__12145),
            .I(beamYZ0Z_7));
    Odrv4 I__2455 (
            .O(N__12142),
            .I(beamYZ0Z_7));
    Odrv12 I__2454 (
            .O(N__12137),
            .I(beamYZ0Z_7));
    LocalMux I__2453 (
            .O(N__12132),
            .I(beamYZ0Z_7));
    LocalMux I__2452 (
            .O(N__12127),
            .I(beamYZ0Z_7));
    LocalMux I__2451 (
            .O(N__12122),
            .I(beamYZ0Z_7));
    InMux I__2450 (
            .O(N__12109),
            .I(un21_beamy_cry_6));
    InMux I__2449 (
            .O(N__12106),
            .I(N__12099));
    InMux I__2448 (
            .O(N__12105),
            .I(N__12094));
    InMux I__2447 (
            .O(N__12104),
            .I(N__12094));
    InMux I__2446 (
            .O(N__12103),
            .I(N__12089));
    InMux I__2445 (
            .O(N__12102),
            .I(N__12086));
    LocalMux I__2444 (
            .O(N__12099),
            .I(N__12081));
    LocalMux I__2443 (
            .O(N__12094),
            .I(N__12081));
    CascadeMux I__2442 (
            .O(N__12093),
            .I(N__12073));
    InMux I__2441 (
            .O(N__12092),
            .I(N__12070));
    LocalMux I__2440 (
            .O(N__12089),
            .I(N__12067));
    LocalMux I__2439 (
            .O(N__12086),
            .I(N__12064));
    Span4Mux_h I__2438 (
            .O(N__12081),
            .I(N__12061));
    InMux I__2437 (
            .O(N__12080),
            .I(N__12058));
    InMux I__2436 (
            .O(N__12079),
            .I(N__12051));
    InMux I__2435 (
            .O(N__12078),
            .I(N__12051));
    InMux I__2434 (
            .O(N__12077),
            .I(N__12051));
    InMux I__2433 (
            .O(N__12076),
            .I(N__12046));
    InMux I__2432 (
            .O(N__12073),
            .I(N__12046));
    LocalMux I__2431 (
            .O(N__12070),
            .I(beamYZ0Z_8));
    Odrv4 I__2430 (
            .O(N__12067),
            .I(beamYZ0Z_8));
    Odrv12 I__2429 (
            .O(N__12064),
            .I(beamYZ0Z_8));
    Odrv4 I__2428 (
            .O(N__12061),
            .I(beamYZ0Z_8));
    LocalMux I__2427 (
            .O(N__12058),
            .I(beamYZ0Z_8));
    LocalMux I__2426 (
            .O(N__12051),
            .I(beamYZ0Z_8));
    LocalMux I__2425 (
            .O(N__12046),
            .I(beamYZ0Z_8));
    InMux I__2424 (
            .O(N__12031),
            .I(un21_beamy_cry_7));
    InMux I__2423 (
            .O(N__12028),
            .I(N__12025));
    LocalMux I__2422 (
            .O(N__12025),
            .I(un5_visibley_3_29));
    CascadeMux I__2421 (
            .O(N__12022),
            .I(g1_8_1_cascade_));
    CascadeMux I__2420 (
            .O(N__12019),
            .I(N__12015));
    InMux I__2419 (
            .O(N__12018),
            .I(N__12011));
    InMux I__2418 (
            .O(N__12015),
            .I(N__12006));
    InMux I__2417 (
            .O(N__12014),
            .I(N__12006));
    LocalMux I__2416 (
            .O(N__12011),
            .I(N__11999));
    LocalMux I__2415 (
            .O(N__12006),
            .I(N__11996));
    InMux I__2414 (
            .O(N__12005),
            .I(N__11985));
    InMux I__2413 (
            .O(N__12004),
            .I(N__11985));
    InMux I__2412 (
            .O(N__12003),
            .I(N__11985));
    InMux I__2411 (
            .O(N__12002),
            .I(N__11980));
    Span4Mux_h I__2410 (
            .O(N__11999),
            .I(N__11977));
    Span4Mux_h I__2409 (
            .O(N__11996),
            .I(N__11974));
    InMux I__2408 (
            .O(N__11995),
            .I(N__11967));
    InMux I__2407 (
            .O(N__11994),
            .I(N__11967));
    InMux I__2406 (
            .O(N__11993),
            .I(N__11967));
    InMux I__2405 (
            .O(N__11992),
            .I(N__11964));
    LocalMux I__2404 (
            .O(N__11985),
            .I(N__11961));
    InMux I__2403 (
            .O(N__11984),
            .I(N__11958));
    InMux I__2402 (
            .O(N__11983),
            .I(N__11955));
    LocalMux I__2401 (
            .O(N__11980),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    Odrv4 I__2400 (
            .O(N__11977),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    Odrv4 I__2399 (
            .O(N__11974),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    LocalMux I__2398 (
            .O(N__11967),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    LocalMux I__2397 (
            .O(N__11964),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    Odrv4 I__2396 (
            .O(N__11961),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    LocalMux I__2395 (
            .O(N__11958),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    LocalMux I__2394 (
            .O(N__11955),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    InMux I__2393 (
            .O(N__11938),
            .I(N__11935));
    LocalMux I__2392 (
            .O(N__11935),
            .I(N__11932));
    Odrv4 I__2391 (
            .O(N__11932),
            .I(g1_3_0));
    CascadeMux I__2390 (
            .O(N__11929),
            .I(N__11926));
    InMux I__2389 (
            .O(N__11926),
            .I(N__11923));
    LocalMux I__2388 (
            .O(N__11923),
            .I(N__11920));
    Odrv12 I__2387 (
            .O(N__11920),
            .I(un5_visibley_1_0_28));
    CascadeMux I__2386 (
            .O(N__11917),
            .I(beamY_RNIJ0H2Z0Z_4_cascade_));
    CascadeMux I__2385 (
            .O(N__11914),
            .I(N__11911));
    InMux I__2384 (
            .O(N__11911),
            .I(N__11908));
    LocalMux I__2383 (
            .O(N__11908),
            .I(un5_visibley_c5));
    InMux I__2382 (
            .O(N__11905),
            .I(N__11902));
    LocalMux I__2381 (
            .O(N__11902),
            .I(un5_visibley_c6_0_0_0));
    CascadeMux I__2380 (
            .O(N__11899),
            .I(un5_visibley_c6_0_0_0_cascade_));
    InMux I__2379 (
            .O(N__11896),
            .I(N__11892));
    InMux I__2378 (
            .O(N__11895),
            .I(N__11889));
    LocalMux I__2377 (
            .O(N__11892),
            .I(un5_visibley_c3));
    LocalMux I__2376 (
            .O(N__11889),
            .I(un5_visibley_c3));
    CascadeMux I__2375 (
            .O(N__11884),
            .I(un19_slaveselectlt5_0_cascade_));
    InMux I__2374 (
            .O(N__11881),
            .I(N__11875));
    InMux I__2373 (
            .O(N__11880),
            .I(N__11875));
    LocalMux I__2372 (
            .O(N__11875),
            .I(un19_slaveselectlt5_0));
    CascadeMux I__2371 (
            .O(N__11872),
            .I(counter_RNI4HQB1Z0Z_5_cascade_));
    CascadeMux I__2370 (
            .O(N__11869),
            .I(beamY_RNI4FVGVZ0Z_4_cascade_));
    InMux I__2369 (
            .O(N__11866),
            .I(N__11857));
    InMux I__2368 (
            .O(N__11865),
            .I(N__11857));
    InMux I__2367 (
            .O(N__11864),
            .I(N__11852));
    InMux I__2366 (
            .O(N__11863),
            .I(N__11852));
    InMux I__2365 (
            .O(N__11862),
            .I(N__11849));
    LocalMux I__2364 (
            .O(N__11857),
            .I(N__11846));
    LocalMux I__2363 (
            .O(N__11852),
            .I(N__11843));
    LocalMux I__2362 (
            .O(N__11849),
            .I(N__11840));
    Span4Mux_h I__2361 (
            .O(N__11846),
            .I(N__11837));
    Span4Mux_h I__2360 (
            .O(N__11843),
            .I(N__11834));
    Odrv4 I__2359 (
            .O(N__11840),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    Odrv4 I__2358 (
            .O(N__11837),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    Odrv4 I__2357 (
            .O(N__11834),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    InMux I__2356 (
            .O(N__11827),
            .I(N__11824));
    LocalMux I__2355 (
            .O(N__11824),
            .I(N__11821));
    Span4Mux_h I__2354 (
            .O(N__11821),
            .I(N__11818));
    Odrv4 I__2353 (
            .O(N__11818),
            .I(N_596_2));
    CascadeMux I__2352 (
            .O(N__11815),
            .I(un5_visibley_4_28_cascade_));
    CascadeMux I__2351 (
            .O(N__11812),
            .I(N__11809));
    InMux I__2350 (
            .O(N__11809),
            .I(N__11805));
    CascadeMux I__2349 (
            .O(N__11808),
            .I(N__11802));
    LocalMux I__2348 (
            .O(N__11805),
            .I(N__11799));
    InMux I__2347 (
            .O(N__11802),
            .I(N__11796));
    Span4Mux_h I__2346 (
            .O(N__11799),
            .I(N__11793));
    LocalMux I__2345 (
            .O(N__11796),
            .I(content_ram12_0));
    Odrv4 I__2344 (
            .O(N__11793),
            .I(content_ram12_0));
    InMux I__2343 (
            .O(N__11788),
            .I(N__11785));
    LocalMux I__2342 (
            .O(N__11785),
            .I(content_awe0_0_a2_0));
    CascadeMux I__2341 (
            .O(N__11782),
            .I(content_awe0_0_a2_0_cascade_));
    InMux I__2340 (
            .O(N__11779),
            .I(N__11776));
    LocalMux I__2339 (
            .O(N__11776),
            .I(N__11772));
    InMux I__2338 (
            .O(N__11775),
            .I(N__11769));
    Span4Mux_h I__2337 (
            .O(N__11772),
            .I(N__11766));
    LocalMux I__2336 (
            .O(N__11769),
            .I(content_ram4_0));
    Odrv4 I__2335 (
            .O(N__11766),
            .I(content_ram4_0));
    InMux I__2334 (
            .O(N__11761),
            .I(N__11752));
    InMux I__2333 (
            .O(N__11760),
            .I(N__11752));
    InMux I__2332 (
            .O(N__11759),
            .I(N__11752));
    LocalMux I__2331 (
            .O(N__11752),
            .I(content_N_36));
    CascadeMux I__2330 (
            .O(N__11749),
            .I(content_N_36_cascade_));
    CascadeMux I__2329 (
            .O(N__11746),
            .I(content_awe7_1_cascade_));
    InMux I__2328 (
            .O(N__11743),
            .I(N__11739));
    InMux I__2327 (
            .O(N__11742),
            .I(N__11736));
    LocalMux I__2326 (
            .O(N__11739),
            .I(N__11733));
    LocalMux I__2325 (
            .O(N__11736),
            .I(content_ram6_0));
    Odrv4 I__2324 (
            .O(N__11733),
            .I(content_ram6_0));
    InMux I__2323 (
            .O(N__11728),
            .I(N__11725));
    LocalMux I__2322 (
            .O(N__11725),
            .I(content_awe7_1));
    CascadeMux I__2321 (
            .O(N__11722),
            .I(N__11718));
    InMux I__2320 (
            .O(N__11721),
            .I(N__11715));
    InMux I__2319 (
            .O(N__11718),
            .I(N__11712));
    LocalMux I__2318 (
            .O(N__11715),
            .I(N__11709));
    LocalMux I__2317 (
            .O(N__11712),
            .I(N__11704));
    Span4Mux_v I__2316 (
            .O(N__11709),
            .I(N__11704));
    Odrv4 I__2315 (
            .O(N__11704),
            .I(content_ram7_0));
    SRMux I__2314 (
            .O(N__11701),
            .I(N__11698));
    LocalMux I__2313 (
            .O(N__11698),
            .I(nCS1_0_sqmuxa));
    CascadeMux I__2312 (
            .O(N__11695),
            .I(content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_));
    CascadeMux I__2311 (
            .O(N__11692),
            .I(N__11688));
    CascadeMux I__2310 (
            .O(N__11691),
            .I(N__11685));
    InMux I__2309 (
            .O(N__11688),
            .I(N__11679));
    InMux I__2308 (
            .O(N__11685),
            .I(N__11679));
    CascadeMux I__2307 (
            .O(N__11684),
            .I(N__11676));
    LocalMux I__2306 (
            .O(N__11679),
            .I(N__11673));
    InMux I__2305 (
            .O(N__11676),
            .I(N__11670));
    Span4Mux_h I__2304 (
            .O(N__11673),
            .I(N__11665));
    LocalMux I__2303 (
            .O(N__11670),
            .I(N__11665));
    Span4Mux_v I__2302 (
            .O(N__11665),
            .I(N__11662));
    Odrv4 I__2301 (
            .O(N__11662),
            .I(content_N_19));
    InMux I__2300 (
            .O(N__11659),
            .I(N__11654));
    InMux I__2299 (
            .O(N__11658),
            .I(N__11647));
    InMux I__2298 (
            .O(N__11657),
            .I(N__11647));
    LocalMux I__2297 (
            .O(N__11654),
            .I(N__11638));
    InMux I__2296 (
            .O(N__11653),
            .I(N__11633));
    InMux I__2295 (
            .O(N__11652),
            .I(N__11633));
    LocalMux I__2294 (
            .O(N__11647),
            .I(N__11630));
    InMux I__2293 (
            .O(N__11646),
            .I(N__11623));
    InMux I__2292 (
            .O(N__11645),
            .I(N__11623));
    InMux I__2291 (
            .O(N__11644),
            .I(N__11623));
    InMux I__2290 (
            .O(N__11643),
            .I(N__11620));
    InMux I__2289 (
            .O(N__11642),
            .I(N__11617));
    InMux I__2288 (
            .O(N__11641),
            .I(N__11614));
    Odrv4 I__2287 (
            .O(N__11638),
            .I(content_column_1_i_2_2));
    LocalMux I__2286 (
            .O(N__11633),
            .I(content_column_1_i_2_2));
    Odrv4 I__2285 (
            .O(N__11630),
            .I(content_column_1_i_2_2));
    LocalMux I__2284 (
            .O(N__11623),
            .I(content_column_1_i_2_2));
    LocalMux I__2283 (
            .O(N__11620),
            .I(content_column_1_i_2_2));
    LocalMux I__2282 (
            .O(N__11617),
            .I(content_column_1_i_2_2));
    LocalMux I__2281 (
            .O(N__11614),
            .I(content_column_1_i_2_2));
    CascadeMux I__2280 (
            .O(N__11599),
            .I(N__11594));
    CascadeMux I__2279 (
            .O(N__11598),
            .I(N__11591));
    InMux I__2278 (
            .O(N__11597),
            .I(N__11586));
    InMux I__2277 (
            .O(N__11594),
            .I(N__11581));
    InMux I__2276 (
            .O(N__11591),
            .I(N__11581));
    InMux I__2275 (
            .O(N__11590),
            .I(N__11576));
    InMux I__2274 (
            .O(N__11589),
            .I(N__11576));
    LocalMux I__2273 (
            .O(N__11586),
            .I(N__11567));
    LocalMux I__2272 (
            .O(N__11581),
            .I(N__11564));
    LocalMux I__2271 (
            .O(N__11576),
            .I(N__11561));
    InMux I__2270 (
            .O(N__11575),
            .I(N__11552));
    InMux I__2269 (
            .O(N__11574),
            .I(N__11552));
    InMux I__2268 (
            .O(N__11573),
            .I(N__11552));
    InMux I__2267 (
            .O(N__11572),
            .I(N__11552));
    InMux I__2266 (
            .O(N__11571),
            .I(N__11549));
    InMux I__2265 (
            .O(N__11570),
            .I(N__11546));
    Odrv4 I__2264 (
            .O(N__11567),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    Odrv12 I__2263 (
            .O(N__11564),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    Odrv4 I__2262 (
            .O(N__11561),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    LocalMux I__2261 (
            .O(N__11552),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    LocalMux I__2260 (
            .O(N__11549),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    LocalMux I__2259 (
            .O(N__11546),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    InMux I__2258 (
            .O(N__11533),
            .I(N__11530));
    LocalMux I__2257 (
            .O(N__11530),
            .I(content_content_ram10__e_0_RNIOLNMN1Z0Z_0));
    CascadeMux I__2256 (
            .O(N__11527),
            .I(N__11522));
    InMux I__2255 (
            .O(N__11526),
            .I(N__11517));
    InMux I__2254 (
            .O(N__11525),
            .I(N__11517));
    InMux I__2253 (
            .O(N__11522),
            .I(N__11514));
    LocalMux I__2252 (
            .O(N__11517),
            .I(N__11511));
    LocalMux I__2251 (
            .O(N__11514),
            .I(content_ram3_0));
    Odrv4 I__2250 (
            .O(N__11511),
            .I(content_ram3_0));
    CEMux I__2249 (
            .O(N__11506),
            .I(N__11503));
    LocalMux I__2248 (
            .O(N__11503),
            .I(content_awe9));
    CascadeMux I__2247 (
            .O(N__11500),
            .I(N__11496));
    InMux I__2246 (
            .O(N__11499),
            .I(N__11493));
    InMux I__2245 (
            .O(N__11496),
            .I(N__11490));
    LocalMux I__2244 (
            .O(N__11493),
            .I(N__11487));
    LocalMux I__2243 (
            .O(N__11490),
            .I(content_ram0_0));
    Odrv4 I__2242 (
            .O(N__11487),
            .I(content_ram0_0));
    CEMux I__2241 (
            .O(N__11482),
            .I(N__11479));
    LocalMux I__2240 (
            .O(N__11479),
            .I(N__11476));
    Span4Mux_h I__2239 (
            .O(N__11476),
            .I(N__11473));
    Odrv4 I__2238 (
            .O(N__11473),
            .I(content_awe8));
    CEMux I__2237 (
            .O(N__11470),
            .I(N__11467));
    LocalMux I__2236 (
            .O(N__11467),
            .I(N__11464));
    Odrv4 I__2235 (
            .O(N__11464),
            .I(content_awe11));
    CascadeMux I__2234 (
            .O(N__11461),
            .I(N__11457));
    InMux I__2233 (
            .O(N__11460),
            .I(N__11454));
    InMux I__2232 (
            .O(N__11457),
            .I(N__11451));
    LocalMux I__2231 (
            .O(N__11454),
            .I(N__11448));
    LocalMux I__2230 (
            .O(N__11451),
            .I(content_ram5_0));
    Odrv4 I__2229 (
            .O(N__11448),
            .I(content_ram5_0));
    InMux I__2228 (
            .O(N__11443),
            .I(N__11440));
    LocalMux I__2227 (
            .O(N__11440),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__2226 (
            .O(N__11437),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__2225 (
            .O(N__11434),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__2224 (
            .O(N__11431),
            .I(N__11427));
    InMux I__2223 (
            .O(N__11430),
            .I(N__11418));
    InMux I__2222 (
            .O(N__11427),
            .I(N__11418));
    InMux I__2221 (
            .O(N__11426),
            .I(N__11418));
    InMux I__2220 (
            .O(N__11425),
            .I(N__11415));
    LocalMux I__2219 (
            .O(N__11418),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4));
    LocalMux I__2218 (
            .O(N__11415),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4));
    CascadeMux I__2217 (
            .O(N__11410),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_));
    InMux I__2216 (
            .O(N__11407),
            .I(N__11404));
    LocalMux I__2215 (
            .O(N__11404),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__2214 (
            .O(N__11401),
            .I(N__11398));
    LocalMux I__2213 (
            .O(N__11398),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54));
    CascadeMux I__2212 (
            .O(N__11395),
            .I(N__11392));
    InMux I__2211 (
            .O(N__11392),
            .I(N__11389));
    LocalMux I__2210 (
            .O(N__11389),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0));
    CascadeMux I__2209 (
            .O(N__11386),
            .I(N__11383));
    InMux I__2208 (
            .O(N__11383),
            .I(N__11380));
    LocalMux I__2207 (
            .O(N__11380),
            .I(N__11377));
    Odrv12 I__2206 (
            .O(N__11377),
            .I(CO4_1));
    InMux I__2205 (
            .O(N__11374),
            .I(N__11371));
    LocalMux I__2204 (
            .O(N__11371),
            .I(N__11368));
    Odrv12 I__2203 (
            .O(N__11368),
            .I(row_1_if_generate_plus_mult1_un47_sum_cZ0Z5));
    InMux I__2202 (
            .O(N__11365),
            .I(N__11362));
    LocalMux I__2201 (
            .O(N__11362),
            .I(N__11359));
    Span4Mux_h I__2200 (
            .O(N__11359),
            .I(N__11356));
    Odrv4 I__2199 (
            .O(N__11356),
            .I(content_ram8_0));
    CascadeMux I__2198 (
            .O(N__11353),
            .I(N__11350));
    InMux I__2197 (
            .O(N__11350),
            .I(N__11347));
    LocalMux I__2196 (
            .O(N__11347),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28));
    InMux I__2195 (
            .O(N__11344),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__2194 (
            .O(N__11341),
            .I(N__11338));
    LocalMux I__2193 (
            .O(N__11338),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__2192 (
            .O(N__11335),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__2191 (
            .O(N__11332),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__2190 (
            .O(N__11329),
            .I(N__11324));
    CascadeMux I__2189 (
            .O(N__11328),
            .I(N__11320));
    InMux I__2188 (
            .O(N__11327),
            .I(N__11316));
    InMux I__2187 (
            .O(N__11324),
            .I(N__11307));
    InMux I__2186 (
            .O(N__11323),
            .I(N__11307));
    InMux I__2185 (
            .O(N__11320),
            .I(N__11307));
    InMux I__2184 (
            .O(N__11319),
            .I(N__11307));
    LocalMux I__2183 (
            .O(N__11316),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0));
    LocalMux I__2182 (
            .O(N__11307),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0));
    CascadeMux I__2181 (
            .O(N__11302),
            .I(N__11299));
    InMux I__2180 (
            .O(N__11299),
            .I(N__11296));
    LocalMux I__2179 (
            .O(N__11296),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__2178 (
            .O(N__11293),
            .I(N__11290));
    LocalMux I__2177 (
            .O(N__11290),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2));
    InMux I__2176 (
            .O(N__11287),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__2175 (
            .O(N__11284),
            .I(N__11281));
    InMux I__2174 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__2173 (
            .O(N__11278),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193));
    InMux I__2172 (
            .O(N__11275),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__2171 (
            .O(N__11272),
            .I(N__11269));
    InMux I__2170 (
            .O(N__11269),
            .I(N__11266));
    LocalMux I__2169 (
            .O(N__11266),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3));
    InMux I__2168 (
            .O(N__11263),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2167 (
            .O(N__11260),
            .I(un5_beamx_2_0_cascade_));
    InMux I__2166 (
            .O(N__11257),
            .I(N__11254));
    LocalMux I__2165 (
            .O(N__11254),
            .I(un5_beamx_3));
    CascadeMux I__2164 (
            .O(N__11251),
            .I(un5_visibley_ac0_11_0_1_cascade_));
    CascadeMux I__2163 (
            .O(N__11248),
            .I(N__11245));
    InMux I__2162 (
            .O(N__11245),
            .I(N__11242));
    LocalMux I__2161 (
            .O(N__11242),
            .I(beamY_RNI8325_0Z0Z_6));
    CascadeMux I__2160 (
            .O(N__11239),
            .I(N__11235));
    InMux I__2159 (
            .O(N__11238),
            .I(N__11230));
    InMux I__2158 (
            .O(N__11235),
            .I(N__11230));
    LocalMux I__2157 (
            .O(N__11230),
            .I(N__11225));
    InMux I__2156 (
            .O(N__11229),
            .I(N__11222));
    InMux I__2155 (
            .O(N__11228),
            .I(N__11219));
    Odrv4 I__2154 (
            .O(N__11225),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    LocalMux I__2153 (
            .O(N__11222),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    LocalMux I__2152 (
            .O(N__11219),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    CascadeMux I__2151 (
            .O(N__11212),
            .I(N__11209));
    InMux I__2150 (
            .O(N__11209),
            .I(N__11206));
    LocalMux I__2149 (
            .O(N__11206),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4));
    InMux I__2148 (
            .O(N__11203),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__2147 (
            .O(N__11200),
            .I(N__11197));
    LocalMux I__2146 (
            .O(N__11197),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7));
    InMux I__2145 (
            .O(N__11194),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__2144 (
            .O(N__11191),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_));
    InMux I__2143 (
            .O(N__11188),
            .I(N__11185));
    LocalMux I__2142 (
            .O(N__11185),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0));
    CascadeMux I__2141 (
            .O(N__11182),
            .I(N__11176));
    InMux I__2140 (
            .O(N__11181),
            .I(N__11171));
    InMux I__2139 (
            .O(N__11180),
            .I(N__11171));
    InMux I__2138 (
            .O(N__11179),
            .I(N__11168));
    InMux I__2137 (
            .O(N__11176),
            .I(N__11164));
    LocalMux I__2136 (
            .O(N__11171),
            .I(N__11159));
    LocalMux I__2135 (
            .O(N__11168),
            .I(N__11159));
    InMux I__2134 (
            .O(N__11167),
            .I(N__11156));
    LocalMux I__2133 (
            .O(N__11164),
            .I(N__11152));
    Span4Mux_v I__2132 (
            .O(N__11159),
            .I(N__11147));
    LocalMux I__2131 (
            .O(N__11156),
            .I(N__11147));
    InMux I__2130 (
            .O(N__11155),
            .I(N__11144));
    Odrv4 I__2129 (
            .O(N__11152),
            .I(beamY_RNIVMI9D5Z0Z_3));
    Odrv4 I__2128 (
            .O(N__11147),
            .I(beamY_RNIVMI9D5Z0Z_3));
    LocalMux I__2127 (
            .O(N__11144),
            .I(beamY_RNIVMI9D5Z0Z_3));
    CascadeMux I__2126 (
            .O(N__11137),
            .I(N__11134));
    InMux I__2125 (
            .O(N__11134),
            .I(N__11131));
    LocalMux I__2124 (
            .O(N__11131),
            .I(un5_visibley_1_29));
    CascadeMux I__2123 (
            .O(N__11128),
            .I(N__11124));
    CascadeMux I__2122 (
            .O(N__11127),
            .I(N__11120));
    InMux I__2121 (
            .O(N__11124),
            .I(N__11116));
    InMux I__2120 (
            .O(N__11123),
            .I(N__11111));
    InMux I__2119 (
            .O(N__11120),
            .I(N__11111));
    CascadeMux I__2118 (
            .O(N__11119),
            .I(N__11106));
    LocalMux I__2117 (
            .O(N__11116),
            .I(N__11103));
    LocalMux I__2116 (
            .O(N__11111),
            .I(N__11100));
    InMux I__2115 (
            .O(N__11110),
            .I(N__11095));
    InMux I__2114 (
            .O(N__11109),
            .I(N__11095));
    InMux I__2113 (
            .O(N__11106),
            .I(N__11092));
    Span4Mux_v I__2112 (
            .O(N__11103),
            .I(N__11085));
    Span4Mux_v I__2111 (
            .O(N__11100),
            .I(N__11085));
    LocalMux I__2110 (
            .O(N__11095),
            .I(N__11085));
    LocalMux I__2109 (
            .O(N__11092),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    Odrv4 I__2108 (
            .O(N__11085),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    CascadeMux I__2107 (
            .O(N__11080),
            .I(beamY_RNI8325Z0Z_6_cascade_));
    CascadeMux I__2106 (
            .O(N__11077),
            .I(un5_visibley_c5_cascade_));
    InMux I__2105 (
            .O(N__11074),
            .I(N__11071));
    LocalMux I__2104 (
            .O(N__11071),
            .I(un1_beamylto9_1));
    CascadeMux I__2103 (
            .O(N__11068),
            .I(un5_visibley_c3_cascade_));
    CascadeMux I__2102 (
            .O(N__11065),
            .I(content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_));
    InMux I__2101 (
            .O(N__11062),
            .I(N__11059));
    LocalMux I__2100 (
            .O(N__11059),
            .I(content_content_ram9__e_0_RNIFBHPN1Z0Z_0));
    CascadeMux I__2099 (
            .O(N__11056),
            .I(N__11053));
    InMux I__2098 (
            .O(N__11053),
            .I(N__11050));
    LocalMux I__2097 (
            .O(N__11050),
            .I(content_content_ram5__RNIEM2QF3Z0Z_0));
    CascadeMux I__2096 (
            .O(N__11047),
            .I(N__11044));
    InMux I__2095 (
            .O(N__11044),
            .I(N__11038));
    InMux I__2094 (
            .O(N__11043),
            .I(N__11038));
    LocalMux I__2093 (
            .O(N__11038),
            .I(content_ram9_0));
    CascadeMux I__2092 (
            .O(N__11035),
            .I(N__11031));
    CascadeMux I__2091 (
            .O(N__11034),
            .I(N__11028));
    InMux I__2090 (
            .O(N__11031),
            .I(N__11023));
    InMux I__2089 (
            .O(N__11028),
            .I(N__11023));
    LocalMux I__2088 (
            .O(N__11023),
            .I(content_ram11_0));
    IoInMux I__2087 (
            .O(N__11020),
            .I(N__11016));
    IoInMux I__2086 (
            .O(N__11019),
            .I(N__11013));
    LocalMux I__2085 (
            .O(N__11016),
            .I(N__11008));
    LocalMux I__2084 (
            .O(N__11013),
            .I(N__11008));
    IoSpan4Mux I__2083 (
            .O(N__11008),
            .I(N__11005));
    Span4Mux_s2_h I__2082 (
            .O(N__11005),
            .I(N__11001));
    InMux I__2081 (
            .O(N__11004),
            .I(N__10998));
    Odrv4 I__2080 (
            .O(N__11001),
            .I(nCS1_c));
    LocalMux I__2079 (
            .O(N__10998),
            .I(nCS1_c));
    InMux I__2078 (
            .O(N__10993),
            .I(N__10987));
    InMux I__2077 (
            .O(N__10992),
            .I(N__10987));
    LocalMux I__2076 (
            .O(N__10987),
            .I(un5_visibley_2_28));
    InMux I__2075 (
            .O(N__10984),
            .I(N__10981));
    LocalMux I__2074 (
            .O(N__10981),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__2073 (
            .O(N__10978),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__2072 (
            .O(N__10975),
            .I(N__10969));
    InMux I__2071 (
            .O(N__10974),
            .I(N__10969));
    LocalMux I__2070 (
            .O(N__10969),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0));
    InMux I__2069 (
            .O(N__10966),
            .I(N__10963));
    LocalMux I__2068 (
            .O(N__10963),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0));
    InMux I__2067 (
            .O(N__10960),
            .I(N__10957));
    LocalMux I__2066 (
            .O(N__10957),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4));
    CascadeMux I__2065 (
            .O(N__10954),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_));
    InMux I__2064 (
            .O(N__10951),
            .I(N__10947));
    InMux I__2063 (
            .O(N__10950),
            .I(N__10944));
    LocalMux I__2062 (
            .O(N__10947),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0));
    LocalMux I__2061 (
            .O(N__10944),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0));
    InMux I__2060 (
            .O(N__10939),
            .I(N__10936));
    LocalMux I__2059 (
            .O(N__10936),
            .I(N__10933));
    Span4Mux_h I__2058 (
            .O(N__10933),
            .I(N__10930));
    Odrv4 I__2057 (
            .O(N__10930),
            .I(chessboardpixel_un178_pixel_26));
    InMux I__2056 (
            .O(N__10927),
            .I(N__10924));
    LocalMux I__2055 (
            .O(N__10924),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__2054 (
            .O(N__10921),
            .I(N__10918));
    LocalMux I__2053 (
            .O(N__10918),
            .I(N__10915));
    Span4Mux_h I__2052 (
            .O(N__10915),
            .I(N__10912));
    Odrv4 I__2051 (
            .O(N__10912),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z5));
    CascadeMux I__2050 (
            .O(N__10909),
            .I(N__10906));
    InMux I__2049 (
            .O(N__10906),
            .I(N__10903));
    LocalMux I__2048 (
            .O(N__10903),
            .I(row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3));
    InMux I__2047 (
            .O(N__10900),
            .I(N__10896));
    InMux I__2046 (
            .O(N__10899),
            .I(N__10893));
    LocalMux I__2045 (
            .O(N__10896),
            .I(N__10890));
    LocalMux I__2044 (
            .O(N__10893),
            .I(N__10887));
    Span4Mux_h I__2043 (
            .O(N__10890),
            .I(N__10882));
    Span4Mux_h I__2042 (
            .O(N__10887),
            .I(N__10879));
    InMux I__2041 (
            .O(N__10886),
            .I(N__10874));
    InMux I__2040 (
            .O(N__10885),
            .I(N__10874));
    Odrv4 I__2039 (
            .O(N__10882),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    Odrv4 I__2038 (
            .O(N__10879),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    LocalMux I__2037 (
            .O(N__10874),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    CascadeMux I__2036 (
            .O(N__10867),
            .I(row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_));
    InMux I__2035 (
            .O(N__10864),
            .I(N__10861));
    LocalMux I__2034 (
            .O(N__10861),
            .I(N__10858));
    Odrv4 I__2033 (
            .O(N__10858),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0));
    CascadeMux I__2032 (
            .O(N__10855),
            .I(chessboardpixel_un200_pixellto4_1_cascade_));
    InMux I__2031 (
            .O(N__10852),
            .I(N__10849));
    LocalMux I__2030 (
            .O(N__10849),
            .I(N__10846));
    Span4Mux_v I__2029 (
            .O(N__10846),
            .I(N__10843));
    Odrv4 I__2028 (
            .O(N__10843),
            .I(chessboardpixel_un200_pixellt10));
    CascadeMux I__2027 (
            .O(N__10840),
            .I(N__10835));
    InMux I__2026 (
            .O(N__10839),
            .I(N__10832));
    InMux I__2025 (
            .O(N__10838),
            .I(N__10829));
    InMux I__2024 (
            .O(N__10835),
            .I(N__10826));
    LocalMux I__2023 (
            .O(N__10832),
            .I(un8_beamy_3));
    LocalMux I__2022 (
            .O(N__10829),
            .I(un8_beamy_3));
    LocalMux I__2021 (
            .O(N__10826),
            .I(un8_beamy_3));
    CascadeMux I__2020 (
            .O(N__10819),
            .I(beamY_i_2_cascade_));
    CascadeMux I__2019 (
            .O(N__10816),
            .I(N__10811));
    InMux I__2018 (
            .O(N__10815),
            .I(N__10807));
    InMux I__2017 (
            .O(N__10814),
            .I(N__10802));
    InMux I__2016 (
            .O(N__10811),
            .I(N__10802));
    InMux I__2015 (
            .O(N__10810),
            .I(N__10799));
    LocalMux I__2014 (
            .O(N__10807),
            .I(beamY_i_2));
    LocalMux I__2013 (
            .O(N__10802),
            .I(beamY_i_2));
    LocalMux I__2012 (
            .O(N__10799),
            .I(beamY_i_2));
    InMux I__2011 (
            .O(N__10792),
            .I(N__10786));
    InMux I__2010 (
            .O(N__10791),
            .I(N__10786));
    LocalMux I__2009 (
            .O(N__10786),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0));
    InMux I__2008 (
            .O(N__10783),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__2007 (
            .O(N__10780),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__2006 (
            .O(N__10777),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__2005 (
            .O(N__10774),
            .I(N__10771));
    LocalMux I__2004 (
            .O(N__10771),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1));
    CascadeMux I__2003 (
            .O(N__10768),
            .I(g2_0_cascade_));
    CascadeMux I__2002 (
            .O(N__10765),
            .I(N__10762));
    InMux I__2001 (
            .O(N__10762),
            .I(N__10759));
    LocalMux I__2000 (
            .O(N__10759),
            .I(N__10756));
    Odrv4 I__1999 (
            .O(N__10756),
            .I(chary_if_generate_plus_mult1_un68_sum_1_5));
    IoInMux I__1998 (
            .O(N__10753),
            .I(N__10750));
    LocalMux I__1997 (
            .O(N__10750),
            .I(N__10747));
    Span4Mux_s3_v I__1996 (
            .O(N__10747),
            .I(N__10744));
    Odrv4 I__1995 (
            .O(N__10744),
            .I(VSync_c));
    CascadeMux I__1994 (
            .O(N__10741),
            .I(N__10738));
    InMux I__1993 (
            .O(N__10738),
            .I(N__10735));
    LocalMux I__1992 (
            .O(N__10735),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3));
    CascadeMux I__1991 (
            .O(N__10732),
            .I(N__10729));
    InMux I__1990 (
            .O(N__10729),
            .I(N__10726));
    LocalMux I__1989 (
            .O(N__10726),
            .I(un5_visibley_3_28));
    CascadeMux I__1988 (
            .O(N__10723),
            .I(un5_visibley_3_28_cascade_));
    CascadeMux I__1987 (
            .O(N__10720),
            .I(g1_3_cascade_));
    InMux I__1986 (
            .O(N__10717),
            .I(N__10714));
    LocalMux I__1985 (
            .O(N__10714),
            .I(g2_0_1));
    InMux I__1984 (
            .O(N__10711),
            .I(N__10708));
    LocalMux I__1983 (
            .O(N__10708),
            .I(N__10705));
    Odrv4 I__1982 (
            .O(N__10705),
            .I(un1_beamylto9_2));
    InMux I__1981 (
            .O(N__10702),
            .I(N__10696));
    InMux I__1980 (
            .O(N__10701),
            .I(N__10696));
    LocalMux I__1979 (
            .O(N__10696),
            .I(un5_visibley_1_28));
    CascadeMux I__1978 (
            .O(N__10693),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_));
    InMux I__1977 (
            .O(N__10690),
            .I(N__10687));
    LocalMux I__1976 (
            .O(N__10687),
            .I(chary_if_generate_plus_mult1_un68_sum_2_5));
    InMux I__1975 (
            .O(N__10684),
            .I(N__10681));
    LocalMux I__1974 (
            .O(N__10681),
            .I(un5_visibley_2_29));
    InMux I__1973 (
            .O(N__10678),
            .I(N__10675));
    LocalMux I__1972 (
            .O(N__10675),
            .I(g2_0_0));
    InMux I__1971 (
            .O(N__10672),
            .I(N__10669));
    LocalMux I__1970 (
            .O(N__10669),
            .I(beamY_RNIMSO1N7Z0Z_2));
    CascadeMux I__1969 (
            .O(N__10666),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_));
    InMux I__1968 (
            .O(N__10663),
            .I(N__10660));
    LocalMux I__1967 (
            .O(N__10660),
            .I(N__10657));
    Odrv12 I__1966 (
            .O(N__10657),
            .I(chary_if_generate_plus_mult1_un68_sum_1_0_5));
    InMux I__1965 (
            .O(N__10654),
            .I(N__10651));
    LocalMux I__1964 (
            .O(N__10651),
            .I(N__10648));
    Odrv4 I__1963 (
            .O(N__10648),
            .I(g2_0));
    CascadeMux I__1962 (
            .O(N__10645),
            .I(N__10642));
    InMux I__1961 (
            .O(N__10642),
            .I(N__10639));
    LocalMux I__1960 (
            .O(N__10639),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__1959 (
            .O(N__10636),
            .I(N__10633));
    LocalMux I__1958 (
            .O(N__10633),
            .I(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__1957 (
            .O(N__10630),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__1956 (
            .O(N__10627),
            .I(N__10624));
    LocalMux I__1955 (
            .O(N__10624),
            .I(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__1954 (
            .O(N__10621),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1953 (
            .O(N__10618),
            .I(content_column_1_i_2_2_cascade_));
    InMux I__1952 (
            .O(N__10615),
            .I(N__10611));
    InMux I__1951 (
            .O(N__10614),
            .I(N__10608));
    LocalMux I__1950 (
            .O(N__10611),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    LocalMux I__1949 (
            .O(N__10608),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    CascadeMux I__1948 (
            .O(N__10603),
            .I(N__10600));
    InMux I__1947 (
            .O(N__10600),
            .I(N__10597));
    LocalMux I__1946 (
            .O(N__10597),
            .I(if_generate_plus_mult1_un75_sum_axb_4_l_fx));
    InMux I__1945 (
            .O(N__10594),
            .I(N__10586));
    InMux I__1944 (
            .O(N__10593),
            .I(N__10586));
    InMux I__1943 (
            .O(N__10592),
            .I(N__10582));
    CascadeMux I__1942 (
            .O(N__10591),
            .I(N__10579));
    LocalMux I__1941 (
            .O(N__10586),
            .I(N__10576));
    InMux I__1940 (
            .O(N__10585),
            .I(N__10573));
    LocalMux I__1939 (
            .O(N__10582),
            .I(N__10570));
    InMux I__1938 (
            .O(N__10579),
            .I(N__10567));
    Span4Mux_h I__1937 (
            .O(N__10576),
            .I(N__10564));
    LocalMux I__1936 (
            .O(N__10573),
            .I(N__10561));
    Span4Mux_v I__1935 (
            .O(N__10570),
            .I(N__10556));
    LocalMux I__1934 (
            .O(N__10567),
            .I(N__10556));
    Odrv4 I__1933 (
            .O(N__10564),
            .I(chessboardpixel_un152_pixel_24));
    Odrv4 I__1932 (
            .O(N__10561),
            .I(chessboardpixel_un152_pixel_24));
    Odrv4 I__1931 (
            .O(N__10556),
            .I(chessboardpixel_un152_pixel_24));
    InMux I__1930 (
            .O(N__10549),
            .I(N__10546));
    LocalMux I__1929 (
            .O(N__10546),
            .I(column_1_if_generate_plus_mult1_un68_sum_iZ0));
    CascadeMux I__1928 (
            .O(N__10543),
            .I(content_m7_ns_1_cascade_));
    InMux I__1927 (
            .O(N__10540),
            .I(N__10533));
    InMux I__1926 (
            .O(N__10539),
            .I(N__10533));
    InMux I__1925 (
            .O(N__10538),
            .I(N__10530));
    LocalMux I__1924 (
            .O(N__10533),
            .I(N__10527));
    LocalMux I__1923 (
            .O(N__10530),
            .I(N__10524));
    Span4Mux_v I__1922 (
            .O(N__10527),
            .I(N__10521));
    Span4Mux_h I__1921 (
            .O(N__10524),
            .I(N__10518));
    Odrv4 I__1920 (
            .O(N__10521),
            .I(content_N_8));
    Odrv4 I__1919 (
            .O(N__10518),
            .I(content_N_8));
    CascadeMux I__1918 (
            .O(N__10513),
            .I(content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_));
    InMux I__1917 (
            .O(N__10510),
            .I(N__10507));
    LocalMux I__1916 (
            .O(N__10507),
            .I(N__10504));
    Odrv4 I__1915 (
            .O(N__10504),
            .I(content_content_ram7__RNI6B0NG3Z0Z_0));
    InMux I__1914 (
            .O(N__10501),
            .I(N__10498));
    LocalMux I__1913 (
            .O(N__10498),
            .I(content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0));
    CascadeMux I__1912 (
            .O(N__10495),
            .I(N__10492));
    InMux I__1911 (
            .O(N__10492),
            .I(N__10489));
    LocalMux I__1910 (
            .O(N__10489),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__1909 (
            .O(N__10486),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__1908 (
            .O(N__10483),
            .I(N__10480));
    LocalMux I__1907 (
            .O(N__10480),
            .I(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__1906 (
            .O(N__10477),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__1905 (
            .O(N__10474),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1904 (
            .O(N__10471),
            .I(N__10468));
    InMux I__1903 (
            .O(N__10468),
            .I(N__10465));
    LocalMux I__1902 (
            .O(N__10465),
            .I(content_column_1_i_2_i_2));
    InMux I__1901 (
            .O(N__10462),
            .I(N__10454));
    InMux I__1900 (
            .O(N__10461),
            .I(N__10454));
    InMux I__1899 (
            .O(N__10460),
            .I(N__10449));
    InMux I__1898 (
            .O(N__10459),
            .I(N__10449));
    LocalMux I__1897 (
            .O(N__10454),
            .I(N__10440));
    LocalMux I__1896 (
            .O(N__10449),
            .I(N__10440));
    InMux I__1895 (
            .O(N__10448),
            .I(N__10437));
    InMux I__1894 (
            .O(N__10447),
            .I(N__10432));
    InMux I__1893 (
            .O(N__10446),
            .I(N__10432));
    InMux I__1892 (
            .O(N__10445),
            .I(N__10429));
    Odrv4 I__1891 (
            .O(N__10440),
            .I(un6_rowlto1));
    LocalMux I__1890 (
            .O(N__10437),
            .I(un6_rowlto1));
    LocalMux I__1889 (
            .O(N__10432),
            .I(un6_rowlto1));
    LocalMux I__1888 (
            .O(N__10429),
            .I(un6_rowlto1));
    InMux I__1887 (
            .O(N__10420),
            .I(N__10414));
    InMux I__1886 (
            .O(N__10419),
            .I(N__10414));
    LocalMux I__1885 (
            .O(N__10414),
            .I(N__10411));
    Span4Mux_h I__1884 (
            .O(N__10411),
            .I(N__10408));
    Odrv4 I__1883 (
            .O(N__10408),
            .I(content_N_25));
    CascadeMux I__1882 (
            .O(N__10405),
            .I(N__10402));
    InMux I__1881 (
            .O(N__10402),
            .I(N__10399));
    LocalMux I__1880 (
            .O(N__10399),
            .I(column_1_if_generate_plus_mult1_un61_sum_iZ0));
    CascadeMux I__1879 (
            .O(N__10396),
            .I(N__10393));
    InMux I__1878 (
            .O(N__10393),
            .I(N__10390));
    LocalMux I__1877 (
            .O(N__10390),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    InMux I__1876 (
            .O(N__10387),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__1875 (
            .O(N__10384),
            .I(N__10381));
    InMux I__1874 (
            .O(N__10381),
            .I(N__10378));
    LocalMux I__1873 (
            .O(N__10378),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__1872 (
            .O(N__10375),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1871 (
            .O(N__10372),
            .I(N__10366));
    InMux I__1870 (
            .O(N__10371),
            .I(N__10366));
    LocalMux I__1869 (
            .O(N__10366),
            .I(column_1_if_generate_plus_mult1_un61_sum_i_5));
    IoInMux I__1868 (
            .O(N__10363),
            .I(N__10360));
    LocalMux I__1867 (
            .O(N__10360),
            .I(N__10357));
    IoSpan4Mux I__1866 (
            .O(N__10357),
            .I(N__10354));
    Sp12to4 I__1865 (
            .O(N__10354),
            .I(N__10351));
    Span12Mux_s7_v I__1864 (
            .O(N__10351),
            .I(N__10348));
    Odrv12 I__1863 (
            .O(N__10348),
            .I(GB_BUFFER_Clock12MHz_c_g_THRU_CO));
    CascadeMux I__1862 (
            .O(N__10345),
            .I(N__10338));
    InMux I__1861 (
            .O(N__10344),
            .I(N__10334));
    CascadeMux I__1860 (
            .O(N__10343),
            .I(N__10331));
    CascadeMux I__1859 (
            .O(N__10342),
            .I(N__10327));
    InMux I__1858 (
            .O(N__10341),
            .I(N__10323));
    InMux I__1857 (
            .O(N__10338),
            .I(N__10318));
    InMux I__1856 (
            .O(N__10337),
            .I(N__10318));
    LocalMux I__1855 (
            .O(N__10334),
            .I(N__10315));
    InMux I__1854 (
            .O(N__10331),
            .I(N__10308));
    InMux I__1853 (
            .O(N__10330),
            .I(N__10308));
    InMux I__1852 (
            .O(N__10327),
            .I(N__10308));
    InMux I__1851 (
            .O(N__10326),
            .I(N__10305));
    LocalMux I__1850 (
            .O(N__10323),
            .I(N__10300));
    LocalMux I__1849 (
            .O(N__10318),
            .I(N__10300));
    Span4Mux_v I__1848 (
            .O(N__10315),
            .I(N__10297));
    LocalMux I__1847 (
            .O(N__10308),
            .I(N__10292));
    LocalMux I__1846 (
            .O(N__10305),
            .I(N__10292));
    Span4Mux_v I__1845 (
            .O(N__10300),
            .I(N__10289));
    Span4Mux_h I__1844 (
            .O(N__10297),
            .I(N__10284));
    Span4Mux_v I__1843 (
            .O(N__10292),
            .I(N__10284));
    Odrv4 I__1842 (
            .O(N__10289),
            .I(charx_if_generate_plus_mult1_un75_sum));
    Odrv4 I__1841 (
            .O(N__10284),
            .I(charx_if_generate_plus_mult1_un75_sum));
    InMux I__1840 (
            .O(N__10279),
            .I(N__10273));
    InMux I__1839 (
            .O(N__10278),
            .I(N__10273));
    LocalMux I__1838 (
            .O(N__10273),
            .I(G_383));
    InMux I__1837 (
            .O(N__10270),
            .I(column_1_if_generate_plus_mult1_un82_sum_cry_4));
    InMux I__1836 (
            .O(N__10267),
            .I(N__10257));
    InMux I__1835 (
            .O(N__10266),
            .I(N__10257));
    InMux I__1834 (
            .O(N__10265),
            .I(N__10257));
    CascadeMux I__1833 (
            .O(N__10264),
            .I(N__10254));
    LocalMux I__1832 (
            .O(N__10257),
            .I(N__10250));
    InMux I__1831 (
            .O(N__10254),
            .I(N__10245));
    InMux I__1830 (
            .O(N__10253),
            .I(N__10245));
    Odrv4 I__1829 (
            .O(N__10250),
            .I(un6_rowlto0));
    LocalMux I__1828 (
            .O(N__10245),
            .I(un6_rowlto0));
    CascadeMux I__1827 (
            .O(N__10240),
            .I(N__10237));
    InMux I__1826 (
            .O(N__10237),
            .I(N__10234));
    LocalMux I__1825 (
            .O(N__10234),
            .I(column_1_if_generate_plus_mult1_un75_sum_iZ0));
    InMux I__1824 (
            .O(N__10231),
            .I(N__10227));
    InMux I__1823 (
            .O(N__10230),
            .I(N__10224));
    LocalMux I__1822 (
            .O(N__10227),
            .I(N__10218));
    LocalMux I__1821 (
            .O(N__10224),
            .I(N__10218));
    InMux I__1820 (
            .O(N__10223),
            .I(N__10215));
    Span4Mux_v I__1819 (
            .O(N__10218),
            .I(N__10209));
    LocalMux I__1818 (
            .O(N__10215),
            .I(N__10209));
    InMux I__1817 (
            .O(N__10214),
            .I(N__10206));
    Span4Mux_h I__1816 (
            .O(N__10209),
            .I(N__10201));
    LocalMux I__1815 (
            .O(N__10206),
            .I(N__10201));
    Odrv4 I__1814 (
            .O(N__10201),
            .I(charx_if_generate_plus_mult1_un68_sum));
    CascadeMux I__1813 (
            .O(N__10198),
            .I(N__10195));
    InMux I__1812 (
            .O(N__10195),
            .I(N__10192));
    LocalMux I__1811 (
            .O(N__10192),
            .I(if_generate_plus_mult1_un75_sum_cry_2_s));
    InMux I__1810 (
            .O(N__10189),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_1));
    CascadeMux I__1809 (
            .O(N__10186),
            .I(N__10182));
    InMux I__1808 (
            .O(N__10185),
            .I(N__10177));
    InMux I__1807 (
            .O(N__10182),
            .I(N__10177));
    LocalMux I__1806 (
            .O(N__10177),
            .I(un5_visibley_0_28));
    InMux I__1805 (
            .O(N__10174),
            .I(N__10171));
    LocalMux I__1804 (
            .O(N__10171),
            .I(g2));
    InMux I__1803 (
            .O(N__10168),
            .I(N__10165));
    LocalMux I__1802 (
            .O(N__10165),
            .I(N__10162));
    Odrv4 I__1801 (
            .O(N__10162),
            .I(un5_visibley_0_29));
    CascadeMux I__1800 (
            .O(N__10159),
            .I(N__10156));
    InMux I__1799 (
            .O(N__10156),
            .I(N__10153));
    LocalMux I__1798 (
            .O(N__10153),
            .I(N__10150));
    Odrv4 I__1797 (
            .O(N__10150),
            .I(Pixel_RNOZ0Z_67));
    CascadeMux I__1796 (
            .O(N__10147),
            .I(un4_beamylt6_cascade_));
    CascadeMux I__1795 (
            .O(N__10144),
            .I(N__10141));
    InMux I__1794 (
            .O(N__10141),
            .I(N__10138));
    LocalMux I__1793 (
            .O(N__10138),
            .I(N__10135));
    Odrv4 I__1792 (
            .O(N__10135),
            .I(un4_beamylt8_0));
    InMux I__1791 (
            .O(N__10132),
            .I(N__10129));
    LocalMux I__1790 (
            .O(N__10129),
            .I(chary_0_24));
    CascadeMux I__1789 (
            .O(N__10126),
            .I(N__10121));
    InMux I__1788 (
            .O(N__10125),
            .I(N__10112));
    InMux I__1787 (
            .O(N__10124),
            .I(N__10112));
    InMux I__1786 (
            .O(N__10121),
            .I(N__10107));
    InMux I__1785 (
            .O(N__10120),
            .I(N__10107));
    InMux I__1784 (
            .O(N__10119),
            .I(N__10100));
    InMux I__1783 (
            .O(N__10118),
            .I(N__10100));
    InMux I__1782 (
            .O(N__10117),
            .I(N__10100));
    LocalMux I__1781 (
            .O(N__10112),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_1));
    LocalMux I__1780 (
            .O(N__10107),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_1));
    LocalMux I__1779 (
            .O(N__10100),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_1));
    CascadeMux I__1778 (
            .O(N__10093),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_));
    InMux I__1777 (
            .O(N__10090),
            .I(N__10087));
    LocalMux I__1776 (
            .O(N__10087),
            .I(g1_2_0));
    CascadeMux I__1775 (
            .O(N__10084),
            .I(beamY_RNIMSO1N7_0Z0Z_2_cascade_));
    InMux I__1774 (
            .O(N__10081),
            .I(N__10075));
    InMux I__1773 (
            .O(N__10080),
            .I(N__10075));
    LocalMux I__1772 (
            .O(N__10075),
            .I(g4_0));
    InMux I__1771 (
            .O(N__10072),
            .I(N__10069));
    LocalMux I__1770 (
            .O(N__10069),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0));
    CascadeMux I__1769 (
            .O(N__10066),
            .I(g2_1_0_cascade_));
    InMux I__1768 (
            .O(N__10063),
            .I(N__10060));
    LocalMux I__1767 (
            .O(N__10060),
            .I(chary_if_generate_plus_mult1_un68_sum_0_5));
    InMux I__1766 (
            .O(N__10057),
            .I(N__10054));
    LocalMux I__1765 (
            .O(N__10054),
            .I(Pixel_RNOZ0Z_66));
    CascadeMux I__1764 (
            .O(N__10051),
            .I(N__10048));
    InMux I__1763 (
            .O(N__10048),
            .I(N__10045));
    LocalMux I__1762 (
            .O(N__10045),
            .I(N__10042));
    Odrv4 I__1761 (
            .O(N__10042),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    InMux I__1760 (
            .O(N__10039),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__1759 (
            .O(N__10036),
            .I(N__10033));
    InMux I__1758 (
            .O(N__10033),
            .I(N__10030));
    LocalMux I__1757 (
            .O(N__10030),
            .I(N__10027));
    Odrv4 I__1756 (
            .O(N__10027),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__1755 (
            .O(N__10024),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__1754 (
            .O(N__10021),
            .I(N__10018));
    LocalMux I__1753 (
            .O(N__10018),
            .I(N__10015));
    Odrv4 I__1752 (
            .O(N__10015),
            .I(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__1751 (
            .O(N__10012),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__1750 (
            .O(N__10009),
            .I(if_generate_plus_mult1_un61_sum_s_5_cascade_));
    InMux I__1749 (
            .O(N__10006),
            .I(N__9998));
    InMux I__1748 (
            .O(N__10005),
            .I(N__9998));
    InMux I__1747 (
            .O(N__10004),
            .I(N__9992));
    InMux I__1746 (
            .O(N__10003),
            .I(N__9989));
    LocalMux I__1745 (
            .O(N__9998),
            .I(N__9986));
    InMux I__1744 (
            .O(N__9997),
            .I(N__9983));
    InMux I__1743 (
            .O(N__9996),
            .I(N__9978));
    InMux I__1742 (
            .O(N__9995),
            .I(N__9978));
    LocalMux I__1741 (
            .O(N__9992),
            .I(N__9973));
    LocalMux I__1740 (
            .O(N__9989),
            .I(N__9973));
    Span4Mux_v I__1739 (
            .O(N__9986),
            .I(N__9970));
    LocalMux I__1738 (
            .O(N__9983),
            .I(N__9967));
    LocalMux I__1737 (
            .O(N__9978),
            .I(N__9964));
    Span4Mux_h I__1736 (
            .O(N__9973),
            .I(N__9961));
    Odrv4 I__1735 (
            .O(N__9970),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1734 (
            .O(N__9967),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1733 (
            .O(N__9964),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1732 (
            .O(N__9961),
            .I(charx_if_generate_plus_mult1_un54_sum));
    InMux I__1731 (
            .O(N__9952),
            .I(N__9946));
    InMux I__1730 (
            .O(N__9951),
            .I(N__9943));
    InMux I__1729 (
            .O(N__9950),
            .I(N__9940));
    InMux I__1728 (
            .O(N__9949),
            .I(N__9937));
    LocalMux I__1727 (
            .O(N__9946),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__1726 (
            .O(N__9943),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__1725 (
            .O(N__9940),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__1724 (
            .O(N__9937),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    InMux I__1723 (
            .O(N__9928),
            .I(N__9925));
    LocalMux I__1722 (
            .O(N__9925),
            .I(column_1_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__1721 (
            .O(N__9922),
            .I(N__9919));
    LocalMux I__1720 (
            .O(N__9919),
            .I(N__9916));
    Span4Mux_h I__1719 (
            .O(N__9916),
            .I(N__9913));
    Odrv4 I__1718 (
            .O(N__9913),
            .I(chary_2_24));
    CascadeMux I__1717 (
            .O(N__9910),
            .I(N__9906));
    InMux I__1716 (
            .O(N__9909),
            .I(N__9903));
    InMux I__1715 (
            .O(N__9906),
            .I(N__9898));
    LocalMux I__1714 (
            .O(N__9903),
            .I(N__9895));
    CascadeMux I__1713 (
            .O(N__9902),
            .I(N__9891));
    CascadeMux I__1712 (
            .O(N__9901),
            .I(N__9888));
    LocalMux I__1711 (
            .O(N__9898),
            .I(N__9884));
    Span12Mux_s5_h I__1710 (
            .O(N__9895),
            .I(N__9881));
    InMux I__1709 (
            .O(N__9894),
            .I(N__9878));
    InMux I__1708 (
            .O(N__9891),
            .I(N__9875));
    InMux I__1707 (
            .O(N__9888),
            .I(N__9870));
    InMux I__1706 (
            .O(N__9887),
            .I(N__9870));
    Span12Mux_s5_h I__1705 (
            .O(N__9884),
            .I(N__9867));
    Odrv12 I__1704 (
            .O(N__9881),
            .I(beamY_RNI539IG9Z0Z_3));
    LocalMux I__1703 (
            .O(N__9878),
            .I(beamY_RNI539IG9Z0Z_3));
    LocalMux I__1702 (
            .O(N__9875),
            .I(beamY_RNI539IG9Z0Z_3));
    LocalMux I__1701 (
            .O(N__9870),
            .I(beamY_RNI539IG9Z0Z_3));
    Odrv12 I__1700 (
            .O(N__9867),
            .I(beamY_RNI539IG9Z0Z_3));
    CascadeMux I__1699 (
            .O(N__9856),
            .I(beamY_RNI539IG9Z0Z_3_cascade_));
    InMux I__1698 (
            .O(N__9853),
            .I(N__9850));
    LocalMux I__1697 (
            .O(N__9850),
            .I(g4));
    InMux I__1696 (
            .O(N__9847),
            .I(N__9843));
    InMux I__1695 (
            .O(N__9846),
            .I(N__9836));
    LocalMux I__1694 (
            .O(N__9843),
            .I(N__9833));
    InMux I__1693 (
            .O(N__9842),
            .I(N__9830));
    InMux I__1692 (
            .O(N__9841),
            .I(N__9827));
    InMux I__1691 (
            .O(N__9840),
            .I(N__9824));
    InMux I__1690 (
            .O(N__9839),
            .I(N__9821));
    LocalMux I__1689 (
            .O(N__9836),
            .I(N__9818));
    Span4Mux_v I__1688 (
            .O(N__9833),
            .I(N__9813));
    LocalMux I__1687 (
            .O(N__9830),
            .I(N__9813));
    LocalMux I__1686 (
            .O(N__9827),
            .I(N__9808));
    LocalMux I__1685 (
            .O(N__9824),
            .I(N__9808));
    LocalMux I__1684 (
            .O(N__9821),
            .I(N__9805));
    Span4Mux_h I__1683 (
            .O(N__9818),
            .I(N__9802));
    Span4Mux_h I__1682 (
            .O(N__9813),
            .I(N__9799));
    Odrv12 I__1681 (
            .O(N__9808),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1680 (
            .O(N__9805),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1679 (
            .O(N__9802),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1678 (
            .O(N__9799),
            .I(charx_if_generate_plus_mult1_un47_sum));
    CascadeMux I__1677 (
            .O(N__9790),
            .I(N__9787));
    InMux I__1676 (
            .O(N__9787),
            .I(N__9784));
    LocalMux I__1675 (
            .O(N__9784),
            .I(N__9781));
    Odrv12 I__1674 (
            .O(N__9781),
            .I(charx_if_generate_plus_mult1_un40_sum_i));
    InMux I__1673 (
            .O(N__9778),
            .I(N__9775));
    LocalMux I__1672 (
            .O(N__9775),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1));
    InMux I__1671 (
            .O(N__9772),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1));
    InMux I__1670 (
            .O(N__9769),
            .I(N__9765));
    InMux I__1669 (
            .O(N__9768),
            .I(N__9762));
    LocalMux I__1668 (
            .O(N__9765),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    LocalMux I__1667 (
            .O(N__9762),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    CascadeMux I__1666 (
            .O(N__9757),
            .I(N__9754));
    InMux I__1665 (
            .O(N__9754),
            .I(N__9751));
    LocalMux I__1664 (
            .O(N__9751),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0));
    CascadeMux I__1663 (
            .O(N__9748),
            .I(N__9744));
    InMux I__1662 (
            .O(N__9747),
            .I(N__9739));
    InMux I__1661 (
            .O(N__9744),
            .I(N__9739));
    LocalMux I__1660 (
            .O(N__9739),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2));
    InMux I__1659 (
            .O(N__9736),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__1658 (
            .O(N__9733),
            .I(N__9727));
    InMux I__1657 (
            .O(N__9732),
            .I(N__9727));
    LocalMux I__1656 (
            .O(N__9727),
            .I(charx_if_generate_plus_mult1_un40_sum_i_5));
    CascadeMux I__1655 (
            .O(N__9724),
            .I(N__9721));
    InMux I__1654 (
            .O(N__9721),
            .I(N__9718));
    LocalMux I__1653 (
            .O(N__9718),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1));
    InMux I__1652 (
            .O(N__9715),
            .I(N__9712));
    LocalMux I__1651 (
            .O(N__9712),
            .I(charx_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__1650 (
            .O(N__9709),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__1649 (
            .O(N__9706),
            .I(N__9703));
    LocalMux I__1648 (
            .O(N__9703),
            .I(charx_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__1647 (
            .O(N__9700),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__1646 (
            .O(N__9697),
            .I(N__9693));
    InMux I__1645 (
            .O(N__9696),
            .I(N__9689));
    InMux I__1644 (
            .O(N__9693),
            .I(N__9684));
    InMux I__1643 (
            .O(N__9692),
            .I(N__9684));
    LocalMux I__1642 (
            .O(N__9689),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    LocalMux I__1641 (
            .O(N__9684),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    CascadeMux I__1640 (
            .O(N__9679),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_));
    InMux I__1639 (
            .O(N__9676),
            .I(N__9673));
    LocalMux I__1638 (
            .O(N__9673),
            .I(charx_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__1637 (
            .O(N__9670),
            .I(N__9667));
    LocalMux I__1636 (
            .O(N__9667),
            .I(un5_visiblex_i_27));
    CascadeMux I__1635 (
            .O(N__9664),
            .I(N__9661));
    InMux I__1634 (
            .O(N__9661),
            .I(N__9658));
    LocalMux I__1633 (
            .O(N__9658),
            .I(N__9654));
    InMux I__1632 (
            .O(N__9657),
            .I(N__9651));
    Odrv4 I__1631 (
            .O(N__9654),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO));
    LocalMux I__1630 (
            .O(N__9651),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO));
    InMux I__1629 (
            .O(N__9646),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__1628 (
            .O(N__9643),
            .I(N__9640));
    LocalMux I__1627 (
            .O(N__9640),
            .I(content_content_ram0__RNIR1C2R81_0Z0Z_0));
    InMux I__1626 (
            .O(N__9637),
            .I(N__9634));
    LocalMux I__1625 (
            .O(N__9634),
            .I(un6_rowlt7_0));
    CascadeMux I__1624 (
            .O(N__9631),
            .I(N__9628));
    InMux I__1623 (
            .O(N__9628),
            .I(N__9625));
    LocalMux I__1622 (
            .O(N__9625),
            .I(N__9622));
    Odrv12 I__1621 (
            .O(N__9622),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3));
    InMux I__1620 (
            .O(N__9619),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1));
    CascadeMux I__1619 (
            .O(N__9616),
            .I(N__9613));
    InMux I__1618 (
            .O(N__9613),
            .I(N__9610));
    LocalMux I__1617 (
            .O(N__9610),
            .I(N__9607));
    Odrv4 I__1616 (
            .O(N__9607),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5));
    InMux I__1615 (
            .O(N__9604),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__1614 (
            .O(N__9601),
            .I(N__9598));
    LocalMux I__1613 (
            .O(N__9598),
            .I(N__9595));
    Odrv4 I__1612 (
            .O(N__9595),
            .I(charx_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__1611 (
            .O(N__9592),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__1610 (
            .O(N__9589),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__1609 (
            .O(N__9586),
            .I(N__9583));
    LocalMux I__1608 (
            .O(N__9583),
            .I(N__9578));
    InMux I__1607 (
            .O(N__9582),
            .I(N__9575));
    InMux I__1606 (
            .O(N__9581),
            .I(N__9572));
    Odrv4 I__1605 (
            .O(N__9578),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7));
    LocalMux I__1604 (
            .O(N__9575),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7));
    LocalMux I__1603 (
            .O(N__9572),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7));
    CascadeMux I__1602 (
            .O(N__9565),
            .I(N__9562));
    InMux I__1601 (
            .O(N__9562),
            .I(N__9559));
    LocalMux I__1600 (
            .O(N__9559),
            .I(charx_if_generate_plus_mult1_un47_sum_i));
    InMux I__1599 (
            .O(N__9556),
            .I(N__9553));
    LocalMux I__1598 (
            .O(N__9553),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6));
    InMux I__1597 (
            .O(N__9550),
            .I(N__9547));
    LocalMux I__1596 (
            .O(N__9547),
            .I(g4_1));
    InMux I__1595 (
            .O(N__9544),
            .I(N__9541));
    LocalMux I__1594 (
            .O(N__9541),
            .I(N__9538));
    Span4Mux_h I__1593 (
            .O(N__9538),
            .I(N__9535));
    Odrv4 I__1592 (
            .O(N__9535),
            .I(g0_0_a3_5));
    CascadeMux I__1591 (
            .O(N__9532),
            .I(m4_rn_1_cascade_));
    InMux I__1590 (
            .O(N__9529),
            .I(N__9526));
    LocalMux I__1589 (
            .O(N__9526),
            .I(N__9523));
    Span4Mux_h I__1588 (
            .O(N__9523),
            .I(N__9520));
    Odrv4 I__1587 (
            .O(N__9520),
            .I(Pixel_RNOZ0Z_40));
    CascadeMux I__1586 (
            .O(N__9517),
            .I(content_content_ram0__RNIR1C2R81Z0Z_0_cascade_));
    InMux I__1585 (
            .O(N__9514),
            .I(N__9505));
    InMux I__1584 (
            .O(N__9513),
            .I(N__9499));
    InMux I__1583 (
            .O(N__9512),
            .I(N__9496));
    InMux I__1582 (
            .O(N__9511),
            .I(N__9493));
    InMux I__1581 (
            .O(N__9510),
            .I(N__9488));
    InMux I__1580 (
            .O(N__9509),
            .I(N__9483));
    InMux I__1579 (
            .O(N__9508),
            .I(N__9483));
    LocalMux I__1578 (
            .O(N__9505),
            .I(N__9480));
    InMux I__1577 (
            .O(N__9504),
            .I(N__9473));
    InMux I__1576 (
            .O(N__9503),
            .I(N__9473));
    InMux I__1575 (
            .O(N__9502),
            .I(N__9473));
    LocalMux I__1574 (
            .O(N__9499),
            .I(N__9468));
    LocalMux I__1573 (
            .O(N__9496),
            .I(N__9468));
    LocalMux I__1572 (
            .O(N__9493),
            .I(N__9464));
    InMux I__1571 (
            .O(N__9492),
            .I(N__9459));
    InMux I__1570 (
            .O(N__9491),
            .I(N__9459));
    LocalMux I__1569 (
            .O(N__9488),
            .I(N__9455));
    LocalMux I__1568 (
            .O(N__9483),
            .I(N__9446));
    Span4Mux_h I__1567 (
            .O(N__9480),
            .I(N__9446));
    LocalMux I__1566 (
            .O(N__9473),
            .I(N__9446));
    Span4Mux_h I__1565 (
            .O(N__9468),
            .I(N__9446));
    InMux I__1564 (
            .O(N__9467),
            .I(N__9443));
    Span4Mux_s3_v I__1563 (
            .O(N__9464),
            .I(N__9438));
    LocalMux I__1562 (
            .O(N__9459),
            .I(N__9438));
    InMux I__1561 (
            .O(N__9458),
            .I(N__9435));
    Odrv12 I__1560 (
            .O(N__9455),
            .I(N_331_i));
    Odrv4 I__1559 (
            .O(N__9446),
            .I(N_331_i));
    LocalMux I__1558 (
            .O(N__9443),
            .I(N_331_i));
    Odrv4 I__1557 (
            .O(N__9438),
            .I(N_331_i));
    LocalMux I__1556 (
            .O(N__9435),
            .I(N_331_i));
    CascadeMux I__1555 (
            .O(N__9424),
            .I(un4_row_m7_ns_1_cascade_));
    CascadeMux I__1554 (
            .O(N__9421),
            .I(N__9418));
    InMux I__1553 (
            .O(N__9418),
            .I(N__9415));
    LocalMux I__1552 (
            .O(N__9415),
            .I(beamY_RNIPAQ91Z0Z_6));
    InMux I__1551 (
            .O(N__9412),
            .I(N__9409));
    LocalMux I__1550 (
            .O(N__9409),
            .I(un4_beamy_0));
    InMux I__1549 (
            .O(N__9406),
            .I(N__9403));
    LocalMux I__1548 (
            .O(N__9403),
            .I(m4_sn));
    CascadeMux I__1547 (
            .O(N__9400),
            .I(chary_1_24_cascade_));
    InMux I__1546 (
            .O(N__9397),
            .I(N__9394));
    LocalMux I__1545 (
            .O(N__9394),
            .I(N_1737_0));
    CascadeMux I__1544 (
            .O(N__9391),
            .I(chary_1_0_24_cascade_));
    CascadeMux I__1543 (
            .O(N__9388),
            .I(g2_3_cascade_));
    InMux I__1542 (
            .O(N__9385),
            .I(N__9382));
    LocalMux I__1541 (
            .O(N__9382),
            .I(g1_1_1));
    InMux I__1540 (
            .O(N__9379),
            .I(N__9376));
    LocalMux I__1539 (
            .O(N__9376),
            .I(un116_pixel_0_0_0));
    InMux I__1538 (
            .O(N__9373),
            .I(N__9370));
    LocalMux I__1537 (
            .O(N__9370),
            .I(N_5_1));
    InMux I__1536 (
            .O(N__9367),
            .I(N__9364));
    LocalMux I__1535 (
            .O(N__9364),
            .I(N__9361));
    Span4Mux_h I__1534 (
            .O(N__9361),
            .I(N__9358));
    Odrv4 I__1533 (
            .O(N__9358),
            .I(g0_0_a3_4));
    CascadeMux I__1532 (
            .O(N__9355),
            .I(un8_beamylto9_1_cascade_));
    InMux I__1531 (
            .O(N__9352),
            .I(N__9349));
    LocalMux I__1530 (
            .O(N__9349),
            .I(un8_beamy));
    InMux I__1529 (
            .O(N__9346),
            .I(N__9343));
    LocalMux I__1528 (
            .O(N__9343),
            .I(N_134_0));
    CascadeMux I__1527 (
            .O(N__9340),
            .I(font_un28_pixel_29_cascade_));
    InMux I__1526 (
            .O(N__9337),
            .I(N__9334));
    LocalMux I__1525 (
            .O(N__9334),
            .I(N__9331));
    Odrv4 I__1524 (
            .O(N__9331),
            .I(beamY_RNIDA2GGA3Z0Z_0));
    InMux I__1523 (
            .O(N__9328),
            .I(N__9325));
    LocalMux I__1522 (
            .O(N__9325),
            .I(N__9322));
    Odrv12 I__1521 (
            .O(N__9322),
            .I(g0_1));
    InMux I__1520 (
            .O(N__9319),
            .I(N__9312));
    InMux I__1519 (
            .O(N__9318),
            .I(N__9309));
    InMux I__1518 (
            .O(N__9317),
            .I(N__9300));
    InMux I__1517 (
            .O(N__9316),
            .I(N__9300));
    CascadeMux I__1516 (
            .O(N__9315),
            .I(N__9297));
    LocalMux I__1515 (
            .O(N__9312),
            .I(N__9291));
    LocalMux I__1514 (
            .O(N__9309),
            .I(N__9288));
    InMux I__1513 (
            .O(N__9308),
            .I(N__9285));
    InMux I__1512 (
            .O(N__9307),
            .I(N__9278));
    InMux I__1511 (
            .O(N__9306),
            .I(N__9278));
    InMux I__1510 (
            .O(N__9305),
            .I(N__9278));
    LocalMux I__1509 (
            .O(N__9300),
            .I(N__9275));
    InMux I__1508 (
            .O(N__9297),
            .I(N__9270));
    InMux I__1507 (
            .O(N__9296),
            .I(N__9270));
    InMux I__1506 (
            .O(N__9295),
            .I(N__9265));
    InMux I__1505 (
            .O(N__9294),
            .I(N__9265));
    Span4Mux_h I__1504 (
            .O(N__9291),
            .I(N__9262));
    Odrv12 I__1503 (
            .O(N__9288),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__1502 (
            .O(N__9285),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__1501 (
            .O(N__9278),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    Odrv4 I__1500 (
            .O(N__9275),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__1499 (
            .O(N__9270),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__1498 (
            .O(N__9265),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    Odrv4 I__1497 (
            .O(N__9262),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    CascadeMux I__1496 (
            .O(N__9247),
            .I(beamY_RNIDA2GGA3Z0Z_0_cascade_));
    InMux I__1495 (
            .O(N__9244),
            .I(N__9241));
    LocalMux I__1494 (
            .O(N__9241),
            .I(N_19_0_0));
    InMux I__1493 (
            .O(N__9238),
            .I(N__9235));
    LocalMux I__1492 (
            .O(N__9235),
            .I(font_un28_pixel_30));
    InMux I__1491 (
            .O(N__9232),
            .I(N__9228));
    InMux I__1490 (
            .O(N__9231),
            .I(N__9225));
    LocalMux I__1489 (
            .O(N__9228),
            .I(N__9222));
    LocalMux I__1488 (
            .O(N__9225),
            .I(font_un28_pixel_29));
    Odrv4 I__1487 (
            .O(N__9222),
            .I(font_un28_pixel_29));
    InMux I__1486 (
            .O(N__9217),
            .I(N__9214));
    LocalMux I__1485 (
            .O(N__9214),
            .I(N_15_i));
    CascadeMux I__1484 (
            .O(N__9211),
            .I(Pixel_RNOZ0Z_28_cascade_));
    InMux I__1483 (
            .O(N__9208),
            .I(N__9205));
    LocalMux I__1482 (
            .O(N__9205),
            .I(N__9202));
    Odrv4 I__1481 (
            .O(N__9202),
            .I(Pixel_RNOZ0Z_9));
    InMux I__1480 (
            .O(N__9199),
            .I(N__9193));
    InMux I__1479 (
            .O(N__9198),
            .I(N__9193));
    LocalMux I__1478 (
            .O(N__9193),
            .I(N__9189));
    InMux I__1477 (
            .O(N__9192),
            .I(N__9185));
    Span4Mux_v I__1476 (
            .O(N__9189),
            .I(N__9182));
    InMux I__1475 (
            .O(N__9188),
            .I(N__9179));
    LocalMux I__1474 (
            .O(N__9185),
            .I(chary_24));
    Odrv4 I__1473 (
            .O(N__9182),
            .I(chary_24));
    LocalMux I__1472 (
            .O(N__9179),
            .I(chary_24));
    InMux I__1471 (
            .O(N__9172),
            .I(N__9169));
    LocalMux I__1470 (
            .O(N__9169),
            .I(N__9165));
    InMux I__1469 (
            .O(N__9168),
            .I(N__9161));
    Span4Mux_h I__1468 (
            .O(N__9165),
            .I(N__9158));
    InMux I__1467 (
            .O(N__9164),
            .I(N__9155));
    LocalMux I__1466 (
            .O(N__9161),
            .I(N__9152));
    Odrv4 I__1465 (
            .O(N__9158),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    LocalMux I__1464 (
            .O(N__9155),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    Odrv4 I__1463 (
            .O(N__9152),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    InMux I__1462 (
            .O(N__9145),
            .I(N__9139));
    InMux I__1461 (
            .O(N__9144),
            .I(N__9139));
    LocalMux I__1460 (
            .O(N__9139),
            .I(charx_if_generate_plus_mult1_un33_sum_i_5));
    InMux I__1459 (
            .O(N__9136),
            .I(N__9127));
    InMux I__1458 (
            .O(N__9135),
            .I(N__9127));
    CascadeMux I__1457 (
            .O(N__9134),
            .I(N__9123));
    CascadeMux I__1456 (
            .O(N__9133),
            .I(N__9120));
    InMux I__1455 (
            .O(N__9132),
            .I(N__9116));
    LocalMux I__1454 (
            .O(N__9127),
            .I(N__9113));
    InMux I__1453 (
            .O(N__9126),
            .I(N__9110));
    InMux I__1452 (
            .O(N__9123),
            .I(N__9105));
    InMux I__1451 (
            .O(N__9120),
            .I(N__9105));
    CascadeMux I__1450 (
            .O(N__9119),
            .I(N__9101));
    LocalMux I__1449 (
            .O(N__9116),
            .I(N__9095));
    Span4Mux_h I__1448 (
            .O(N__9113),
            .I(N__9092));
    LocalMux I__1447 (
            .O(N__9110),
            .I(N__9087));
    LocalMux I__1446 (
            .O(N__9105),
            .I(N__9087));
    InMux I__1445 (
            .O(N__9104),
            .I(N__9084));
    InMux I__1444 (
            .O(N__9101),
            .I(N__9081));
    InMux I__1443 (
            .O(N__9100),
            .I(N__9074));
    InMux I__1442 (
            .O(N__9099),
            .I(N__9074));
    InMux I__1441 (
            .O(N__9098),
            .I(N__9074));
    Odrv4 I__1440 (
            .O(N__9095),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    Odrv4 I__1439 (
            .O(N__9092),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    Odrv4 I__1438 (
            .O(N__9087),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    LocalMux I__1437 (
            .O(N__9084),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    LocalMux I__1436 (
            .O(N__9081),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    LocalMux I__1435 (
            .O(N__9074),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3));
    CascadeMux I__1434 (
            .O(N__9061),
            .I(N__9058));
    InMux I__1433 (
            .O(N__9058),
            .I(N__9055));
    LocalMux I__1432 (
            .O(N__9055),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i));
    InMux I__1431 (
            .O(N__9052),
            .I(N__9049));
    LocalMux I__1430 (
            .O(N__9049),
            .I(N__9046));
    Odrv4 I__1429 (
            .O(N__9046),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO));
    InMux I__1428 (
            .O(N__9043),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6));
    InMux I__1427 (
            .O(N__9040),
            .I(N__9033));
    InMux I__1426 (
            .O(N__9039),
            .I(N__9033));
    InMux I__1425 (
            .O(N__9038),
            .I(N__9030));
    LocalMux I__1424 (
            .O(N__9033),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0));
    LocalMux I__1423 (
            .O(N__9030),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0));
    InMux I__1422 (
            .O(N__9025),
            .I(N__9019));
    InMux I__1421 (
            .O(N__9024),
            .I(N__9019));
    LocalMux I__1420 (
            .O(N__9019),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8));
    InMux I__1419 (
            .O(N__9016),
            .I(N__9013));
    LocalMux I__1418 (
            .O(N__9013),
            .I(N__9010));
    Odrv12 I__1417 (
            .O(N__9010),
            .I(Pixel_RNOZ0Z_14));
    InMux I__1416 (
            .O(N__9007),
            .I(N__9004));
    LocalMux I__1415 (
            .O(N__9004),
            .I(N__9001));
    Odrv12 I__1414 (
            .O(N__9001),
            .I(font_un126_pixel_5_a0_1));
    InMux I__1413 (
            .O(N__8998),
            .I(N__8995));
    LocalMux I__1412 (
            .O(N__8995),
            .I(N__8992));
    Span12Mux_s3_v I__1411 (
            .O(N__8992),
            .I(N__8989));
    Odrv12 I__1410 (
            .O(N__8989),
            .I(N_1740_0));
    CascadeMux I__1409 (
            .O(N__8986),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_));
    InMux I__1408 (
            .O(N__8983),
            .I(N__8980));
    LocalMux I__1407 (
            .O(N__8980),
            .I(N__8974));
    InMux I__1406 (
            .O(N__8979),
            .I(N__8969));
    InMux I__1405 (
            .O(N__8978),
            .I(N__8969));
    InMux I__1404 (
            .O(N__8977),
            .I(N__8964));
    Span4Mux_v I__1403 (
            .O(N__8974),
            .I(N__8956));
    LocalMux I__1402 (
            .O(N__8969),
            .I(N__8956));
    InMux I__1401 (
            .O(N__8968),
            .I(N__8953));
    CascadeMux I__1400 (
            .O(N__8967),
            .I(N__8950));
    LocalMux I__1399 (
            .O(N__8964),
            .I(N__8947));
    InMux I__1398 (
            .O(N__8963),
            .I(N__8940));
    InMux I__1397 (
            .O(N__8962),
            .I(N__8940));
    InMux I__1396 (
            .O(N__8961),
            .I(N__8940));
    Span4Mux_h I__1395 (
            .O(N__8956),
            .I(N__8937));
    LocalMux I__1394 (
            .O(N__8953),
            .I(N__8934));
    InMux I__1393 (
            .O(N__8950),
            .I(N__8931));
    Odrv12 I__1392 (
            .O(N__8947),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__1391 (
            .O(N__8940),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv4 I__1390 (
            .O(N__8937),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv12 I__1389 (
            .O(N__8934),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__1388 (
            .O(N__8931),
            .I(charx_if_generate_plus_mult1_un33_sum));
    CascadeMux I__1387 (
            .O(N__8920),
            .I(N__8917));
    InMux I__1386 (
            .O(N__8917),
            .I(N__8914));
    LocalMux I__1385 (
            .O(N__8914),
            .I(charx_if_generate_plus_mult1_un33_sum_i));
    CascadeMux I__1384 (
            .O(N__8911),
            .I(N__8908));
    InMux I__1383 (
            .O(N__8908),
            .I(N__8895));
    InMux I__1382 (
            .O(N__8907),
            .I(N__8895));
    InMux I__1381 (
            .O(N__8906),
            .I(N__8895));
    InMux I__1380 (
            .O(N__8905),
            .I(N__8888));
    InMux I__1379 (
            .O(N__8904),
            .I(N__8888));
    InMux I__1378 (
            .O(N__8903),
            .I(N__8888));
    InMux I__1377 (
            .O(N__8902),
            .I(N__8885));
    LocalMux I__1376 (
            .O(N__8895),
            .I(N__8880));
    LocalMux I__1375 (
            .O(N__8888),
            .I(N__8880));
    LocalMux I__1374 (
            .O(N__8885),
            .I(N__8875));
    Span4Mux_h I__1373 (
            .O(N__8880),
            .I(N__8872));
    InMux I__1372 (
            .O(N__8879),
            .I(N__8869));
    InMux I__1371 (
            .O(N__8878),
            .I(N__8866));
    Odrv4 I__1370 (
            .O(N__8875),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1369 (
            .O(N__8872),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1368 (
            .O(N__8869),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1367 (
            .O(N__8866),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    CascadeMux I__1366 (
            .O(N__8857),
            .I(N__8854));
    InMux I__1365 (
            .O(N__8854),
            .I(N__8851));
    LocalMux I__1364 (
            .O(N__8851),
            .I(N__8848));
    Odrv12 I__1363 (
            .O(N__8848),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421));
    InMux I__1362 (
            .O(N__8845),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__1361 (
            .O(N__8842),
            .I(N__8839));
    InMux I__1360 (
            .O(N__8839),
            .I(N__8836));
    LocalMux I__1359 (
            .O(N__8836),
            .I(N__8833));
    Span4Mux_v I__1358 (
            .O(N__8833),
            .I(N__8830));
    Odrv4 I__1357 (
            .O(N__8830),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0));
    CascadeMux I__1356 (
            .O(N__8827),
            .I(N__8824));
    InMux I__1355 (
            .O(N__8824),
            .I(N__8821));
    LocalMux I__1354 (
            .O(N__8821),
            .I(N__8818));
    Odrv12 I__1353 (
            .O(N__8818),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1));
    InMux I__1352 (
            .O(N__8815),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    CascadeMux I__1351 (
            .O(N__8812),
            .I(N__8809));
    InMux I__1350 (
            .O(N__8809),
            .I(N__8806));
    LocalMux I__1349 (
            .O(N__8806),
            .I(N__8803));
    Span4Mux_h I__1348 (
            .O(N__8803),
            .I(N__8800));
    Odrv4 I__1347 (
            .O(N__8800),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0));
    InMux I__1346 (
            .O(N__8797),
            .I(N__8794));
    LocalMux I__1345 (
            .O(N__8794),
            .I(N__8791));
    Odrv12 I__1344 (
            .O(N__8791),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__1343 (
            .O(N__8788),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__1342 (
            .O(N__8785),
            .I(N__8782));
    LocalMux I__1341 (
            .O(N__8782),
            .I(N__8779));
    Span4Mux_h I__1340 (
            .O(N__8779),
            .I(N__8776));
    Odrv4 I__1339 (
            .O(N__8776),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__1338 (
            .O(N__8773),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__1337 (
            .O(N__8770),
            .I(N__8767));
    LocalMux I__1336 (
            .O(N__8767),
            .I(N__8762));
    InMux I__1335 (
            .O(N__8766),
            .I(N__8759));
    InMux I__1334 (
            .O(N__8765),
            .I(N__8756));
    Span4Mux_h I__1333 (
            .O(N__8762),
            .I(N__8751));
    LocalMux I__1332 (
            .O(N__8759),
            .I(N__8751));
    LocalMux I__1331 (
            .O(N__8756),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1));
    Odrv4 I__1330 (
            .O(N__8751),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1));
    InMux I__1329 (
            .O(N__8746),
            .I(N__8743));
    LocalMux I__1328 (
            .O(N__8743),
            .I(un4_row_9_0));
    CascadeMux I__1327 (
            .O(N__8740),
            .I(N__8737));
    InMux I__1326 (
            .O(N__8737),
            .I(N__8734));
    LocalMux I__1325 (
            .O(N__8734),
            .I(N__8731));
    Odrv4 I__1324 (
            .O(N__8731),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__1323 (
            .O(N__8728),
            .I(N__8723));
    InMux I__1322 (
            .O(N__8727),
            .I(N__8718));
    InMux I__1321 (
            .O(N__8726),
            .I(N__8718));
    LocalMux I__1320 (
            .O(N__8723),
            .I(column_1_if_generate_plus_mult1_un47_sum_cZ0Z5));
    LocalMux I__1319 (
            .O(N__8718),
            .I(column_1_if_generate_plus_mult1_un47_sum_cZ0Z5));
    CascadeMux I__1318 (
            .O(N__8713),
            .I(N__8710));
    InMux I__1317 (
            .O(N__8710),
            .I(N__8707));
    LocalMux I__1316 (
            .O(N__8707),
            .I(N__8701));
    InMux I__1315 (
            .O(N__8706),
            .I(N__8698));
    InMux I__1314 (
            .O(N__8705),
            .I(N__8692));
    InMux I__1313 (
            .O(N__8704),
            .I(N__8692));
    Span4Mux_v I__1312 (
            .O(N__8701),
            .I(N__8686));
    LocalMux I__1311 (
            .O(N__8698),
            .I(N__8686));
    InMux I__1310 (
            .O(N__8697),
            .I(N__8680));
    LocalMux I__1309 (
            .O(N__8692),
            .I(N__8677));
    InMux I__1308 (
            .O(N__8691),
            .I(N__8674));
    Span4Mux_h I__1307 (
            .O(N__8686),
            .I(N__8671));
    InMux I__1306 (
            .O(N__8685),
            .I(N__8664));
    InMux I__1305 (
            .O(N__8684),
            .I(N__8664));
    InMux I__1304 (
            .O(N__8683),
            .I(N__8664));
    LocalMux I__1303 (
            .O(N__8680),
            .I(N__8661));
    Odrv12 I__1302 (
            .O(N__8677),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__1301 (
            .O(N__8674),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__1300 (
            .O(N__8671),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__1299 (
            .O(N__8664),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv12 I__1298 (
            .O(N__8661),
            .I(charx_if_generate_plus_mult1_un40_sum));
    InMux I__1297 (
            .O(N__8650),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1));
    CascadeMux I__1296 (
            .O(N__8647),
            .I(N__8644));
    InMux I__1295 (
            .O(N__8644),
            .I(N__8641));
    LocalMux I__1294 (
            .O(N__8641),
            .I(N__8638));
    Span4Mux_v I__1293 (
            .O(N__8638),
            .I(N__8635));
    Odrv4 I__1292 (
            .O(N__8635),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0));
    InMux I__1291 (
            .O(N__8632),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__1290 (
            .O(N__8629),
            .I(N__8626));
    InMux I__1289 (
            .O(N__8626),
            .I(N__8623));
    LocalMux I__1288 (
            .O(N__8623),
            .I(N__8620));
    Span4Mux_h I__1287 (
            .O(N__8620),
            .I(N__8617));
    Odrv4 I__1286 (
            .O(N__8617),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0));
    InMux I__1285 (
            .O(N__8614),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__1284 (
            .O(N__8611),
            .I(N__8608));
    LocalMux I__1283 (
            .O(N__8608),
            .I(N__8605));
    Span4Mux_h I__1282 (
            .O(N__8605),
            .I(N__8602));
    Odrv4 I__1281 (
            .O(N__8602),
            .I(charx_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__1280 (
            .O(N__8599),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__1279 (
            .O(N__8596),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__1278 (
            .O(N__8593),
            .I(N__8590));
    LocalMux I__1277 (
            .O(N__8590),
            .I(N__8587));
    Span4Mux_v I__1276 (
            .O(N__8587),
            .I(N__8584));
    Odrv4 I__1275 (
            .O(N__8584),
            .I(if_generate_plus_mult1_un54_sum_axb_3_l_ofx));
    CascadeMux I__1274 (
            .O(N__8581),
            .I(N__8578));
    InMux I__1273 (
            .O(N__8578),
            .I(N__8575));
    LocalMux I__1272 (
            .O(N__8575),
            .I(N__8572));
    Span4Mux_h I__1271 (
            .O(N__8572),
            .I(N__8569));
    Odrv4 I__1270 (
            .O(N__8569),
            .I(column_1_if_generate_plus_mult1_un47_sum_c5_iZ0));
    InMux I__1269 (
            .O(N__8566),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__1268 (
            .O(N__8563),
            .I(N__8560));
    InMux I__1267 (
            .O(N__8560),
            .I(N__8557));
    LocalMux I__1266 (
            .O(N__8557),
            .I(N__8554));
    Span4Mux_h I__1265 (
            .O(N__8554),
            .I(N__8551));
    Odrv4 I__1264 (
            .O(N__8551),
            .I(if_generate_plus_mult1_un54_sum_axb_4_l_ofx));
    InMux I__1263 (
            .O(N__8548),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__1262 (
            .O(N__8545),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__1261 (
            .O(N__8542),
            .I(N__8536));
    InMux I__1260 (
            .O(N__8541),
            .I(N__8536));
    LocalMux I__1259 (
            .O(N__8536),
            .I(N__8533));
    Odrv4 I__1258 (
            .O(N__8533),
            .I(charx_if_generate_plus_mult1_un54_sum_i_5));
    CascadeMux I__1257 (
            .O(N__8530),
            .I(N__8527));
    InMux I__1256 (
            .O(N__8527),
            .I(N__8524));
    LocalMux I__1255 (
            .O(N__8524),
            .I(un5_visiblex_i_26));
    InMux I__1254 (
            .O(N__8521),
            .I(N__8515));
    InMux I__1253 (
            .O(N__8520),
            .I(N__8515));
    LocalMux I__1252 (
            .O(N__8515),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__1251 (
            .O(N__8512),
            .I(un4_row_9_2_cascade_));
    InMux I__1250 (
            .O(N__8509),
            .I(N__8506));
    LocalMux I__1249 (
            .O(N__8506),
            .I(N__8503));
    Odrv4 I__1248 (
            .O(N__8503),
            .I(un4_row_9_5));
    CascadeMux I__1247 (
            .O(N__8500),
            .I(N__8496));
    InMux I__1246 (
            .O(N__8499),
            .I(N__8491));
    InMux I__1245 (
            .O(N__8496),
            .I(N__8491));
    LocalMux I__1244 (
            .O(N__8491),
            .I(N__8488));
    Span4Mux_v I__1243 (
            .O(N__8488),
            .I(N__8483));
    InMux I__1242 (
            .O(N__8487),
            .I(N__8478));
    InMux I__1241 (
            .O(N__8486),
            .I(N__8478));
    Span4Mux_v I__1240 (
            .O(N__8483),
            .I(N__8475));
    LocalMux I__1239 (
            .O(N__8478),
            .I(beamXZ0Z_10));
    Odrv4 I__1238 (
            .O(N__8475),
            .I(beamXZ0Z_10));
    CascadeMux I__1237 (
            .O(N__8470),
            .I(N__8466));
    InMux I__1236 (
            .O(N__8469),
            .I(N__8462));
    InMux I__1235 (
            .O(N__8466),
            .I(N__8459));
    InMux I__1234 (
            .O(N__8465),
            .I(N__8456));
    LocalMux I__1233 (
            .O(N__8462),
            .I(N__8451));
    LocalMux I__1232 (
            .O(N__8459),
            .I(N__8451));
    LocalMux I__1231 (
            .O(N__8456),
            .I(N__8448));
    Span4Mux_v I__1230 (
            .O(N__8451),
            .I(N__8445));
    Odrv4 I__1229 (
            .O(N__8448),
            .I(un1_beamx_2));
    Odrv4 I__1228 (
            .O(N__8445),
            .I(un1_beamx_2));
    CascadeMux I__1227 (
            .O(N__8440),
            .I(N__8436));
    CascadeMux I__1226 (
            .O(N__8439),
            .I(N__8431));
    InMux I__1225 (
            .O(N__8436),
            .I(N__8424));
    InMux I__1224 (
            .O(N__8435),
            .I(N__8424));
    InMux I__1223 (
            .O(N__8434),
            .I(N__8421));
    InMux I__1222 (
            .O(N__8431),
            .I(N__8417));
    InMux I__1221 (
            .O(N__8430),
            .I(N__8414));
    InMux I__1220 (
            .O(N__8429),
            .I(N__8411));
    LocalMux I__1219 (
            .O(N__8424),
            .I(N__8406));
    LocalMux I__1218 (
            .O(N__8421),
            .I(N__8406));
    CascadeMux I__1217 (
            .O(N__8420),
            .I(N__8402));
    LocalMux I__1216 (
            .O(N__8417),
            .I(N__8397));
    LocalMux I__1215 (
            .O(N__8414),
            .I(N__8397));
    LocalMux I__1214 (
            .O(N__8411),
            .I(N__8394));
    Span4Mux_s2_v I__1213 (
            .O(N__8406),
            .I(N__8391));
    InMux I__1212 (
            .O(N__8405),
            .I(N__8387));
    InMux I__1211 (
            .O(N__8402),
            .I(N__8384));
    Span12Mux_s9_v I__1210 (
            .O(N__8397),
            .I(N__8381));
    Span4Mux_h I__1209 (
            .O(N__8394),
            .I(N__8376));
    Span4Mux_v I__1208 (
            .O(N__8391),
            .I(N__8376));
    InMux I__1207 (
            .O(N__8390),
            .I(N__8373));
    LocalMux I__1206 (
            .O(N__8387),
            .I(beamXZ0Z_7));
    LocalMux I__1205 (
            .O(N__8384),
            .I(beamXZ0Z_7));
    Odrv12 I__1204 (
            .O(N__8381),
            .I(beamXZ0Z_7));
    Odrv4 I__1203 (
            .O(N__8376),
            .I(beamXZ0Z_7));
    LocalMux I__1202 (
            .O(N__8373),
            .I(beamXZ0Z_7));
    InMux I__1201 (
            .O(N__8362),
            .I(N__8359));
    LocalMux I__1200 (
            .O(N__8359),
            .I(N__8356));
    Odrv12 I__1199 (
            .O(N__8356),
            .I(un1_beamxlt10_0));
    IoInMux I__1198 (
            .O(N__8353),
            .I(N__8350));
    LocalMux I__1197 (
            .O(N__8350),
            .I(N__8347));
    Span4Mux_s3_v I__1196 (
            .O(N__8347),
            .I(N__8344));
    Span4Mux_h I__1195 (
            .O(N__8344),
            .I(N__8341));
    Odrv4 I__1194 (
            .O(N__8341),
            .I(HSync_c));
    InMux I__1193 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__1192 (
            .O(N__8335),
            .I(N__8331));
    InMux I__1191 (
            .O(N__8334),
            .I(N__8328));
    Span4Mux_s2_v I__1190 (
            .O(N__8331),
            .I(N__8322));
    LocalMux I__1189 (
            .O(N__8328),
            .I(N__8319));
    InMux I__1188 (
            .O(N__8327),
            .I(N__8314));
    InMux I__1187 (
            .O(N__8326),
            .I(N__8314));
    InMux I__1186 (
            .O(N__8325),
            .I(N__8311));
    Span4Mux_v I__1185 (
            .O(N__8322),
            .I(N__8308));
    Span4Mux_s3_h I__1184 (
            .O(N__8319),
            .I(N__8303));
    LocalMux I__1183 (
            .O(N__8314),
            .I(N__8303));
    LocalMux I__1182 (
            .O(N__8311),
            .I(N__8300));
    Odrv4 I__1181 (
            .O(N__8308),
            .I(un4_row));
    Odrv4 I__1180 (
            .O(N__8303),
            .I(un4_row));
    Odrv4 I__1179 (
            .O(N__8300),
            .I(un4_row));
    CascadeMux I__1178 (
            .O(N__8293),
            .I(N__8290));
    InMux I__1177 (
            .O(N__8290),
            .I(N__8287));
    LocalMux I__1176 (
            .O(N__8287),
            .I(N__8284));
    Odrv12 I__1175 (
            .O(N__8284),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1));
    InMux I__1174 (
            .O(N__8281),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__1173 (
            .O(N__8278),
            .I(N__8275));
    InMux I__1172 (
            .O(N__8275),
            .I(N__8272));
    LocalMux I__1171 (
            .O(N__8272),
            .I(N__8269));
    Odrv4 I__1170 (
            .O(N__8269),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2));
    InMux I__1169 (
            .O(N__8266),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__1168 (
            .O(N__8263),
            .I(N__8260));
    LocalMux I__1167 (
            .O(N__8260),
            .I(N__8257));
    Odrv4 I__1166 (
            .O(N__8257),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__1165 (
            .O(N__8254),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__1164 (
            .O(N__8251),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__1163 (
            .O(N__8248),
            .I(N__8245));
    LocalMux I__1162 (
            .O(N__8245),
            .I(N__8240));
    InMux I__1161 (
            .O(N__8244),
            .I(N__8237));
    InMux I__1160 (
            .O(N__8243),
            .I(N__8234));
    Span4Mux_s1_h I__1159 (
            .O(N__8240),
            .I(N__8227));
    LocalMux I__1158 (
            .O(N__8237),
            .I(N__8227));
    LocalMux I__1157 (
            .O(N__8234),
            .I(N__8227));
    Odrv4 I__1156 (
            .O(N__8227),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2));
    CascadeMux I__1155 (
            .O(N__8224),
            .I(beamY_RNINKIU27Z0Z_0_cascade_));
    CascadeMux I__1154 (
            .O(N__8221),
            .I(Pixel_RNOZ0Z_29_cascade_));
    InMux I__1153 (
            .O(N__8218),
            .I(N__8215));
    LocalMux I__1152 (
            .O(N__8215),
            .I(N_10));
    InMux I__1151 (
            .O(N__8212),
            .I(N__8209));
    LocalMux I__1150 (
            .O(N__8209),
            .I(N__8206));
    Odrv4 I__1149 (
            .O(N__8206),
            .I(chessboardpixel_un152_pixel_27));
    CascadeMux I__1148 (
            .O(N__8203),
            .I(N__8200));
    InMux I__1147 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__1146 (
            .O(N__8197),
            .I(N__8194));
    Odrv12 I__1145 (
            .O(N__8194),
            .I(chessboardpixel_un174_pixellt10));
    InMux I__1144 (
            .O(N__8191),
            .I(N__8188));
    LocalMux I__1143 (
            .O(N__8188),
            .I(N__8185));
    Span4Mux_s3_h I__1142 (
            .O(N__8185),
            .I(N__8180));
    InMux I__1141 (
            .O(N__8184),
            .I(N__8175));
    InMux I__1140 (
            .O(N__8183),
            .I(N__8175));
    Odrv4 I__1139 (
            .O(N__8180),
            .I(chessboardpixel_un175_pixel));
    LocalMux I__1138 (
            .O(N__8175),
            .I(chessboardpixel_un175_pixel));
    InMux I__1137 (
            .O(N__8170),
            .I(N__8167));
    LocalMux I__1136 (
            .O(N__8167),
            .I(N__8164));
    Span4Mux_h I__1135 (
            .O(N__8164),
            .I(N__8161));
    Odrv4 I__1134 (
            .O(N__8161),
            .I(g1_2_1));
    CascadeMux I__1133 (
            .O(N__8158),
            .I(chessboardpixel_un175_pixel_cascade_));
    InMux I__1132 (
            .O(N__8155),
            .I(N__8152));
    LocalMux I__1131 (
            .O(N__8152),
            .I(N__8149));
    Span4Mux_s3_h I__1130 (
            .O(N__8149),
            .I(N__8146));
    Odrv4 I__1129 (
            .O(N__8146),
            .I(g2_3_0_0));
    InMux I__1128 (
            .O(N__8143),
            .I(N__8136));
    InMux I__1127 (
            .O(N__8142),
            .I(N__8136));
    InMux I__1126 (
            .O(N__8141),
            .I(N__8133));
    LocalMux I__1125 (
            .O(N__8136),
            .I(N__8130));
    LocalMux I__1124 (
            .O(N__8133),
            .I(N__8127));
    Odrv12 I__1123 (
            .O(N__8130),
            .I(un13_beamylt7));
    Odrv4 I__1122 (
            .O(N__8127),
            .I(un13_beamylt7));
    InMux I__1121 (
            .O(N__8122),
            .I(N__8118));
    InMux I__1120 (
            .O(N__8121),
            .I(N__8115));
    LocalMux I__1119 (
            .O(N__8118),
            .I(un15_beamy));
    LocalMux I__1118 (
            .O(N__8115),
            .I(un15_beamy));
    InMux I__1117 (
            .O(N__8110),
            .I(N__8107));
    LocalMux I__1116 (
            .O(N__8107),
            .I(N__8104));
    Odrv4 I__1115 (
            .O(N__8104),
            .I(un18_beamylt10_0));
    InMux I__1114 (
            .O(N__8101),
            .I(N__8097));
    InMux I__1113 (
            .O(N__8100),
            .I(N__8094));
    LocalMux I__1112 (
            .O(N__8097),
            .I(N__8089));
    LocalMux I__1111 (
            .O(N__8094),
            .I(N__8089));
    Span4Mux_s3_h I__1110 (
            .O(N__8089),
            .I(N__8084));
    InMux I__1109 (
            .O(N__8088),
            .I(N__8079));
    InMux I__1108 (
            .O(N__8087),
            .I(N__8079));
    Odrv4 I__1107 (
            .O(N__8084),
            .I(un15_beamy_2));
    LocalMux I__1106 (
            .O(N__8079),
            .I(un15_beamy_2));
    CascadeMux I__1105 (
            .O(N__8074),
            .I(Pixel_RNOZ0Z_44_cascade_));
    InMux I__1104 (
            .O(N__8071),
            .I(N__8068));
    LocalMux I__1103 (
            .O(N__8068),
            .I(N__8065));
    Span12Mux_s3_h I__1102 (
            .O(N__8065),
            .I(N__8062));
    Odrv12 I__1101 (
            .O(N__8062),
            .I(N_10_0_0));
    InMux I__1100 (
            .O(N__8059),
            .I(N__8056));
    LocalMux I__1099 (
            .O(N__8056),
            .I(N__8053));
    Span4Mux_h I__1098 (
            .O(N__8053),
            .I(N__8050));
    Odrv4 I__1097 (
            .O(N__8050),
            .I(N_20));
    CascadeMux I__1096 (
            .O(N__8047),
            .I(g0_4_cascade_));
    InMux I__1095 (
            .O(N__8044),
            .I(N__8041));
    LocalMux I__1094 (
            .O(N__8041),
            .I(N__8038));
    Odrv4 I__1093 (
            .O(N__8038),
            .I(G_21_i_2));
    IoInMux I__1092 (
            .O(N__8035),
            .I(N__8032));
    LocalMux I__1091 (
            .O(N__8032),
            .I(N__8029));
    Span4Mux_s1_v I__1090 (
            .O(N__8029),
            .I(N__8026));
    Span4Mux_h I__1089 (
            .O(N__8026),
            .I(N__8023));
    Odrv4 I__1088 (
            .O(N__8023),
            .I(Pixel_c));
    InMux I__1087 (
            .O(N__8020),
            .I(N__8017));
    LocalMux I__1086 (
            .O(N__8017),
            .I(g1_1_0));
    InMux I__1085 (
            .O(N__8014),
            .I(N__8011));
    LocalMux I__1084 (
            .O(N__8011),
            .I(N__8008));
    Odrv12 I__1083 (
            .O(N__8008),
            .I(g0_2_0));
    CascadeMux I__1082 (
            .O(N__8005),
            .I(g1_1_cascade_));
    InMux I__1081 (
            .O(N__8002),
            .I(N__7999));
    LocalMux I__1080 (
            .O(N__7999),
            .I(g3_1));
    InMux I__1079 (
            .O(N__7996),
            .I(N__7993));
    LocalMux I__1078 (
            .O(N__7993),
            .I(g0_5));
    InMux I__1077 (
            .O(N__7990),
            .I(N__7986));
    InMux I__1076 (
            .O(N__7989),
            .I(N__7983));
    LocalMux I__1075 (
            .O(N__7986),
            .I(g1_0_0));
    LocalMux I__1074 (
            .O(N__7983),
            .I(g1_0_0));
    CascadeMux I__1073 (
            .O(N__7978),
            .I(N__7975));
    InMux I__1072 (
            .O(N__7975),
            .I(N__7972));
    LocalMux I__1071 (
            .O(N__7972),
            .I(N__7969));
    Odrv12 I__1070 (
            .O(N__7969),
            .I(g0_0_a3_0));
    InMux I__1069 (
            .O(N__7966),
            .I(N__7957));
    InMux I__1068 (
            .O(N__7965),
            .I(N__7952));
    InMux I__1067 (
            .O(N__7964),
            .I(N__7952));
    CascadeMux I__1066 (
            .O(N__7963),
            .I(N__7949));
    InMux I__1065 (
            .O(N__7962),
            .I(N__7945));
    InMux I__1064 (
            .O(N__7961),
            .I(N__7940));
    InMux I__1063 (
            .O(N__7960),
            .I(N__7940));
    LocalMux I__1062 (
            .O(N__7957),
            .I(N__7934));
    LocalMux I__1061 (
            .O(N__7952),
            .I(N__7934));
    InMux I__1060 (
            .O(N__7949),
            .I(N__7931));
    InMux I__1059 (
            .O(N__7948),
            .I(N__7927));
    LocalMux I__1058 (
            .O(N__7945),
            .I(N__7922));
    LocalMux I__1057 (
            .O(N__7940),
            .I(N__7922));
    InMux I__1056 (
            .O(N__7939),
            .I(N__7919));
    Span4Mux_s2_v I__1055 (
            .O(N__7934),
            .I(N__7914));
    LocalMux I__1054 (
            .O(N__7931),
            .I(N__7914));
    CascadeMux I__1053 (
            .O(N__7930),
            .I(N__7910));
    LocalMux I__1052 (
            .O(N__7927),
            .I(N__7903));
    Span4Mux_s2_v I__1051 (
            .O(N__7922),
            .I(N__7903));
    LocalMux I__1050 (
            .O(N__7919),
            .I(N__7903));
    Span4Mux_v I__1049 (
            .O(N__7914),
            .I(N__7900));
    CascadeMux I__1048 (
            .O(N__7913),
            .I(N__7896));
    InMux I__1047 (
            .O(N__7910),
            .I(N__7890));
    Span4Mux_v I__1046 (
            .O(N__7903),
            .I(N__7887));
    Span4Mux_v I__1045 (
            .O(N__7900),
            .I(N__7884));
    InMux I__1044 (
            .O(N__7899),
            .I(N__7875));
    InMux I__1043 (
            .O(N__7896),
            .I(N__7875));
    InMux I__1042 (
            .O(N__7895),
            .I(N__7875));
    InMux I__1041 (
            .O(N__7894),
            .I(N__7875));
    InMux I__1040 (
            .O(N__7893),
            .I(N__7872));
    LocalMux I__1039 (
            .O(N__7890),
            .I(beamXZ0Z_0));
    Odrv4 I__1038 (
            .O(N__7887),
            .I(beamXZ0Z_0));
    Odrv4 I__1037 (
            .O(N__7884),
            .I(beamXZ0Z_0));
    LocalMux I__1036 (
            .O(N__7875),
            .I(beamXZ0Z_0));
    LocalMux I__1035 (
            .O(N__7872),
            .I(beamXZ0Z_0));
    CascadeMux I__1034 (
            .O(N__7861),
            .I(N__7858));
    InMux I__1033 (
            .O(N__7858),
            .I(N__7855));
    LocalMux I__1032 (
            .O(N__7855),
            .I(N__7852));
    Odrv4 I__1031 (
            .O(N__7852),
            .I(N_35));
    InMux I__1030 (
            .O(N__7849),
            .I(N__7846));
    LocalMux I__1029 (
            .O(N__7846),
            .I(N__7843));
    Odrv4 I__1028 (
            .O(N__7843),
            .I(N_58_mux));
    InMux I__1027 (
            .O(N__7840),
            .I(N__7834));
    InMux I__1026 (
            .O(N__7839),
            .I(N__7831));
    InMux I__1025 (
            .O(N__7838),
            .I(N__7826));
    InMux I__1024 (
            .O(N__7837),
            .I(N__7826));
    LocalMux I__1023 (
            .O(N__7834),
            .I(N__7816));
    LocalMux I__1022 (
            .O(N__7831),
            .I(N__7816));
    LocalMux I__1021 (
            .O(N__7826),
            .I(N__7809));
    CascadeMux I__1020 (
            .O(N__7825),
            .I(N__7805));
    InMux I__1019 (
            .O(N__7824),
            .I(N__7800));
    InMux I__1018 (
            .O(N__7823),
            .I(N__7800));
    InMux I__1017 (
            .O(N__7822),
            .I(N__7795));
    InMux I__1016 (
            .O(N__7821),
            .I(N__7795));
    Span4Mux_s3_v I__1015 (
            .O(N__7816),
            .I(N__7792));
    InMux I__1014 (
            .O(N__7815),
            .I(N__7783));
    InMux I__1013 (
            .O(N__7814),
            .I(N__7783));
    InMux I__1012 (
            .O(N__7813),
            .I(N__7783));
    InMux I__1011 (
            .O(N__7812),
            .I(N__7783));
    Span4Mux_h I__1010 (
            .O(N__7809),
            .I(N__7780));
    InMux I__1009 (
            .O(N__7808),
            .I(N__7775));
    InMux I__1008 (
            .O(N__7805),
            .I(N__7775));
    LocalMux I__1007 (
            .O(N__7800),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__1006 (
            .O(N__7795),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    Odrv4 I__1005 (
            .O(N__7792),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__1004 (
            .O(N__7783),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    Odrv4 I__1003 (
            .O(N__7780),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__1002 (
            .O(N__7775),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    CascadeMux I__1001 (
            .O(N__7762),
            .I(beamY_RNIDQG2Z0Z_0_cascade_));
    InMux I__1000 (
            .O(N__7759),
            .I(N__7753));
    InMux I__999 (
            .O(N__7758),
            .I(N__7748));
    InMux I__998 (
            .O(N__7757),
            .I(N__7748));
    InMux I__997 (
            .O(N__7756),
            .I(N__7742));
    LocalMux I__996 (
            .O(N__7753),
            .I(N__7734));
    LocalMux I__995 (
            .O(N__7748),
            .I(N__7731));
    InMux I__994 (
            .O(N__7747),
            .I(N__7724));
    InMux I__993 (
            .O(N__7746),
            .I(N__7724));
    InMux I__992 (
            .O(N__7745),
            .I(N__7724));
    LocalMux I__991 (
            .O(N__7742),
            .I(N__7721));
    InMux I__990 (
            .O(N__7741),
            .I(N__7714));
    InMux I__989 (
            .O(N__7740),
            .I(N__7714));
    InMux I__988 (
            .O(N__7739),
            .I(N__7714));
    InMux I__987 (
            .O(N__7738),
            .I(N__7709));
    InMux I__986 (
            .O(N__7737),
            .I(N__7709));
    Span4Mux_h I__985 (
            .O(N__7734),
            .I(N__7706));
    Span4Mux_h I__984 (
            .O(N__7731),
            .I(N__7703));
    LocalMux I__983 (
            .O(N__7724),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    Odrv4 I__982 (
            .O(N__7721),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    LocalMux I__981 (
            .O(N__7714),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    LocalMux I__980 (
            .O(N__7709),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    Odrv4 I__979 (
            .O(N__7706),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    Odrv4 I__978 (
            .O(N__7703),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    InMux I__977 (
            .O(N__7690),
            .I(N__7687));
    LocalMux I__976 (
            .O(N__7687),
            .I(N__7684));
    Odrv4 I__975 (
            .O(N__7684),
            .I(beamY_RNINKIU27Z0Z_0));
    InMux I__974 (
            .O(N__7681),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7));
    CascadeMux I__973 (
            .O(N__7678),
            .I(g2_1_cascade_));
    CascadeMux I__972 (
            .O(N__7675),
            .I(N_7_cascade_));
    InMux I__971 (
            .O(N__7672),
            .I(N__7669));
    LocalMux I__970 (
            .O(N__7669),
            .I(g2_1));
    CascadeMux I__969 (
            .O(N__7666),
            .I(g0_1_0_cascade_));
    CascadeMux I__968 (
            .O(N__7663),
            .I(g0_1_3_cascade_));
    CascadeMux I__967 (
            .O(N__7660),
            .I(g3_2_2_cascade_));
    CascadeMux I__966 (
            .O(N__7657),
            .I(N__7654));
    InMux I__965 (
            .O(N__7654),
            .I(N__7651));
    LocalMux I__964 (
            .O(N__7651),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538));
    InMux I__963 (
            .O(N__7648),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__962 (
            .O(N__7645),
            .I(N__7642));
    LocalMux I__961 (
            .O(N__7642),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO));
    InMux I__960 (
            .O(N__7639),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__959 (
            .O(N__7636),
            .I(N__7633));
    InMux I__958 (
            .O(N__7633),
            .I(N__7630));
    LocalMux I__957 (
            .O(N__7630),
            .I(un5_visiblex_i_24));
    InMux I__956 (
            .O(N__7627),
            .I(N__7624));
    LocalMux I__955 (
            .O(N__7624),
            .I(charx_if_generate_plus_mult1_un26_sum_i_5));
    InMux I__954 (
            .O(N__7621),
            .I(N__7615));
    InMux I__953 (
            .O(N__7620),
            .I(N__7615));
    LocalMux I__952 (
            .O(N__7615),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    InMux I__951 (
            .O(N__7612),
            .I(N__7603));
    InMux I__950 (
            .O(N__7611),
            .I(N__7603));
    InMux I__949 (
            .O(N__7610),
            .I(N__7603));
    LocalMux I__948 (
            .O(N__7603),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    InMux I__947 (
            .O(N__7600),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__946 (
            .O(N__7597),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__945 (
            .O(N__7594),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__944 (
            .O(N__7591),
            .I(un8_beamx_cry_9));
    CascadeMux I__943 (
            .O(N__7588),
            .I(N__7585));
    InMux I__942 (
            .O(N__7585),
            .I(N__7579));
    InMux I__941 (
            .O(N__7584),
            .I(N__7575));
    CascadeMux I__940 (
            .O(N__7583),
            .I(N__7571));
    InMux I__939 (
            .O(N__7582),
            .I(N__7568));
    LocalMux I__938 (
            .O(N__7579),
            .I(N__7565));
    InMux I__937 (
            .O(N__7578),
            .I(N__7562));
    LocalMux I__936 (
            .O(N__7575),
            .I(N__7559));
    InMux I__935 (
            .O(N__7574),
            .I(N__7555));
    InMux I__934 (
            .O(N__7571),
            .I(N__7552));
    LocalMux I__933 (
            .O(N__7568),
            .I(N__7549));
    Span4Mux_h I__932 (
            .O(N__7565),
            .I(N__7542));
    LocalMux I__931 (
            .O(N__7562),
            .I(N__7542));
    Span4Mux_s1_h I__930 (
            .O(N__7559),
            .I(N__7542));
    InMux I__929 (
            .O(N__7558),
            .I(N__7539));
    LocalMux I__928 (
            .O(N__7555),
            .I(beamXZ0Z_4));
    LocalMux I__927 (
            .O(N__7552),
            .I(beamXZ0Z_4));
    Odrv12 I__926 (
            .O(N__7549),
            .I(beamXZ0Z_4));
    Odrv4 I__925 (
            .O(N__7542),
            .I(beamXZ0Z_4));
    LocalMux I__924 (
            .O(N__7539),
            .I(beamXZ0Z_4));
    CascadeMux I__923 (
            .O(N__7528),
            .I(N__7525));
    InMux I__922 (
            .O(N__7525),
            .I(N__7518));
    InMux I__921 (
            .O(N__7524),
            .I(N__7514));
    InMux I__920 (
            .O(N__7523),
            .I(N__7511));
    InMux I__919 (
            .O(N__7522),
            .I(N__7508));
    InMux I__918 (
            .O(N__7521),
            .I(N__7505));
    LocalMux I__917 (
            .O(N__7518),
            .I(N__7502));
    InMux I__916 (
            .O(N__7517),
            .I(N__7498));
    LocalMux I__915 (
            .O(N__7514),
            .I(N__7491));
    LocalMux I__914 (
            .O(N__7511),
            .I(N__7491));
    LocalMux I__913 (
            .O(N__7508),
            .I(N__7491));
    LocalMux I__912 (
            .O(N__7505),
            .I(N__7486));
    Span12Mux_s9_v I__911 (
            .O(N__7502),
            .I(N__7486));
    InMux I__910 (
            .O(N__7501),
            .I(N__7483));
    LocalMux I__909 (
            .O(N__7498),
            .I(beamXZ0Z_6));
    Odrv12 I__908 (
            .O(N__7491),
            .I(beamXZ0Z_6));
    Odrv12 I__907 (
            .O(N__7486),
            .I(beamXZ0Z_6));
    LocalMux I__906 (
            .O(N__7483),
            .I(beamXZ0Z_6));
    InMux I__905 (
            .O(N__7474),
            .I(N__7471));
    LocalMux I__904 (
            .O(N__7471),
            .I(un3_beamx_5));
    InMux I__903 (
            .O(N__7468),
            .I(N__7465));
    LocalMux I__902 (
            .O(N__7465),
            .I(N__7462));
    Odrv4 I__901 (
            .O(N__7462),
            .I(un3_beamx_7));
    InMux I__900 (
            .O(N__7459),
            .I(N__7453));
    InMux I__899 (
            .O(N__7458),
            .I(N__7448));
    InMux I__898 (
            .O(N__7457),
            .I(N__7448));
    InMux I__897 (
            .O(N__7456),
            .I(N__7445));
    LocalMux I__896 (
            .O(N__7453),
            .I(beamXZ0Z_2));
    LocalMux I__895 (
            .O(N__7448),
            .I(beamXZ0Z_2));
    LocalMux I__894 (
            .O(N__7445),
            .I(beamXZ0Z_2));
    InMux I__893 (
            .O(N__7438),
            .I(N__7432));
    CascadeMux I__892 (
            .O(N__7437),
            .I(N__7429));
    CascadeMux I__891 (
            .O(N__7436),
            .I(N__7426));
    InMux I__890 (
            .O(N__7435),
            .I(N__7422));
    LocalMux I__889 (
            .O(N__7432),
            .I(N__7419));
    InMux I__888 (
            .O(N__7429),
            .I(N__7416));
    InMux I__887 (
            .O(N__7426),
            .I(N__7413));
    InMux I__886 (
            .O(N__7425),
            .I(N__7410));
    LocalMux I__885 (
            .O(N__7422),
            .I(beamXZ0Z_3));
    Odrv12 I__884 (
            .O(N__7419),
            .I(beamXZ0Z_3));
    LocalMux I__883 (
            .O(N__7416),
            .I(beamXZ0Z_3));
    LocalMux I__882 (
            .O(N__7413),
            .I(beamXZ0Z_3));
    LocalMux I__881 (
            .O(N__7410),
            .I(beamXZ0Z_3));
    CascadeMux I__880 (
            .O(N__7399),
            .I(N__7395));
    CascadeMux I__879 (
            .O(N__7398),
            .I(N__7392));
    InMux I__878 (
            .O(N__7395),
            .I(N__7388));
    InMux I__877 (
            .O(N__7392),
            .I(N__7385));
    InMux I__876 (
            .O(N__7391),
            .I(N__7382));
    LocalMux I__875 (
            .O(N__7388),
            .I(N__7375));
    LocalMux I__874 (
            .O(N__7385),
            .I(N__7375));
    LocalMux I__873 (
            .O(N__7382),
            .I(N__7375));
    Span4Mux_v I__872 (
            .O(N__7375),
            .I(N__7372));
    Odrv4 I__871 (
            .O(N__7372),
            .I(un18_beamylt4));
    InMux I__870 (
            .O(N__7369),
            .I(N__7362));
    InMux I__869 (
            .O(N__7368),
            .I(N__7355));
    InMux I__868 (
            .O(N__7367),
            .I(N__7355));
    InMux I__867 (
            .O(N__7366),
            .I(N__7355));
    InMux I__866 (
            .O(N__7365),
            .I(N__7352));
    LocalMux I__865 (
            .O(N__7362),
            .I(beamXZ0Z_1));
    LocalMux I__864 (
            .O(N__7355),
            .I(beamXZ0Z_1));
    LocalMux I__863 (
            .O(N__7352),
            .I(beamXZ0Z_1));
    InMux I__862 (
            .O(N__7345),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1));
    CascadeMux I__861 (
            .O(N__7342),
            .I(N__7339));
    InMux I__860 (
            .O(N__7339),
            .I(N__7336));
    LocalMux I__859 (
            .O(N__7336),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328));
    InMux I__858 (
            .O(N__7333),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__857 (
            .O(N__7330),
            .I(un8_beamx_cry_1));
    InMux I__856 (
            .O(N__7327),
            .I(un8_beamx_cry_2));
    InMux I__855 (
            .O(N__7324),
            .I(un8_beamx_cry_3));
    InMux I__854 (
            .O(N__7321),
            .I(N__7315));
    InMux I__853 (
            .O(N__7320),
            .I(N__7310));
    InMux I__852 (
            .O(N__7319),
            .I(N__7307));
    InMux I__851 (
            .O(N__7318),
            .I(N__7304));
    LocalMux I__850 (
            .O(N__7315),
            .I(N__7301));
    InMux I__849 (
            .O(N__7314),
            .I(N__7297));
    InMux I__848 (
            .O(N__7313),
            .I(N__7294));
    LocalMux I__847 (
            .O(N__7310),
            .I(N__7289));
    LocalMux I__846 (
            .O(N__7307),
            .I(N__7289));
    LocalMux I__845 (
            .O(N__7304),
            .I(N__7284));
    Span4Mux_s1_h I__844 (
            .O(N__7301),
            .I(N__7284));
    InMux I__843 (
            .O(N__7300),
            .I(N__7281));
    LocalMux I__842 (
            .O(N__7297),
            .I(beamXZ0Z_5));
    LocalMux I__841 (
            .O(N__7294),
            .I(beamXZ0Z_5));
    Odrv12 I__840 (
            .O(N__7289),
            .I(beamXZ0Z_5));
    Odrv4 I__839 (
            .O(N__7284),
            .I(beamXZ0Z_5));
    LocalMux I__838 (
            .O(N__7281),
            .I(beamXZ0Z_5));
    InMux I__837 (
            .O(N__7270),
            .I(un8_beamx_cry_4));
    InMux I__836 (
            .O(N__7267),
            .I(un8_beamx_cry_5));
    InMux I__835 (
            .O(N__7264),
            .I(un8_beamx_cry_6));
    InMux I__834 (
            .O(N__7261),
            .I(N__7252));
    InMux I__833 (
            .O(N__7260),
            .I(N__7252));
    InMux I__832 (
            .O(N__7259),
            .I(N__7249));
    InMux I__831 (
            .O(N__7258),
            .I(N__7244));
    InMux I__830 (
            .O(N__7257),
            .I(N__7244));
    LocalMux I__829 (
            .O(N__7252),
            .I(N__7239));
    LocalMux I__828 (
            .O(N__7249),
            .I(N__7239));
    LocalMux I__827 (
            .O(N__7244),
            .I(N__7232));
    Span4Mux_v I__826 (
            .O(N__7239),
            .I(N__7232));
    InMux I__825 (
            .O(N__7238),
            .I(N__7229));
    InMux I__824 (
            .O(N__7237),
            .I(N__7226));
    Span4Mux_v I__823 (
            .O(N__7232),
            .I(N__7221));
    LocalMux I__822 (
            .O(N__7229),
            .I(N__7221));
    LocalMux I__821 (
            .O(N__7226),
            .I(beamXZ0Z_8));
    Odrv4 I__820 (
            .O(N__7221),
            .I(beamXZ0Z_8));
    InMux I__819 (
            .O(N__7216),
            .I(un8_beamx_cry_7));
    InMux I__818 (
            .O(N__7213),
            .I(N__7204));
    InMux I__817 (
            .O(N__7212),
            .I(N__7204));
    InMux I__816 (
            .O(N__7211),
            .I(N__7201));
    InMux I__815 (
            .O(N__7210),
            .I(N__7195));
    InMux I__814 (
            .O(N__7209),
            .I(N__7195));
    LocalMux I__813 (
            .O(N__7204),
            .I(N__7190));
    LocalMux I__812 (
            .O(N__7201),
            .I(N__7190));
    InMux I__811 (
            .O(N__7200),
            .I(N__7186));
    LocalMux I__810 (
            .O(N__7195),
            .I(N__7181));
    Sp12to4 I__809 (
            .O(N__7190),
            .I(N__7181));
    InMux I__808 (
            .O(N__7189),
            .I(N__7178));
    LocalMux I__807 (
            .O(N__7186),
            .I(beamXZ0Z_9));
    Odrv12 I__806 (
            .O(N__7181),
            .I(beamXZ0Z_9));
    LocalMux I__805 (
            .O(N__7178),
            .I(beamXZ0Z_9));
    InMux I__804 (
            .O(N__7171),
            .I(bfn_2_11_0_));
    InMux I__803 (
            .O(N__7168),
            .I(N__7162));
    InMux I__802 (
            .O(N__7167),
            .I(N__7162));
    LocalMux I__801 (
            .O(N__7162),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__800 (
            .O(N__7159),
            .I(N__7156));
    InMux I__799 (
            .O(N__7156),
            .I(N__7153));
    LocalMux I__798 (
            .O(N__7153),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7));
    InMux I__797 (
            .O(N__7150),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1));
    CascadeMux I__796 (
            .O(N__7147),
            .I(N__7144));
    InMux I__795 (
            .O(N__7144),
            .I(N__7141));
    LocalMux I__794 (
            .O(N__7141),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0));
    InMux I__793 (
            .O(N__7138),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__792 (
            .O(N__7135),
            .I(N__7132));
    LocalMux I__791 (
            .O(N__7132),
            .I(charx_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__790 (
            .O(N__7129),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__789 (
            .O(N__7126),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__788 (
            .O(N__7123),
            .I(N__7119));
    InMux I__787 (
            .O(N__7122),
            .I(N__7116));
    LocalMux I__786 (
            .O(N__7119),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0));
    LocalMux I__785 (
            .O(N__7116),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0));
    CascadeMux I__784 (
            .O(N__7111),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_));
    InMux I__783 (
            .O(N__7108),
            .I(N__7102));
    InMux I__782 (
            .O(N__7107),
            .I(N__7102));
    LocalMux I__781 (
            .O(N__7102),
            .I(charx_if_generate_plus_mult1_un61_sum_i_5));
    CascadeMux I__780 (
            .O(N__7099),
            .I(N__7096));
    InMux I__779 (
            .O(N__7096),
            .I(N__7093));
    LocalMux I__778 (
            .O(N__7093),
            .I(charx_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__777 (
            .O(N__7090),
            .I(un13_beamylt7_0_cascade_));
    InMux I__776 (
            .O(N__7087),
            .I(N__7084));
    LocalMux I__775 (
            .O(N__7084),
            .I(N__7081));
    Odrv4 I__774 (
            .O(N__7081),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0));
    InMux I__773 (
            .O(N__7078),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__772 (
            .O(N__7075),
            .I(N__7072));
    InMux I__771 (
            .O(N__7072),
            .I(N__7069));
    LocalMux I__770 (
            .O(N__7069),
            .I(N__7066));
    Odrv4 I__769 (
            .O(N__7066),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0));
    InMux I__768 (
            .O(N__7063),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__767 (
            .O(N__7060),
            .I(N__7057));
    LocalMux I__766 (
            .O(N__7057),
            .I(N__7054));
    Odrv4 I__765 (
            .O(N__7054),
            .I(charx_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__764 (
            .O(N__7051),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__763 (
            .O(N__7048),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__762 (
            .O(N__7045),
            .I(N__7042));
    InMux I__761 (
            .O(N__7042),
            .I(N__7035));
    InMux I__760 (
            .O(N__7041),
            .I(N__7035));
    InMux I__759 (
            .O(N__7040),
            .I(N__7032));
    LocalMux I__758 (
            .O(N__7035),
            .I(N__7029));
    LocalMux I__757 (
            .O(N__7032),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0));
    Odrv4 I__756 (
            .O(N__7029),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0));
    CascadeMux I__755 (
            .O(N__7024),
            .I(N__7021));
    InMux I__754 (
            .O(N__7021),
            .I(N__7018));
    LocalMux I__753 (
            .O(N__7018),
            .I(charx_if_generate_plus_mult1_un61_sum_i));
    InMux I__752 (
            .O(N__7015),
            .I(N__7012));
    LocalMux I__751 (
            .O(N__7012),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0));
    CascadeMux I__750 (
            .O(N__7009),
            .I(N__7004));
    InMux I__749 (
            .O(N__7008),
            .I(N__6999));
    InMux I__748 (
            .O(N__7007),
            .I(N__6994));
    InMux I__747 (
            .O(N__7004),
            .I(N__6994));
    InMux I__746 (
            .O(N__7003),
            .I(N__6991));
    InMux I__745 (
            .O(N__7002),
            .I(N__6988));
    LocalMux I__744 (
            .O(N__6999),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    LocalMux I__743 (
            .O(N__6994),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    LocalMux I__742 (
            .O(N__6991),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    LocalMux I__741 (
            .O(N__6988),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    InMux I__740 (
            .O(N__6979),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__739 (
            .O(N__6976),
            .I(N__6971));
    InMux I__738 (
            .O(N__6975),
            .I(N__6968));
    InMux I__737 (
            .O(N__6974),
            .I(N__6965));
    LocalMux I__736 (
            .O(N__6971),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1));
    LocalMux I__735 (
            .O(N__6968),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1));
    LocalMux I__734 (
            .O(N__6965),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1));
    InMux I__733 (
            .O(N__6958),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__732 (
            .O(N__6955),
            .I(N__6949));
    InMux I__731 (
            .O(N__6954),
            .I(N__6949));
    LocalMux I__730 (
            .O(N__6949),
            .I(charx_if_generate_plus_mult1_un68_sum_i_5));
    InMux I__729 (
            .O(N__6946),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__728 (
            .O(N__6943),
            .I(N__6940));
    LocalMux I__727 (
            .O(N__6940),
            .I(N__6932));
    InMux I__726 (
            .O(N__6939),
            .I(N__6925));
    InMux I__725 (
            .O(N__6938),
            .I(N__6925));
    InMux I__724 (
            .O(N__6937),
            .I(N__6925));
    InMux I__723 (
            .O(N__6936),
            .I(N__6920));
    InMux I__722 (
            .O(N__6935),
            .I(N__6920));
    Odrv4 I__721 (
            .O(N__6932),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1));
    LocalMux I__720 (
            .O(N__6925),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1));
    LocalMux I__719 (
            .O(N__6920),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1));
    CascadeMux I__718 (
            .O(N__6913),
            .I(N__6910));
    InMux I__717 (
            .O(N__6910),
            .I(N__6907));
    LocalMux I__716 (
            .O(N__6907),
            .I(charx_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__715 (
            .O(N__6904),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_));
    InMux I__714 (
            .O(N__6901),
            .I(N__6898));
    LocalMux I__713 (
            .O(N__6898),
            .I(font_un126_pixel_5_a0_2));
    CascadeMux I__712 (
            .O(N__6895),
            .I(G_19_i_a11_0_1_cascade_));
    InMux I__711 (
            .O(N__6892),
            .I(N__6889));
    LocalMux I__710 (
            .O(N__6889),
            .I(Pixel_RNOZ0Z_36));
    CascadeMux I__709 (
            .O(N__6886),
            .I(g1_1_0_0_cascade_));
    InMux I__708 (
            .O(N__6883),
            .I(N__6880));
    LocalMux I__707 (
            .O(N__6880),
            .I(g0_0));
    InMux I__706 (
            .O(N__6877),
            .I(N__6873));
    InMux I__705 (
            .O(N__6876),
            .I(N__6870));
    LocalMux I__704 (
            .O(N__6873),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    LocalMux I__703 (
            .O(N__6870),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    InMux I__702 (
            .O(N__6865),
            .I(N__6862));
    LocalMux I__701 (
            .O(N__6862),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0));
    CascadeMux I__700 (
            .O(N__6859),
            .I(N__6855));
    CascadeMux I__699 (
            .O(N__6858),
            .I(N__6852));
    InMux I__698 (
            .O(N__6855),
            .I(N__6847));
    InMux I__697 (
            .O(N__6852),
            .I(N__6847));
    LocalMux I__696 (
            .O(N__6847),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0));
    InMux I__695 (
            .O(N__6844),
            .I(N__6838));
    InMux I__694 (
            .O(N__6843),
            .I(N__6838));
    LocalMux I__693 (
            .O(N__6838),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0));
    CascadeMux I__692 (
            .O(N__6835),
            .I(g3_3_cascade_));
    CascadeMux I__691 (
            .O(N__6832),
            .I(g0_0_2_cascade_));
    CascadeMux I__690 (
            .O(N__6829),
            .I(g0_3_cascade_));
    InMux I__689 (
            .O(N__6826),
            .I(N__6823));
    LocalMux I__688 (
            .O(N__6823),
            .I(N_21_0));
    InMux I__687 (
            .O(N__6820),
            .I(N__6817));
    LocalMux I__686 (
            .O(N__6817),
            .I(Pixel_RNOZ0Z_37));
    CascadeMux I__685 (
            .O(N__6814),
            .I(font_un126_pixel_m_2_1_1_cascade_));
    InMux I__684 (
            .O(N__6811),
            .I(N__6808));
    LocalMux I__683 (
            .O(N__6808),
            .I(Pixel_RNOZ0Z_71));
    InMux I__682 (
            .O(N__6805),
            .I(N__6802));
    LocalMux I__681 (
            .O(N__6802),
            .I(g0_0_1));
    InMux I__680 (
            .O(N__6799),
            .I(N__6796));
    LocalMux I__679 (
            .O(N__6796),
            .I(font_un3_pixel_29));
    CascadeMux I__678 (
            .O(N__6793),
            .I(font_un126_pixel_m_2_1_cascade_));
    InMux I__677 (
            .O(N__6790),
            .I(N__6787));
    LocalMux I__676 (
            .O(N__6787),
            .I(g2_2_0_1));
    InMux I__675 (
            .O(N__6784),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__674 (
            .O(N__6781),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__673 (
            .O(N__6778),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4));
    InMux I__672 (
            .O(N__6775),
            .I(N__6772));
    LocalMux I__671 (
            .O(N__6772),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_1));
    InMux I__670 (
            .O(N__6769),
            .I(N__6766));
    LocalMux I__669 (
            .O(N__6766),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3_i));
    CascadeMux I__668 (
            .O(N__6763),
            .I(g1_2_cascade_));
    CascadeMux I__667 (
            .O(N__6760),
            .I(g2_3_0_cascade_));
    InMux I__666 (
            .O(N__6757),
            .I(N__6754));
    LocalMux I__665 (
            .O(N__6754),
            .I(g2_2_0));
    InMux I__664 (
            .O(N__6751),
            .I(un5_visiblex_cry_2));
    InMux I__663 (
            .O(N__6748),
            .I(un5_visiblex_cry_3));
    InMux I__662 (
            .O(N__6745),
            .I(un5_visiblex_cry_4));
    InMux I__661 (
            .O(N__6742),
            .I(un5_visiblex_cry_5));
    InMux I__660 (
            .O(N__6739),
            .I(un5_visiblex_cry_6));
    InMux I__659 (
            .O(N__6736),
            .I(bfn_1_12_0_));
    InMux I__658 (
            .O(N__6733),
            .I(un5_visiblex_cry_8));
    InMux I__657 (
            .O(N__6730),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1));
    CascadeMux I__656 (
            .O(N__6727),
            .I(N__6724));
    InMux I__655 (
            .O(N__6724),
            .I(N__6721));
    LocalMux I__654 (
            .O(N__6721),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__653 (
            .O(N__6718),
            .I(N__6715));
    InMux I__652 (
            .O(N__6715),
            .I(N__6712));
    LocalMux I__651 (
            .O(N__6712),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i));
    InMux I__650 (
            .O(N__6709),
            .I(un5_visiblex_cry_0));
    InMux I__649 (
            .O(N__6706),
            .I(un5_visiblex_cry_1));
    InMux I__648 (
            .O(N__6703),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__647 (
            .O(N__6700),
            .I(N__6695));
    InMux I__646 (
            .O(N__6699),
            .I(N__6692));
    InMux I__645 (
            .O(N__6698),
            .I(N__6689));
    LocalMux I__644 (
            .O(N__6695),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0));
    LocalMux I__643 (
            .O(N__6692),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0));
    LocalMux I__642 (
            .O(N__6689),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0));
    CascadeMux I__641 (
            .O(N__6682),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_));
    InMux I__640 (
            .O(N__6679),
            .I(N__6676));
    LocalMux I__639 (
            .O(N__6676),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__638 (
            .O(N__6673),
            .I(N__6667));
    InMux I__637 (
            .O(N__6672),
            .I(N__6667));
    LocalMux I__636 (
            .O(N__6667),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__635 (
            .O(N__6664),
            .I(N__6661));
    InMux I__634 (
            .O(N__6661),
            .I(N__6658));
    LocalMux I__633 (
            .O(N__6658),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93));
    InMux I__632 (
            .O(N__6655),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__631 (
            .O(N__6652),
            .I(N__6649));
    InMux I__630 (
            .O(N__6649),
            .I(N__6646));
    LocalMux I__629 (
            .O(N__6646),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4));
    InMux I__628 (
            .O(N__6643),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__627 (
            .O(N__6640),
            .I(N__6637));
    LocalMux I__626 (
            .O(N__6637),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__625 (
            .O(N__6634),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__624 (
            .O(N__6631),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__623 (
            .O(N__6628),
            .I(N__6623));
    InMux I__622 (
            .O(N__6627),
            .I(N__6618));
    InMux I__621 (
            .O(N__6626),
            .I(N__6618));
    LocalMux I__620 (
            .O(N__6623),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36));
    LocalMux I__619 (
            .O(N__6618),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36));
    InMux I__618 (
            .O(N__6613),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__617 (
            .O(N__6610),
            .I(N__6607));
    LocalMux I__616 (
            .O(N__6607),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0));
    InMux I__615 (
            .O(N__6604),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__614 (
            .O(N__6601),
            .I(N__6598));
    InMux I__613 (
            .O(N__6598),
            .I(N__6595));
    LocalMux I__612 (
            .O(N__6595),
            .I(N__6592));
    Odrv12 I__611 (
            .O(N__6592),
            .I(un18_beamylto9_2));
    CascadeMux I__610 (
            .O(N__6589),
            .I(N__6586));
    InMux I__609 (
            .O(N__6586),
            .I(N__6583));
    LocalMux I__608 (
            .O(N__6583),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__607 (
            .O(N__6580),
            .I(N__6577));
    InMux I__606 (
            .O(N__6577),
            .I(N__6574));
    LocalMux I__605 (
            .O(N__6574),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6));
    InMux I__604 (
            .O(N__6571),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__603 (
            .O(N__6568),
            .I(N__6565));
    InMux I__602 (
            .O(N__6565),
            .I(N__6562));
    LocalMux I__601 (
            .O(N__6562),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9));
    InMux I__600 (
            .O(N__6559),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__599 (
            .O(N__6556),
            .I(N__6553));
    LocalMux I__598 (
            .O(N__6553),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__597 (
            .O(N__6550),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__596 (
            .O(N__6547),
            .I(N__6544));
    LocalMux I__595 (
            .O(N__6544),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3));
    InMux I__594 (
            .O(N__6541),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1));
    CascadeMux I__593 (
            .O(N__6538),
            .I(N__6535));
    InMux I__592 (
            .O(N__6535),
            .I(N__6532));
    LocalMux I__591 (
            .O(N__6532),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3));
    InMux I__590 (
            .O(N__6529),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2));
    CascadeMux I__589 (
            .O(N__6526),
            .I(N__6523));
    InMux I__588 (
            .O(N__6523),
            .I(N__6520));
    LocalMux I__587 (
            .O(N__6520),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO));
    InMux I__586 (
            .O(N__6517),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3));
    InMux I__585 (
            .O(N__6514),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4));
    CascadeMux I__584 (
            .O(N__6511),
            .I(N__6508));
    InMux I__583 (
            .O(N__6508),
            .I(N__6502));
    InMux I__582 (
            .O(N__6507),
            .I(N__6502));
    LocalMux I__581 (
            .O(N__6502),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO));
    InMux I__580 (
            .O(N__6499),
            .I(N__6496));
    LocalMux I__579 (
            .O(N__6496),
            .I(charx_i_24));
    InMux I__578 (
            .O(N__6493),
            .I(N__6490));
    LocalMux I__577 (
            .O(N__6490),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3));
    InMux I__576 (
            .O(N__6487),
            .I(N__6484));
    LocalMux I__575 (
            .O(N__6484),
            .I(charx_i_23));
    InMux I__574 (
            .O(N__6481),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__573 (
            .O(N__6478),
            .I(N__6475));
    LocalMux I__572 (
            .O(N__6475),
            .I(g1));
    InMux I__571 (
            .O(N__6472),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1));
    InMux I__570 (
            .O(N__6469),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2));
    InMux I__569 (
            .O(N__6466),
            .I(N__6463));
    LocalMux I__568 (
            .O(N__6463),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5));
    InMux I__567 (
            .O(N__6460),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4));
    CascadeMux I__566 (
            .O(N__6457),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_));
    CascadeMux I__565 (
            .O(N__6454),
            .I(N__6450));
    InMux I__564 (
            .O(N__6453),
            .I(N__6442));
    InMux I__563 (
            .O(N__6450),
            .I(N__6442));
    InMux I__562 (
            .O(N__6449),
            .I(N__6442));
    LocalMux I__561 (
            .O(N__6442),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803));
    CascadeMux I__560 (
            .O(N__6439),
            .I(font_un3_pixel_29_cascade_));
    CascadeMux I__559 (
            .O(N__6436),
            .I(Pixel_RNOZ0Z_18_cascade_));
    CascadeMux I__558 (
            .O(N__6433),
            .I(N_1214_0_cascade_));
    IoInMux I__557 (
            .O(N__6430),
            .I(N__6427));
    LocalMux I__556 (
            .O(N__6427),
            .I(N__6424));
    Span4Mux_s1_h I__555 (
            .O(N__6424),
            .I(N__6421));
    Span4Mux_h I__554 (
            .O(N__6421),
            .I(N__6418));
    Sp12to4 I__553 (
            .O(N__6418),
            .I(N__6415));
    Odrv12 I__552 (
            .O(N__6415),
            .I(\Clock50MHz.PixelClock ));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_9_8_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__6430),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam beamX_RNII5M_9_LC_1_2_3.C_ON=1'b0;
    defparam beamX_RNII5M_9_LC_1_2_3.SEQ_MODE=4'b0000;
    defparam beamX_RNII5M_9_LC_1_2_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNII5M_9_LC_1_2_3 (
            .in0(N__7259),
            .in1(N__8434),
            .in2(N__7528),
            .in3(N__7211),
            .lcout(un18_beamylto9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_0_LC_1_3_1.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_0_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_0_LC_1_3_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_0_LC_1_3_1 (
            .in0(N__7821),
            .in1(N__9296),
            .in2(_gnd_net_),
            .in3(N__7737),
            .lcout(font_un3_pixel_29),
            .ltout(font_un3_pixel_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_18_LC_1_3_2.C_ON=1'b0;
    defparam Pixel_RNO_18_LC_1_3_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_18_LC_1_3_2.LUT_INIT=16'b1111001100000011;
    LogicCell40 Pixel_RNO_18_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(N__9513),
            .in2(N__6439),
            .in3(N__9529),
            .lcout(),
            .ltout(Pixel_RNOZ0Z_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_5_LC_1_3_3.C_ON=1'b0;
    defparam Pixel_RNO_5_LC_1_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_5_LC_1_3_3.LUT_INIT=16'b1111000111100000;
    LogicCell40 Pixel_RNO_5_LC_1_3_3 (
            .in0(N__13108),
            .in1(N__6478),
            .in2(N__6436),
            .in3(N__8998),
            .lcout(),
            .ltout(N_1214_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_0_LC_1_3_4.C_ON=1'b0;
    defparam Pixel_RNO_0_LC_1_3_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_0_LC_1_3_4.LUT_INIT=16'b1111111110101110;
    LogicCell40 Pixel_RNO_0_LC_1_3_4 (
            .in0(N__6826),
            .in1(N__6757),
            .in2(N__6433),
            .in3(N__6883),
            .lcout(G_21_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_20_LC_1_3_6.C_ON=1'b0;
    defparam Pixel_RNO_20_LC_1_3_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_20_LC_1_3_6.LUT_INIT=16'b0000111110100101;
    LogicCell40 Pixel_RNO_20_LC_1_3_6 (
            .in0(N__7738),
            .in1(_gnd_net_),
            .in2(N__9315),
            .in3(N__7822),
            .lcout(g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_1_4_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_1_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7825),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_1_4_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_1_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_1_4_1 (
            .in0(_gnd_net_),
            .in1(N__6487),
            .in2(N__6511),
            .in3(N__6472),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_71_LC_1_4_2.C_ON=1'b1;
    defparam Pixel_RNO_71_LC_1_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_71_LC_1_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_71_LC_1_4_2 (
            .in0(_gnd_net_),
            .in1(N__6547),
            .in2(N__6454),
            .in3(N__6469),
            .lcout(Pixel_RNOZ0Z_71),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_1_4_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_1_4_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_1_4_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_1_4_3 (
            .in0(_gnd_net_),
            .in1(N__6466),
            .in2(N__6538),
            .in3(N__6449),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_1_4_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_1_4_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_1_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_1_4_4 (
            .in0(N__6453),
            .in1(N__6877),
            .in2(N__6526),
            .in3(N__6460),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3),
            .ltout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_30_LC_1_4_5.C_ON=1'b0;
    defparam Pixel_RNO_30_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_30_LC_1_4_5.LUT_INIT=16'b0011000000000000;
    LogicCell40 Pixel_RNO_30_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(N__7808),
            .in2(N__6457),
            .in3(N__7939),
            .lcout(g0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_1_4_6.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_1_4_6.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_1_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_1_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6507),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_1_5_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_1_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_1_5_0 (
            .in0(_gnd_net_),
            .in1(N__7015),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_1_5_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_1_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__6499),
            .in2(_gnd_net_),
            .in3(N__6541),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDB3_LC_1_5_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDB3_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDB3_LC_1_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDB3_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(N__6493),
            .in2(N__15585),
            .in3(N__6529),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_1_5_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_1_5_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_1_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_1_5_3 (
            .in0(_gnd_net_),
            .in1(N__6876),
            .in2(_gnd_net_),
            .in3(N__6517),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_1_5_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_1_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_1_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6514),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_1_5_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_1_5_5.LUT_INIT=16'b1100011000110011;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_1_5_5 (
            .in0(N__7003),
            .in1(N__6974),
            .in2(N__10342),
            .in3(N__6937),
            .lcout(charx_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_1_5_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_1_5_6.LUT_INIT=16'b1000101001110101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_1_5_6 (
            .in0(N__6938),
            .in1(N__10330),
            .in2(N__7009),
            .in3(N__6975),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_1_5_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_1_5_7.LUT_INIT=16'b0011110000110011;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_1_5_7 (
            .in0(_gnd_net_),
            .in1(N__7007),
            .in2(N__10343),
            .in3(N__6939),
            .lcout(charx_i_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_1_6_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_1_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(N__9997),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_1_6_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_1_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(N__6679),
            .in2(N__6589),
            .in3(N__6481),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_1_6_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_1_6_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_1_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_1_6_2 (
            .in0(_gnd_net_),
            .in1(N__6700),
            .in2(N__6580),
            .in3(N__6613),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_1_6_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_1_6_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_1_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_1_6_3 (
            .in0(_gnd_net_),
            .in1(N__6610),
            .in2(N__6568),
            .in3(N__6698),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_1_6_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_1_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_1_6_4 (
            .in0(_gnd_net_),
            .in1(N__6556),
            .in2(_gnd_net_),
            .in3(N__6604),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_4_LC_1_6_5.C_ON=1'b0;
    defparam beamX_RNIVEM1_4_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_4_LC_1_6_5.LUT_INIT=16'b1101000011000000;
    LogicCell40 beamX_RNIVEM1_4_LC_1_6_5 (
            .in0(N__7391),
            .in1(N__7321),
            .in2(N__6601),
            .in3(N__7584),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_2_LC_1_6_6.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_2_LC_1_6_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_2_LC_1_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_2_LC_1_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9841),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_1_7_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_1_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_1_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_1_7_0 (
            .in0(_gnd_net_),
            .in1(N__9840),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_1_7_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_1_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_1_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_1_7_1 (
            .in0(_gnd_net_),
            .in1(N__6672),
            .in2(N__6718),
            .in3(N__6571),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_1_7_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_1_7_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_1_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_1_7_2 (
            .in0(_gnd_net_),
            .in1(N__6627),
            .in2(N__6664),
            .in3(N__6559),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_1_7_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_1_7_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_1_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_1_7_3 (
            .in0(N__6699),
            .in1(N__6673),
            .in2(N__6652),
            .in3(N__6550),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_1_7_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_1_7_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_1_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_1_7_4 (
            .in0(_gnd_net_),
            .in1(N__6640),
            .in2(_gnd_net_),
            .in3(N__6703),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0),
            .ltout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_1_7_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_1_7_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_1_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_1_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6682),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_1_7_6.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_1_7_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_1_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_1_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6626),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_1_8_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_1_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(N__8704),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_1_8_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_1_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_1_8_1 (
            .in0(_gnd_net_),
            .in1(N__7167),
            .in2(N__6727),
            .in3(N__6655),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_1_8_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_1_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(N__8248),
            .in2(N__8293),
            .in3(N__6643),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_1_8_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_1_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_1_8_3 (
            .in0(N__6628),
            .in1(N__7168),
            .in2(N__8278),
            .in3(N__6634),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_1_8_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_1_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_1_8_4 (
            .in0(_gnd_net_),
            .in1(N__8263),
            .in2(_gnd_net_),
            .in3(N__6631),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_1_8_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_1_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_1_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8977),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_1_8_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_1_8_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_1_8_7 (
            .in0(N__8705),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_1_9_2.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_1_9_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 beamX_RNI5457_5_LC_1_9_2 (
            .in0(N__8465),
            .in1(N__7468),
            .in2(N__8420),
            .in3(N__7314),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_ofx_LC_1_10_1.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_ofx_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_ofx_LC_1_10_1.LUT_INIT=16'b0100101010110101;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_3_l_ofx_LC_1_10_1 (
            .in0(N__8961),
            .in1(N__8906),
            .in2(N__9133),
            .in3(N__8684),
            .lcout(if_generate_plus_mult1_un54_sum_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_ofx_LC_1_10_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_ofx_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_ofx_LC_1_10_4.LUT_INIT=16'b0010110110111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_l_ofx_LC_1_10_4 (
            .in0(N__9126),
            .in1(N__8691),
            .in2(N__8911),
            .in3(N__8963),
            .lcout(if_generate_plus_mult1_un54_sum_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_i_LC_1_10_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_i_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_i_LC_1_10_5.LUT_INIT=16'b0110001111100111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_c5_i_LC_1_10_5 (
            .in0(N__8962),
            .in1(N__8907),
            .in2(N__9134),
            .in3(N__8685),
            .lcout(column_1_if_generate_plus_mult1_un47_sum_c5_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_1_10_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_1_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8683),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_1_11_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_1_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_1_11_0 (
            .in0(_gnd_net_),
            .in1(N__7893),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_1_11_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_1_11_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(N__7365),
            .in2(_gnd_net_),
            .in3(N__6709),
            .lcout(charx_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_1_11_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_1_11_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_1_11_2 (
            .in0(_gnd_net_),
            .in1(N__7456),
            .in2(_gnd_net_),
            .in3(N__6706),
            .lcout(charx_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_1_11_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_1_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_1_11_3 (
            .in0(_gnd_net_),
            .in1(N__7425),
            .in2(N__15586),
            .in3(N__6751),
            .lcout(chessboardpixel_un152_pixel_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_1_11_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_1_11_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_1_11_4 (
            .in0(_gnd_net_),
            .in1(N__7558),
            .in2(_gnd_net_),
            .in3(N__6748),
            .lcout(charx_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_1_11_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_1_11_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_1_11_5 (
            .in0(_gnd_net_),
            .in1(N__7300),
            .in2(_gnd_net_),
            .in3(N__6745),
            .lcout(charx_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_1_11_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_1_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_1_11_6 (
            .in0(_gnd_net_),
            .in1(N__7501),
            .in2(N__15587),
            .in3(N__6742),
            .lcout(charx_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_1_11_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_1_11_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_1_11_7 (
            .in0(_gnd_net_),
            .in1(N__8390),
            .in2(_gnd_net_),
            .in3(N__6739),
            .lcout(charx_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_1_12_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_1_12_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_1_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_1_12_0 (
            .in0(_gnd_net_),
            .in1(N__7238),
            .in2(N__15596),
            .in3(N__6736),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_1_12_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_1_12_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_1_12_1 (
            .in0(_gnd_net_),
            .in1(N__7189),
            .in2(_gnd_net_),
            .in3(N__6733),
            .lcout(charx_if_generate_plus_mult1_un26_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_1_13_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_1_13_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_1_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_1_13_0 (
            .in0(_gnd_net_),
            .in1(N__8878),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_1_13_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_1_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_1_13_1 (
            .in0(_gnd_net_),
            .in1(N__6769),
            .in2(_gnd_net_),
            .in3(N__6730),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_1_13_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_1_13_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_1_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_1_13_2 (
            .in0(_gnd_net_),
            .in1(N__6775),
            .in2(N__15597),
            .in3(N__6784),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_1_13_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_1_13_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_1_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_1_13_3 (
            .in0(_gnd_net_),
            .in1(N__9100),
            .in2(_gnd_net_),
            .in3(N__6781),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_1_13_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_1_13_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_1_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_1_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6778),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_1_13_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_1_13_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_1_13_6 (
            .in0(N__9099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_1_13_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_1_13_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_1_13_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_2_LC_1_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9098),
            .lcout(charx_if_generate_plus_mult1_un26_sum_axb_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_48_LC_2_2_2.C_ON=1'b0;
    defparam Pixel_RNO_48_LC_2_2_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_48_LC_2_2_2.LUT_INIT=16'b1110111011111110;
    LogicCell40 Pixel_RNO_48_LC_2_2_2 (
            .in0(N__7212),
            .in1(N__7260),
            .in2(N__8440),
            .in3(N__8143),
            .lcout(),
            .ltout(g1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_26_LC_2_2_3.C_ON=1'b0;
    defparam Pixel_RNO_26_LC_2_2_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_26_LC_2_2_3.LUT_INIT=16'b1101111111111111;
    LogicCell40 Pixel_RNO_26_LC_2_2_3 (
            .in0(N__8101),
            .in1(N__8338),
            .in2(N__6763),
            .in3(N__8191),
            .lcout(),
            .ltout(g2_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_7_LC_2_2_4.C_ON=1'b0;
    defparam Pixel_RNO_7_LC_2_2_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_7_LC_2_2_4.LUT_INIT=16'b0000000011000000;
    LogicCell40 Pixel_RNO_7_LC_2_2_4 (
            .in0(_gnd_net_),
            .in1(N__6790),
            .in2(N__6760),
            .in3(N__7962),
            .lcout(g2_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_73_LC_2_2_6.C_ON=1'b0;
    defparam Pixel_RNO_73_LC_2_2_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_73_LC_2_2_6.LUT_INIT=16'b1101110111011101;
    LogicCell40 Pixel_RNO_73_LC_2_2_6 (
            .in0(N__8435),
            .in1(N__8142),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(g3_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_56_LC_2_2_7.C_ON=1'b0;
    defparam Pixel_RNO_56_LC_2_2_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_56_LC_2_2_7.LUT_INIT=16'b1100110010001100;
    LogicCell40 Pixel_RNO_56_LC_2_2_7 (
            .in0(N__7261),
            .in1(N__8100),
            .in2(N__6835),
            .in3(N__7213),
            .lcout(g0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_38_LC_2_3_0.C_ON=1'b0;
    defparam Pixel_RNO_38_LC_2_3_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_38_LC_2_3_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 Pixel_RNO_38_LC_2_3_0 (
            .in0(N__7813),
            .in1(N__7961),
            .in2(_gnd_net_),
            .in3(N__7739),
            .lcout(),
            .ltout(g0_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_17_LC_2_3_1.C_ON=1'b0;
    defparam Pixel_RNO_17_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_17_LC_2_3_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 Pixel_RNO_17_LC_2_3_1 (
            .in0(N__6892),
            .in1(N__8155),
            .in2(N__6832),
            .in3(N__6820),
            .lcout(),
            .ltout(g0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_4_LC_2_3_2.C_ON=1'b0;
    defparam Pixel_RNO_4_LC_2_3_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_4_LC_2_3_2.LUT_INIT=16'b0001000000110000;
    LogicCell40 Pixel_RNO_4_LC_2_3_2 (
            .in0(N__6901),
            .in1(N__9016),
            .in2(N__6829),
            .in3(N__9007),
            .lcout(N_21_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_37_LC_2_3_3.C_ON=1'b0;
    defparam Pixel_RNO_37_LC_2_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_37_LC_2_3_3.LUT_INIT=16'b0000000010111010;
    LogicCell40 Pixel_RNO_37_LC_2_3_3 (
            .in0(N__9295),
            .in1(N__13106),
            .in2(N__13294),
            .in3(N__9512),
            .lcout(Pixel_RNOZ0Z_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_72_LC_2_3_4.C_ON=1'b0;
    defparam Pixel_RNO_72_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_72_LC_2_3_4.LUT_INIT=16'b0001000111101110;
    LogicCell40 Pixel_RNO_72_LC_2_3_4 (
            .in0(N__7812),
            .in1(N__9294),
            .in2(_gnd_net_),
            .in3(N__7960),
            .lcout(),
            .ltout(font_un126_pixel_m_2_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_55_LC_2_3_5.C_ON=1'b0;
    defparam Pixel_RNO_55_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_55_LC_2_3_5.LUT_INIT=16'b0110000000000110;
    LogicCell40 Pixel_RNO_55_LC_2_3_5 (
            .in0(N__7740),
            .in1(N__7814),
            .in2(N__6814),
            .in3(N__6811),
            .lcout(),
            .ltout(font_un126_pixel_m_2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_33_LC_2_3_6.C_ON=1'b0;
    defparam Pixel_RNO_33_LC_2_3_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_33_LC_2_3_6.LUT_INIT=16'b1000101000000000;
    LogicCell40 Pixel_RNO_33_LC_2_3_6 (
            .in0(N__6805),
            .in1(N__6799),
            .in2(N__6793),
            .in3(N__8334),
            .lcout(g0_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_25_LC_2_3_7.C_ON=1'b0;
    defparam Pixel_RNO_25_LC_2_3_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_25_LC_2_3_7.LUT_INIT=16'b0110010001100010;
    LogicCell40 Pixel_RNO_25_LC_2_3_7 (
            .in0(N__7741),
            .in1(N__7815),
            .in2(N__12952),
            .in3(N__9308),
            .lcout(g2_2_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_2_4_0.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_2_4_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_2_4_0.LUT_INIT=16'b1100110000110011;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_2_4_0 (
            .in0(_gnd_net_),
            .in1(N__10341),
            .in2(_gnd_net_),
            .in3(N__6943),
            .lcout(charx_if_generate_plus_mult1_un1_sum_axb1),
            .ltout(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_16_LC_2_4_1.C_ON=1'b0;
    defparam Pixel_RNO_16_LC_2_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_16_LC_2_4_1.LUT_INIT=16'b0000001000110001;
    LogicCell40 Pixel_RNO_16_LC_2_4_1 (
            .in0(N__7745),
            .in1(N__9199),
            .in2(N__6904),
            .in3(N__9305),
            .lcout(font_un126_pixel_5_a0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_8_LC_2_4_2.C_ON=1'b0;
    defparam Pixel_RNO_8_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_8_LC_2_4_2.LUT_INIT=16'b0000000010001000;
    LogicCell40 Pixel_RNO_8_LC_2_4_2 (
            .in0(N__7948),
            .in1(N__7824),
            .in2(_gnd_net_),
            .in3(N__7747),
            .lcout(),
            .ltout(G_19_i_a11_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_1_LC_2_4_3.C_ON=1'b0;
    defparam Pixel_RNO_1_LC_2_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_1_LC_2_4_3.LUT_INIT=16'b0100000001110000;
    LogicCell40 Pixel_RNO_1_LC_2_4_3 (
            .in0(N__9337),
            .in1(N__9307),
            .in2(N__6895),
            .in3(N__9208),
            .lcout(N_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_36_LC_2_4_4.C_ON=1'b0;
    defparam Pixel_RNO_36_LC_2_4_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_36_LC_2_4_4.LUT_INIT=16'b0000000010001000;
    LogicCell40 Pixel_RNO_36_LC_2_4_4 (
            .in0(N__9198),
            .in1(N__13107),
            .in2(_gnd_net_),
            .in3(N__13287),
            .lcout(Pixel_RNOZ0Z_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_24_LC_2_4_6.C_ON=1'b0;
    defparam Pixel_RNO_24_LC_2_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_24_LC_2_4_6.LUT_INIT=16'b0010000001000000;
    LogicCell40 Pixel_RNO_24_LC_2_4_6 (
            .in0(N__9306),
            .in1(N__7823),
            .in2(N__7861),
            .in3(N__7746),
            .lcout(),
            .ltout(g1_1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_6_LC_2_4_7.C_ON=1'b0;
    defparam Pixel_RNO_6_LC_2_4_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_6_LC_2_4_7.LUT_INIT=16'b1111100010001000;
    LogicCell40 Pixel_RNO_6_LC_2_4_7 (
            .in0(N__9367),
            .in1(N__9544),
            .in2(N__6886),
            .in3(N__8071),
            .lcout(g0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_2_5_0.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_2_5_0.LUT_INIT=16'b0011100111001100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_2_5_0 (
            .in0(N__7008),
            .in1(N__6976),
            .in2(N__10345),
            .in3(N__6936),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIL5OEN1_LC_2_5_1.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIL5OEN1_LC_2_5_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIL5OEN1_LC_2_5_1.LUT_INIT=16'b0110001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIL5OEN1_LC_2_5_1 (
            .in0(N__10005),
            .in1(N__6865),
            .in2(N__6858),
            .in3(N__6843),
            .lcout(chessboardpixel_un152_pixel_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAKPE41_LC_2_5_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAKPE41_LC_2_5_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAKPE41_LC_2_5_5.LUT_INIT=16'b1010010011010000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAKPE41_LC_2_5_5 (
            .in0(N__10006),
            .in1(N__10592),
            .in2(N__6859),
            .in3(N__6844),
            .lcout(chessboardpixel_un174_pixellt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_2_5_6.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_2_5_6.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_2_5_6 (
            .in0(N__10337),
            .in1(N__7002),
            .in2(_gnd_net_),
            .in3(N__6935),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI8P51_4_LC_2_5_7.C_ON=1'b0;
    defparam beamX_RNI8P51_4_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam beamX_RNI8P51_4_LC_2_5_7.LUT_INIT=16'b0101000101010101;
    LogicCell40 beamX_RNI8P51_4_LC_2_5_7 (
            .in0(N__7522),
            .in1(N__7319),
            .in2(N__7398),
            .in3(N__7582),
            .lcout(un13_beamylt7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_2_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_2_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_2_6_0 (
            .in0(_gnd_net_),
            .in1(N__10326),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_2_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_2_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_2_6_1 (
            .in0(_gnd_net_),
            .in1(N__6954),
            .in2(N__6913),
            .in3(N__6979),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_2_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_2_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_2_6_2 (
            .in0(_gnd_net_),
            .in1(N__7087),
            .in2(N__7045),
            .in3(N__6958),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_2_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_2_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_2_6_3 (
            .in0(_gnd_net_),
            .in1(N__6955),
            .in2(N__7075),
            .in3(N__7041),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_2_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_2_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_2_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_2_6_4 (
            .in0(_gnd_net_),
            .in1(N__7060),
            .in2(_gnd_net_),
            .in3(N__6946),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_RNO_0_LC_2_6_5.C_ON=1'b0;
    defparam HSync_RNO_0_LC_2_6_5.SEQ_MODE=4'b0000;
    defparam HSync_RNO_0_LC_2_6_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 HSync_RNO_0_LC_2_6_5 (
            .in0(N__7320),
            .in1(N__7438),
            .in2(N__7588),
            .in3(N__7524),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_2_7_0.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_2_7_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_2_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10223),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_2_7_2.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_2_7_2.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_RNIR4B_9_LC_2_7_2 (
            .in0(N__7257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7209),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_77_LC_2_7_6.C_ON=1'b0;
    defparam Pixel_RNO_77_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_77_LC_2_7_6.LUT_INIT=16'b0101000101010101;
    LogicCell40 Pixel_RNO_77_LC_2_7_6 (
            .in0(N__7523),
            .in1(N__7318),
            .in2(N__7399),
            .in3(N__7578),
            .lcout(),
            .ltout(un13_beamylt7_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_61_LC_2_7_7.C_ON=1'b0;
    defparam Pixel_RNO_61_LC_2_7_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_61_LC_2_7_7.LUT_INIT=16'b1110111111101110;
    LogicCell40 Pixel_RNO_61_LC_2_7_7 (
            .in0(N__7210),
            .in1(N__7258),
            .in2(N__7090),
            .in3(N__8429),
            .lcout(g1_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_2_8_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_2_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(N__10214),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_2_8_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_2_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(N__7107),
            .in2(N__7024),
            .in3(N__7078),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_2_8_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_2_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(N__7123),
            .in2(N__7159),
            .in3(N__7063),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_2_8_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_2_8_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_2_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_2_8_3 (
            .in0(N__7040),
            .in1(N__7108),
            .in2(N__7147),
            .in3(N__7051),
            .lcout(charx_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_2_8_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_2_8_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_2_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_2_8_4 (
            .in0(_gnd_net_),
            .in1(N__7135),
            .in2(_gnd_net_),
            .in3(N__7048),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_2_8_5.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_2_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_2_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10585),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_2_8_6.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_2_8_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_2_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_2_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8243),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_2_9_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_2_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_2_9_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_2_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__8541),
            .in2(N__7099),
            .in3(N__7150),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_2_9_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_2_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_2_9_2 (
            .in0(_gnd_net_),
            .in1(N__9586),
            .in2(N__9631),
            .in3(N__7138),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_2_9_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_2_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_2_9_3 (
            .in0(N__7122),
            .in1(N__8542),
            .in2(N__9616),
            .in3(N__7129),
            .lcout(charx_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_2_9_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_2_9_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_2_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_2_9_4 (
            .in0(_gnd_net_),
            .in1(N__9601),
            .in2(_gnd_net_),
            .in3(N__7126),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0),
            .ltout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_2_9_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_2_9_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_2_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7111),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_2_9_7.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_2_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_2_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10004),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_2_10_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_2_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(N__7369),
            .in2(N__7930),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_2_10_1.C_ON=1'b1;
    defparam beamX_2_LC_2_10_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_2_10_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(N__7459),
            .in2(_gnd_net_),
            .in3(N__7330),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_2_10_2.C_ON=1'b1;
    defparam beamX_3_LC_2_10_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_2_10_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(N__7435),
            .in2(_gnd_net_),
            .in3(N__7327),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_2_10_3.C_ON=1'b1;
    defparam beamX_4_LC_2_10_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_2_10_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_2_10_3 (
            .in0(N__13360),
            .in1(N__7574),
            .in2(_gnd_net_),
            .in3(N__7324),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_2_10_4.C_ON=1'b1;
    defparam beamX_5_LC_2_10_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_2_10_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__7313),
            .in2(_gnd_net_),
            .in3(N__7270),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_2_10_5.C_ON=1'b1;
    defparam beamX_6_LC_2_10_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_2_10_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(N__7521),
            .in2(_gnd_net_),
            .in3(N__7267),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_2_10_6.C_ON=1'b1;
    defparam beamX_7_LC_2_10_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_2_10_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_2_10_6 (
            .in0(_gnd_net_),
            .in1(N__8405),
            .in2(_gnd_net_),
            .in3(N__7264),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_2_10_7.C_ON=1'b1;
    defparam beamX_8_LC_2_10_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_2_10_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_2_10_7 (
            .in0(_gnd_net_),
            .in1(N__7237),
            .in2(_gnd_net_),
            .in3(N__7216),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__13418),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_2_11_0.C_ON=1'b1;
    defparam beamX_9_LC_2_11_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_2_11_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_2_11_0 (
            .in0(_gnd_net_),
            .in1(N__7200),
            .in2(_gnd_net_),
            .in3(N__7171),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__13419),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_2_11_1.C_ON=1'b0;
    defparam beamX_10_LC_2_11_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_2_11_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_10_LC_2_11_1 (
            .in0(N__13373),
            .in1(N__8487),
            .in2(_gnd_net_),
            .in3(N__7591),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_10_LC_2_11_3.C_ON=1'b0;
    defparam beamX_RNICPU5_10_LC_2_11_3.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_10_LC_2_11_3.LUT_INIT=16'b0001000000000000;
    LogicCell40 beamX_RNICPU5_10_LC_2_11_3 (
            .in0(N__7367),
            .in1(N__7458),
            .in2(N__7583),
            .in3(N__8486),
            .lcout(un3_beamx_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_2_11_4.C_ON=1'b0;
    defparam beamX_0_LC_2_11_4.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_2_11_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_0_LC_2_11_4 (
            .in0(_gnd_net_),
            .in1(N__13374),
            .in2(_gnd_net_),
            .in3(N__7899),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_3_LC_2_11_5.C_ON=1'b0;
    defparam beamX_RNIKVE6_3_LC_2_11_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_3_LC_2_11_5.LUT_INIT=16'b0000000100000000;
    LogicCell40 beamX_RNIKVE6_3_LC_2_11_5 (
            .in0(N__7895),
            .in1(N__7517),
            .in2(N__7437),
            .in3(N__7474),
            .lcout(un3_beamx_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_2_11_6.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_2_11_6.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_2_11_6.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamX_RNIQCL_1_LC_2_11_6 (
            .in0(N__7457),
            .in1(N__7366),
            .in2(N__7436),
            .in3(N__7894),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_2_11_7.C_ON=1'b0;
    defparam beamX_1_LC_2_11_7.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_2_11_7.LUT_INIT=16'b1010010101011010;
    LogicCell40 beamX_1_LC_2_11_7 (
            .in0(N__7368),
            .in1(_gnd_net_),
            .in2(N__7913),
            .in3(_gnd_net_),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_LC_2_12_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_LC_2_12_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_LC_2_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_1_c_LC_2_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_2_12_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_2_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(N__7621),
            .in2(N__7636),
            .in3(N__7345),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_2_12_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_2_12_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_2_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_2_12_2 (
            .in0(_gnd_net_),
            .in1(N__7611),
            .in2(N__7342),
            .in3(N__7333),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_2_12_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_2_12_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_2_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_2_12_3 (
            .in0(N__9164),
            .in1(N__7627),
            .in2(N__7657),
            .in3(N__7648),
            .lcout(charx_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_2_12_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_2_12_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_2_12_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_2_12_4 (
            .in0(N__7645),
            .in1(N__7612),
            .in2(N__9119),
            .in3(N__7639),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_2_12_5.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_2_12_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_2_12_5.LUT_INIT=16'b0011001100110011;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_2_12_5 (
            .in0(_gnd_net_),
            .in1(N__8879),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_2_12_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_2_12_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_2_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_2_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7610),
            .lcout(charx_if_generate_plus_mult1_un26_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_2_12_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_2_12_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_2_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_2_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7620),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_2_13_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_2_13_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_2_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_2_13_0 (
            .in0(_gnd_net_),
            .in1(N__9104),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_2_13_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_2_13_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_2_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_2_13_1 (
            .in0(_gnd_net_),
            .in1(N__15602),
            .in2(_gnd_net_),
            .in3(N__7600),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_2_13_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_2_13_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_2_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_2_13_2 (
            .in0(_gnd_net_),
            .in1(N__15606),
            .in2(N__15607),
            .in3(N__7597),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_13_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_13_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7594),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_2_13_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_2_13_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_2_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_2_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7681),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_4_2_0.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_4_2_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_4_2_0.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_4_2_0 (
            .in0(N__7837),
            .in1(N__9319),
            .in2(_gnd_net_),
            .in3(N__7757),
            .lcout(g2_1),
            .ltout(g2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_74_LC_4_2_1.C_ON=1'b0;
    defparam Pixel_RNO_74_LC_4_2_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_74_LC_4_2_1.LUT_INIT=16'b1100111100001100;
    LogicCell40 Pixel_RNO_74_LC_4_2_1 (
            .in0(_gnd_net_),
            .in1(N__13109),
            .in2(N__7678),
            .in3(N__13289),
            .lcout(),
            .ltout(N_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_58_LC_4_2_2.C_ON=1'b0;
    defparam Pixel_RNO_58_LC_4_2_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_58_LC_4_2_2.LUT_INIT=16'b1000000001000000;
    LogicCell40 Pixel_RNO_58_LC_4_2_2 (
            .in0(N__7838),
            .in1(N__7965),
            .in2(N__7675),
            .in3(N__7758),
            .lcout(g1_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_76_LC_4_2_4.C_ON=1'b0;
    defparam Pixel_RNO_76_LC_4_2_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_76_LC_4_2_4.LUT_INIT=16'b0101101000000000;
    LogicCell40 Pixel_RNO_76_LC_4_2_4 (
            .in0(N__13290),
            .in1(_gnd_net_),
            .in2(N__13114),
            .in3(N__7964),
            .lcout(),
            .ltout(g0_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_60_LC_4_2_5.C_ON=1'b0;
    defparam Pixel_RNO_60_LC_4_2_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_60_LC_4_2_5.LUT_INIT=16'b0000000010000000;
    LogicCell40 Pixel_RNO_60_LC_4_2_5 (
            .in0(N__7672),
            .in1(N__7989),
            .in2(N__7666),
            .in3(N__9511),
            .lcout(),
            .ltout(g0_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_35_LC_4_2_6.C_ON=1'b0;
    defparam Pixel_RNO_35_LC_4_2_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_35_LC_4_2_6.LUT_INIT=16'b0001000000100000;
    LogicCell40 Pixel_RNO_35_LC_4_2_6 (
            .in0(N__12911),
            .in1(N__9922),
            .in2(N__7663),
            .in3(N__9909),
            .lcout(g3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_13_LC_4_3_0.C_ON=1'b0;
    defparam Pixel_RNO_13_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_13_LC_4_3_0.LUT_INIT=16'b1111110111111111;
    LogicCell40 Pixel_RNO_13_LC_4_3_0 (
            .in0(N__7966),
            .in1(N__13113),
            .in2(N__13296),
            .in3(N__7990),
            .lcout(),
            .ltout(g3_2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_3_LC_4_3_1.C_ON=1'b0;
    defparam Pixel_RNO_3_LC_4_3_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_3_LC_4_3_1.LUT_INIT=16'b0101010000000000;
    LogicCell40 Pixel_RNO_3_LC_4_3_1 (
            .in0(N__9244),
            .in1(N__8218),
            .in2(N__7660),
            .in3(N__7996),
            .lcout(),
            .ltout(g0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_4_3_2.C_ON=1'b0;
    defparam PixelZ0_LC_4_3_2.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_4_3_2.LUT_INIT=16'b0000000010111010;
    LogicCell40 PixelZ0_LC_4_3_2 (
            .in0(N__7849),
            .in1(N__8059),
            .in2(N__8047),
            .in3(N__8044),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_34_LC_4_3_3.C_ON=1'b0;
    defparam Pixel_RNO_34_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_34_LC_4_3_3.LUT_INIT=16'b0000010010001000;
    LogicCell40 Pixel_RNO_34_LC_4_3_3 (
            .in0(N__7690),
            .in1(N__8020),
            .in2(N__7978),
            .in3(N__9514),
            .lcout(),
            .ltout(g1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_12_LC_4_3_4.C_ON=1'b0;
    defparam Pixel_RNO_12_LC_4_3_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_12_LC_4_3_4.LUT_INIT=16'b0000000000001000;
    LogicCell40 Pixel_RNO_12_LC_4_3_4 (
            .in0(N__9217),
            .in1(N__8014),
            .in2(N__8005),
            .in3(N__8002),
            .lcout(g0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI50PU65_LC_4_3_5.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI50PU65_LC_4_3_5.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI50PU65_LC_4_3_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI50PU65_LC_4_3_5 (
            .in0(_gnd_net_),
            .in1(N__7839),
            .in2(_gnd_net_),
            .in3(N__7759),
            .lcout(g1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_57_LC_4_4_0.C_ON=1'b0;
    defparam Pixel_RNO_57_LC_4_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_57_LC_4_4_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 Pixel_RNO_57_LC_4_4_0 (
            .in0(N__13267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13090),
            .lcout(g0_0_a3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_46_LC_4_4_1.C_ON=1'b0;
    defparam Pixel_RNO_46_LC_4_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_46_LC_4_4_1.LUT_INIT=16'b0000101100001111;
    LogicCell40 Pixel_RNO_46_LC_4_4_1 (
            .in0(N__8326),
            .in1(N__8183),
            .in2(N__7963),
            .in3(N__8121),
            .lcout(N_35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_2_LC_4_4_2.C_ON=1'b0;
    defparam Pixel_RNO_2_LC_4_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_2_LC_4_4_2.LUT_INIT=16'b0000000010001000;
    LogicCell40 Pixel_RNO_2_LC_4_4_2 (
            .in0(N__8184),
            .in1(N__8122),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(N_58_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDQG2_0_LC_4_4_4.C_ON=1'b0;
    defparam beamY_RNIDQG2_0_LC_4_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIDQG2_0_LC_4_4_4.LUT_INIT=16'b0101010110101010;
    LogicCell40 beamY_RNIDQG2_0_LC_4_4_4 (
            .in0(N__13266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13089),
            .lcout(),
            .ltout(beamY_RNIDQG2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNINKIU27_0_LC_4_4_5.C_ON=1'b0;
    defparam beamY_RNINKIU27_0_LC_4_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNINKIU27_0_LC_4_4_5.LUT_INIT=16'b0000100100001100;
    LogicCell40 beamY_RNINKIU27_0_LC_4_4_5 (
            .in0(N__7840),
            .in1(N__9316),
            .in2(N__7762),
            .in3(N__7756),
            .lcout(beamY_RNINKIU27Z0Z_0),
            .ltout(beamY_RNINKIU27Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_29_LC_4_4_6.C_ON=1'b0;
    defparam Pixel_RNO_29_LC_4_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_29_LC_4_4_6.LUT_INIT=16'b1010010110101101;
    LogicCell40 Pixel_RNO_29_LC_4_4_6 (
            .in0(N__9508),
            .in1(N__13091),
            .in2(N__8224),
            .in3(N__13297),
            .lcout(),
            .ltout(Pixel_RNOZ0Z_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_10_LC_4_4_7.C_ON=1'b0;
    defparam Pixel_RNO_10_LC_4_4_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_10_LC_4_4_7.LUT_INIT=16'b1111110010111000;
    LogicCell40 Pixel_RNO_10_LC_4_4_7 (
            .in0(N__9231),
            .in1(N__9317),
            .in2(N__8221),
            .in3(N__9509),
            .lcout(N_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGH4H57_1_LC_4_5_0.C_ON=1'b0;
    defparam beamY_RNIGH4H57_1_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIGH4H57_1_LC_4_5_0.LUT_INIT=16'b0000010100110110;
    LogicCell40 beamY_RNIGH4H57_1_LC_4_5_0 (
            .in0(N__8212),
            .in1(N__10939),
            .in2(N__8203),
            .in3(N__10852),
            .lcout(chessboardpixel_un175_pixel),
            .ltout(chessboardpixel_un175_pixel_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_39_LC_4_5_1.C_ON=1'b0;
    defparam Pixel_RNO_39_LC_4_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_39_LC_4_5_1.LUT_INIT=16'b1111111101111111;
    LogicCell40 Pixel_RNO_39_LC_4_5_1 (
            .in0(N__8170),
            .in1(N__8088),
            .in2(N__8158),
            .in3(N__8325),
            .lcout(g2_3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNISO4T_7_LC_4_5_3.C_ON=1'b0;
    defparam beamX_RNISO4T_7_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam beamX_RNISO4T_7_LC_4_5_3.LUT_INIT=16'b0100110000001100;
    LogicCell40 beamX_RNISO4T_7_LC_4_5_3 (
            .in0(N__8141),
            .in1(N__8087),
            .in2(N__8470),
            .in3(N__8430),
            .lcout(un15_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIT9ER_10_LC_4_6_0.C_ON=1'b0;
    defparam beamX_RNIT9ER_10_LC_4_6_0.SEQ_MODE=4'b0000;
    defparam beamX_RNIT9ER_10_LC_4_6_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNIT9ER_10_LC_4_6_0 (
            .in0(N__8110),
            .in1(N__9352),
            .in2(N__8500),
            .in3(N__9412),
            .lcout(un15_beamy_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_44_LC_4_6_1.C_ON=1'b0;
    defparam Pixel_RNO_44_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_44_LC_4_6_1.LUT_INIT=16'b0000000000010100;
    LogicCell40 Pixel_RNO_44_LC_4_6_1 (
            .in0(N__9188),
            .in1(N__12910),
            .in2(N__9910),
            .in3(N__9467),
            .lcout(),
            .ltout(Pixel_RNOZ0Z_44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_21_LC_4_6_2.C_ON=1'b0;
    defparam Pixel_RNO_21_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_21_LC_4_6_2.LUT_INIT=16'b0000001001000110;
    LogicCell40 Pixel_RNO_21_LC_4_6_2 (
            .in0(N__13257),
            .in1(N__13093),
            .in2(N__8074),
            .in3(N__9346),
            .lcout(N_10_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_45_LC_4_6_4.C_ON=1'b0;
    defparam Pixel_RNO_45_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_45_LC_4_6_4.LUT_INIT=16'b0101111101011111;
    LogicCell40 Pixel_RNO_45_LC_4_6_4 (
            .in0(N__13256),
            .in1(_gnd_net_),
            .in2(N__12931),
            .in3(_gnd_net_),
            .lcout(g4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSyncZ0_LC_4_6_6.C_ON=1'b0;
    defparam HSyncZ0_LC_4_6_6.SEQ_MODE=4'b1000;
    defparam HSyncZ0_LC_4_6_6.LUT_INIT=16'b1111111111111011;
    LogicCell40 HSyncZ0_LC_4_6_6 (
            .in0(N__8499),
            .in1(N__8469),
            .in2(N__8439),
            .in3(N__8362),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13420),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI627QC51_6_LC_4_7_1.C_ON=1'b0;
    defparam beamY_RNI627QC51_6_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI627QC51_6_LC_4_7_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 beamY_RNI627QC51_6_LC_4_7_1 (
            .in0(N__10921),
            .in1(N__8509),
            .in2(N__9421),
            .in3(N__9637),
            .lcout(un4_row),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_4_8_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_4_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_4_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_4_8_0 (
            .in0(_gnd_net_),
            .in1(N__8983),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_4_8_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_4_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_4_8_1 (
            .in0(_gnd_net_),
            .in1(N__8520),
            .in2(N__8740),
            .in3(N__8281),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_4_8_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_4_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_4_8_2 (
            .in0(_gnd_net_),
            .in1(N__8770),
            .in2(N__8857),
            .in3(N__8266),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_4_8_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_4_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_4_8_3 (
            .in0(N__8244),
            .in1(N__8521),
            .in2(N__8827),
            .in3(N__8254),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_4_8_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_4_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_4_8_4 (
            .in0(_gnd_net_),
            .in1(N__8797),
            .in2(_gnd_net_),
            .in3(N__8251),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_4_9_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_4_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_4_9_0 (
            .in0(_gnd_net_),
            .in1(N__9846),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_4_9_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_4_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(N__8726),
            .in2(N__8530),
            .in3(N__8596),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(N__8593),
            .in2(N__8581),
            .in3(N__8566),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_4_9_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_4_9_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_4_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_4_9_3 (
            .in0(N__9950),
            .in1(N__8727),
            .in2(N__8563),
            .in3(N__8548),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_LUT4_0_LC_4_9_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_LUT4_0_LC_4_9_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_LUT4_0_LC_4_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_LUT4_0_LC_4_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8545),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_4_9_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_4_9_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_4_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9581),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_2_LC_4_9_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_2_LC_4_9_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_2_LC_4_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_2_LC_4_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8706),
            .lcout(un5_visiblex_i_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_4_9_7.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_4_9_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_4_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_4_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8766),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIOHGI2_LC_4_10_0.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIOHGI2_LC_4_10_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIOHGI2_LC_4_10_0.LUT_INIT=16'b0010001000000000;
    LogicCell40 un5_visiblex_cry_6_c_RNIOHGI2_LC_4_10_0 (
            .in0(N__8746),
            .in1(N__8728),
            .in2(_gnd_net_),
            .in3(N__9952),
            .lcout(),
            .ltout(un4_row_9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNI1GN17_LC_4_10_1.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNI1GN17_LC_4_10_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNI1GN17_LC_4_10_1.LUT_INIT=16'b0100000000000000;
    LogicCell40 un5_visiblex_cry_6_c_RNI1GN17_LC_4_10_1 (
            .in0(N__11374),
            .in1(N__10864),
            .in2(N__8512),
            .in3(N__10899),
            .lcout(un4_row_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_4_10_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_4_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_s_5_LC_4_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9657),
            .lcout(if_generate_plus_mult1_un54_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIK2PQ_LC_4_10_3.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIK2PQ_LC_4_10_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIK2PQ_LC_4_10_3.LUT_INIT=16'b0000000100001111;
    LogicCell40 un5_visiblex_cry_6_c_RNIK2PQ_LC_4_10_3 (
            .in0(N__8979),
            .in1(N__8905),
            .in2(N__11386),
            .in3(N__9136),
            .lcout(un4_row_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_4_10_6.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_4_10_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_4_10_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_1_LC_4_10_6 (
            .in0(N__8904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_LC_4_10_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_LC_4_10_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_c5_LC_4_10_7.LUT_INIT=16'b1001000111001000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_c5_LC_4_10_7 (
            .in0(N__8978),
            .in1(N__8903),
            .in2(N__8713),
            .in3(N__9135),
            .lcout(column_1_if_generate_plus_mult1_un47_sum_cZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_4_11_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_4_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_4_11_0 (
            .in0(_gnd_net_),
            .in1(N__8697),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_4_11_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_4_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_4_11_1 (
            .in0(_gnd_net_),
            .in1(N__9144),
            .in2(N__8920),
            .in3(N__8650),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_4_11_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_4_11_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_4_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_4_11_2 (
            .in0(_gnd_net_),
            .in1(N__9172),
            .in2(N__8647),
            .in3(N__8632),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_4_11_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_4_11_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_4_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_4_11_3 (
            .in0(N__9768),
            .in1(N__9145),
            .in2(N__8629),
            .in3(N__8614),
            .lcout(charx_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_4_11_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_4_11_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_4_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_4_11_4 (
            .in0(_gnd_net_),
            .in1(N__8611),
            .in2(_gnd_net_),
            .in3(N__8599),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1),
            .ltout(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_4_11_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_4_11_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_4_11_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_4_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8986),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_4_11_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_4_11_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_4_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_4_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8968),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_4_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9839),
            .lcout(un5_visiblex_i_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_4_12_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_4_12_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_4_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_4_12_0 (
            .in0(_gnd_net_),
            .in1(N__8902),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_4_12_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_4_12_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_4_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_4_12_1 (
            .in0(_gnd_net_),
            .in1(N__9024),
            .in2(N__9061),
            .in3(N__8845),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_4_12_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_4_12_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_4_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_4_12_2 (
            .in0(_gnd_net_),
            .in1(N__9039),
            .in2(N__8842),
            .in3(N__8815),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_4_12_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_4_12_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_4_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_4_12_3 (
            .in0(N__8765),
            .in1(N__9025),
            .in2(N__8812),
            .in3(N__8788),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_4_12_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_4_12_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_4_12_4.LUT_INIT=16'b0110011010011001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_4_12_4 (
            .in0(N__8785),
            .in1(N__9040),
            .in2(_gnd_net_),
            .in3(N__8773),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_4_12_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_4_12_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_4_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_4_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9168),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_4_12_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_4_12_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_4_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_4_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9132),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_4_13_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_4_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_4_13_0 (
            .in0(_gnd_net_),
            .in1(N__15600),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_4_13_1.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_4_13_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_4_13_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_4_13_1 (
            .in0(_gnd_net_),
            .in1(N__9052),
            .in2(_gnd_net_),
            .in3(N__9043),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_4_13_6.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_4_13_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_4_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_4_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9038),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_14_LC_5_3_0.C_ON=1'b0;
    defparam Pixel_RNO_14_LC_5_3_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_14_LC_5_3_0.LUT_INIT=16'b0000100000000010;
    LogicCell40 Pixel_RNO_14_LC_5_3_0 (
            .in0(N__13092),
            .in1(N__9887),
            .in2(N__13295),
            .in3(N__12913),
            .lcout(Pixel_RNOZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_15_LC_5_3_1.C_ON=1'b0;
    defparam Pixel_RNO_15_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_15_LC_5_3_1.LUT_INIT=16'b0001001000000000;
    LogicCell40 Pixel_RNO_15_LC_5_3_1 (
            .in0(N__12912),
            .in1(N__13283),
            .in2(N__9901),
            .in3(N__9510),
            .lcout(font_un126_pixel_5_a0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_19_LC_5_4_0.C_ON=1'b0;
    defparam Pixel_RNO_19_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_19_LC_5_4_0.LUT_INIT=16'b1111111111010000;
    LogicCell40 Pixel_RNO_19_LC_5_4_0 (
            .in0(N__9853),
            .in1(N__10132),
            .in2(N__13288),
            .in3(N__9504),
            .lcout(N_1740_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_54_LC_5_4_1.C_ON=1'b0;
    defparam Pixel_RNO_54_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_54_LC_5_4_1.LUT_INIT=16'b0001100001000010;
    LogicCell40 Pixel_RNO_54_LC_5_4_1 (
            .in0(N__11181),
            .in1(N__10125),
            .in2(N__12673),
            .in3(N__12917),
            .lcout(font_un28_pixel_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM1QKG9_0_3_LC_5_4_2.C_ON=1'b0;
    defparam beamY_RNIM1QKG9_0_3_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIM1QKG9_0_3_LC_5_4_2.LUT_INIT=16'b0100001000100100;
    LogicCell40 beamY_RNIM1QKG9_0_3_LC_5_4_2 (
            .in0(N__10124),
            .in1(N__12665),
            .in2(N__12932),
            .in3(N__11180),
            .lcout(font_un28_pixel_29),
            .ltout(font_un28_pixel_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDA2GGA3_0_LC_5_4_3.C_ON=1'b0;
    defparam beamY_RNIDA2GGA3_0_LC_5_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIDA2GGA3_0_LC_5_4_3.LUT_INIT=16'b0000100101101100;
    LogicCell40 beamY_RNIDA2GGA3_0_LC_5_4_3 (
            .in0(N__9503),
            .in1(N__13099),
            .in2(N__9340),
            .in3(N__13262),
            .lcout(beamY_RNIDA2GGA3Z0Z_0),
            .ltout(beamY_RNIDA2GGA3Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_11_LC_5_4_4.C_ON=1'b0;
    defparam Pixel_RNO_11_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_11_LC_5_4_4.LUT_INIT=16'b0000001010001010;
    LogicCell40 Pixel_RNO_11_LC_5_4_4 (
            .in0(N__9328),
            .in1(N__9318),
            .in2(N__9247),
            .in3(N__9379),
            .lcout(N_19_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_32_LC_5_4_5.C_ON=1'b0;
    defparam Pixel_RNO_32_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_32_LC_5_4_5.LUT_INIT=16'b0101010101100110;
    LogicCell40 Pixel_RNO_32_LC_5_4_5 (
            .in0(N__9238),
            .in1(N__13263),
            .in2(_gnd_net_),
            .in3(N__9232),
            .lcout(N_15_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_28_LC_5_4_6.C_ON=1'b0;
    defparam Pixel_RNO_28_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_28_LC_5_4_6.LUT_INIT=16'b1110101100010100;
    LogicCell40 Pixel_RNO_28_LC_5_4_6 (
            .in0(N__9192),
            .in1(N__12918),
            .in2(N__9902),
            .in3(N__9502),
            .lcout(),
            .ltout(Pixel_RNOZ0Z_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_9_LC_5_4_7.C_ON=1'b0;
    defparam Pixel_RNO_9_LC_5_4_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_9_LC_5_4_7.LUT_INIT=16'b1111101101000000;
    LogicCell40 Pixel_RNO_9_LC_5_4_7 (
            .in0(N__13276),
            .in1(N__13100),
            .in2(N__9211),
            .in3(N__9397),
            .lcout(Pixel_RNOZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_52_LC_5_5_0.C_ON=1'b0;
    defparam Pixel_RNO_52_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_52_LC_5_5_0.LUT_INIT=16'b0010100000010100;
    LogicCell40 Pixel_RNO_52_LC_5_5_0 (
            .in0(N__12644),
            .in1(N__9894),
            .in2(N__12933),
            .in3(N__10090),
            .lcout(g1_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM1QKG9_3_LC_5_5_1.C_ON=1'b0;
    defparam beamY_RNIM1QKG9_3_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIM1QKG9_3_LC_5_5_1.LUT_INIT=16'b0011110010011001;
    LogicCell40 beamY_RNIM1QKG9_3_LC_5_5_1 (
            .in0(N__10117),
            .in1(N__12643),
            .in2(N__11182),
            .in3(N__12921),
            .lcout(chary_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_50_LC_5_5_2.C_ON=1'b0;
    defparam Pixel_RNO_50_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_50_LC_5_5_2.LUT_INIT=16'b0110110000111001;
    LogicCell40 Pixel_RNO_50_LC_5_5_2 (
            .in0(N__12922),
            .in1(N__12648),
            .in2(N__10765),
            .in3(N__10119),
            .lcout(),
            .ltout(chary_1_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_27_LC_5_5_3.C_ON=1'b0;
    defparam Pixel_RNO_27_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_27_LC_5_5_3.LUT_INIT=16'b0000000001011101;
    LogicCell40 Pixel_RNO_27_LC_5_5_3 (
            .in0(N__11827),
            .in1(N__10081),
            .in2(N__9400),
            .in3(N__9491),
            .lcout(N_1737_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_70_LC_5_5_4.C_ON=1'b0;
    defparam Pixel_RNO_70_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_70_LC_5_5_4.LUT_INIT=16'b0111100000101101;
    LogicCell40 Pixel_RNO_70_LC_5_5_4 (
            .in0(N__12926),
            .in1(N__10663),
            .in2(N__12670),
            .in3(N__10118),
            .lcout(),
            .ltout(chary_1_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_53_LC_5_5_5.C_ON=1'b0;
    defparam Pixel_RNO_53_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_53_LC_5_5_5.LUT_INIT=16'b1001111110011001;
    LogicCell40 Pixel_RNO_53_LC_5_5_5 (
            .in0(N__13264),
            .in1(N__13056),
            .in2(N__9391),
            .in3(N__10080),
            .lcout(),
            .ltout(g2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_31_LC_5_5_6.C_ON=1'b0;
    defparam Pixel_RNO_31_LC_5_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_31_LC_5_5_6.LUT_INIT=16'b0101000101100010;
    LogicCell40 Pixel_RNO_31_LC_5_5_6 (
            .in0(N__9492),
            .in1(N__9373),
            .in2(N__9388),
            .in3(N__9385),
            .lcout(un116_pixel_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_51_LC_5_5_7.C_ON=1'b0;
    defparam Pixel_RNO_51_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_51_LC_5_5_7.LUT_INIT=16'b1111111100110011;
    LogicCell40 Pixel_RNO_51_LC_5_5_7 (
            .in0(_gnd_net_),
            .in1(N__13055),
            .in2(_gnd_net_),
            .in3(N__13258),
            .lcout(N_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_22_LC_5_6_1.C_ON=1'b0;
    defparam Pixel_RNO_22_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_22_LC_5_6_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 Pixel_RNO_22_LC_5_6_1 (
            .in0(N__13481),
            .in1(N__12105),
            .in2(N__12671),
            .in3(N__12172),
            .lcout(g0_0_a3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_4_LC_5_6_2.C_ON=1'b0;
    defparam beamY_RNI2KA6_4_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_4_LC_5_6_2.LUT_INIT=16'b0111000011110000;
    LogicCell40 beamY_RNI2KA6_4_LC_5_6_2 (
            .in0(N__12456),
            .in1(N__12656),
            .in2(N__10840),
            .in3(N__12920),
            .lcout(),
            .ltout(un8_beamylto9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_0_9_LC_5_6_3.C_ON=1'b0;
    defparam beamY_RNISI4A_0_9_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_0_9_LC_5_6_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNISI4A_0_9_LC_5_6_3 (
            .in0(N__13480),
            .in1(N__12104),
            .in2(N__9355),
            .in3(N__12171),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_43_LC_5_6_5.C_ON=1'b0;
    defparam Pixel_RNO_43_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_43_LC_5_6_5.LUT_INIT=16'b0001110111100010;
    LogicCell40 Pixel_RNO_43_LC_5_6_5 (
            .in0(N__10057),
            .in1(N__10174),
            .in2(N__10159),
            .in3(N__9458),
            .lcout(N_134_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_23_LC_5_6_6.C_ON=1'b0;
    defparam Pixel_RNO_23_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_23_LC_5_6_6.LUT_INIT=16'b0000000100000000;
    LogicCell40 Pixel_RNO_23_LC_5_6_6 (
            .in0(N__12457),
            .in1(N__12328),
            .in2(N__12253),
            .in3(N__9550),
            .lcout(g0_0_a3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_62_LC_5_7_0.C_ON=1'b0;
    defparam Pixel_RNO_62_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_62_LC_5_7_0.LUT_INIT=16'b0000110001000100;
    LogicCell40 Pixel_RNO_62_LC_5_7_0 (
            .in0(N__10420),
            .in1(N__13226),
            .in2(N__11692),
            .in3(N__10267),
            .lcout(),
            .ltout(m4_rn_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_40_LC_5_7_1.C_ON=1'b0;
    defparam Pixel_RNO_40_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_40_LC_5_7_1.LUT_INIT=16'b0101010100001111;
    LogicCell40 Pixel_RNO_40_LC_5_7_1 (
            .in0(N__10540),
            .in1(_gnd_net_),
            .in2(N__9532),
            .in3(N__9406),
            .lcout(Pixel_RNOZ0Z_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram0__RNIR1C2R81_0_LC_5_7_2.C_ON=1'b0;
    defparam content_content_ram0__RNIR1C2R81_0_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam content_content_ram0__RNIR1C2R81_0_LC_5_7_2.LUT_INIT=16'b0111001111111011;
    LogicCell40 content_content_ram0__RNIR1C2R81_0_LC_5_7_2 (
            .in0(N__10461),
            .in1(N__10265),
            .in2(N__11691),
            .in3(N__10539),
            .lcout(),
            .ltout(content_content_ram0__RNIR1C2R81Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram0__RNIAENOV03_0_LC_5_7_3.C_ON=1'b0;
    defparam content_content_ram0__RNIAENOV03_0_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam content_content_ram0__RNIAENOV03_0_LC_5_7_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 content_content_ram0__RNIAENOV03_0_LC_5_7_3 (
            .in0(_gnd_net_),
            .in1(N__9643),
            .in2(N__9517),
            .in3(N__10419),
            .lcout(N_331_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0H2_0_4_LC_5_7_4.C_ON=1'b0;
    defparam beamY_RNIJ0H2_0_4_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0H2_0_4_LC_5_7_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIJ0H2_0_4_LC_5_7_4 (
            .in0(N__12642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12455),
            .lcout(),
            .ltout(un4_row_m7_ns_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPAQ91_6_LC_5_7_5.C_ON=1'b0;
    defparam beamY_RNIPAQ91_6_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIPAQ91_6_LC_5_7_5.LUT_INIT=16'b0100000110000010;
    LogicCell40 beamY_RNIPAQ91_6_LC_5_7_5 (
            .in0(N__10900),
            .in1(N__12324),
            .in2(N__9424),
            .in3(N__12243),
            .lcout(beamY_RNIPAQ91Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_9_LC_5_7_6.C_ON=1'b0;
    defparam beamY_RNISI4A_9_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_9_LC_5_7_6.LUT_INIT=16'b1100110011001000;
    LogicCell40 beamY_RNISI4A_9_LC_5_7_6 (
            .in0(N__12102),
            .in1(N__13486),
            .in2(N__10144),
            .in3(N__12164),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_63_LC_5_7_7.C_ON=1'b0;
    defparam Pixel_RNO_63_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_63_LC_5_7_7.LUT_INIT=16'b1010000000000000;
    LogicCell40 Pixel_RNO_63_LC_5_7_7 (
            .in0(N__10266),
            .in1(_gnd_net_),
            .in2(N__13265),
            .in3(N__10462),
            .lcout(m4_sn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram0__RNIR1C2R81_0_0_LC_5_8_1.C_ON=1'b0;
    defparam content_content_ram0__RNIR1C2R81_0_0_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam content_content_ram0__RNIR1C2R81_0_0_LC_5_8_1.LUT_INIT=16'b0100000011001000;
    LogicCell40 content_content_ram0__RNIR1C2R81_0_0_LC_5_8_1 (
            .in0(N__10459),
            .in1(N__10253),
            .in2(N__11684),
            .in3(N__10538),
            .lcout(content_content_ram0__RNIR1C2R81_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un6_rowlto3_LC_5_8_2.C_ON=1'b0;
    defparam un6_rowlto3_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam un6_rowlto3_LC_5_8_2.LUT_INIT=16'b0000000000010101;
    LogicCell40 un6_rowlto3_LC_5_8_2 (
            .in0(N__11659),
            .in1(N__10460),
            .in2(N__10264),
            .in3(N__11597),
            .lcout(un6_rowlt7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_5_9_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_5_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(N__10003),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_5_9_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_5_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(N__9676),
            .in2(N__9565),
            .in3(N__9619),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_5_9_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_5_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(N__9778),
            .in2(N__9697),
            .in3(N__9604),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_5_9_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_5_9_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_5_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_5_9_3 (
            .in0(N__9582),
            .in1(N__9556),
            .in2(N__9748),
            .in3(N__9592),
            .lcout(charx_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_5_9_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_5_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_5_9_4 (
            .in0(_gnd_net_),
            .in1(N__9715),
            .in2(_gnd_net_),
            .in3(N__9589),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_9_6.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9847),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_5_9_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_5_9_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_5_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_5_9_7 (
            .in0(N__9747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9692),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_5_10_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_5_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__9842),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_5_10_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_5_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(N__9732),
            .in2(N__9790),
            .in3(N__9772),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_5_10_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_5_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_5_10_2 (
            .in0(_gnd_net_),
            .in1(N__9769),
            .in2(N__9757),
            .in3(N__9736),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_5_10_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_5_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_5_10_3 (
            .in0(N__9696),
            .in1(N__9733),
            .in2(N__9724),
            .in3(N__9709),
            .lcout(charx_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_5_10_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_5_10_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_5_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(N__9706),
            .in2(_gnd_net_),
            .in3(N__9700),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3),
            .ltout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_5_10_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_5_10_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_5_10_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_5_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9679),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_5_11_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_5_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(N__9995),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_11_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(N__9670),
            .in2(N__9664),
            .in3(N__9646),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(N__9951),
            .in2(N__10051),
            .in3(N__10039),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_5_11_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_5_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_5_11_3 (
            .in0(N__11570),
            .in1(N__9928),
            .in2(N__10036),
            .in3(N__10024),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_5_11_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_5_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_s_5_LC_5_11_4 (
            .in0(_gnd_net_),
            .in1(N__10021),
            .in2(_gnd_net_),
            .in3(N__10012),
            .lcout(if_generate_plus_mult1_un61_sum_s_5),
            .ltout(if_generate_plus_mult1_un61_sum_s_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_5_11_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_5_11_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_5_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10009),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_5_11_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_5_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_i_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9996),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_11_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9949),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_59_LC_6_4_0.C_ON=1'b0;
    defparam Pixel_RNO_59_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_59_LC_6_4_0.LUT_INIT=16'b0110010110101001;
    LogicCell40 Pixel_RNO_59_LC_6_4_0 (
            .in0(N__12664),
            .in1(N__12930),
            .in2(N__10126),
            .in3(N__10690),
            .lcout(chary_2_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI539IG9_3_LC_6_4_2.C_ON=1'b0;
    defparam beamY_RNI539IG9_3_LC_6_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI539IG9_3_LC_6_4_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNI539IG9_3_LC_6_4_2 (
            .in0(N__12018),
            .in1(N__11862),
            .in2(N__11128),
            .in3(N__11179),
            .lcout(beamY_RNI539IG9Z0Z_3),
            .ltout(beamY_RNI539IG9Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_42_LC_6_4_3.C_ON=1'b0;
    defparam Pixel_RNO_42_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_42_LC_6_4_3.LUT_INIT=16'b0000111111110000;
    LogicCell40 Pixel_RNO_42_LC_6_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9856),
            .in3(N__12886),
            .lcout(g4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_41_LC_6_4_7.C_ON=1'b0;
    defparam Pixel_RNO_41_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_41_LC_6_4_7.LUT_INIT=16'b0111100001001011;
    LogicCell40 Pixel_RNO_41_LC_6_4_7 (
            .in0(N__10063),
            .in1(N__12887),
            .in2(N__12672),
            .in3(N__10120),
            .lcout(chary_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6CM834_3_LC_6_5_1.C_ON=1'b0;
    defparam beamY_RNI6CM834_3_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI6CM834_3_LC_6_5_1.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI6CM834_3_LC_6_5_1 (
            .in0(N__11109),
            .in1(N__12003),
            .in2(_gnd_net_),
            .in3(N__11863),
            .lcout(chary_if_generate_plus_mult1_un75_sum_axbxc5_1),
            .ltout(chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_69_LC_6_5_2.C_ON=1'b0;
    defparam Pixel_RNO_69_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_69_LC_6_5_2.LUT_INIT=16'b0110011000001111;
    LogicCell40 Pixel_RNO_69_LC_6_5_2 (
            .in0(N__15059),
            .in1(N__11938),
            .in2(N__10093),
            .in3(N__12888),
            .lcout(g1_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_78_LC_6_5_3.C_ON=1'b0;
    defparam Pixel_RNO_78_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_78_LC_6_5_3.LUT_INIT=16'b1000101000101010;
    LogicCell40 Pixel_RNO_78_LC_6_5_3 (
            .in0(N__14718),
            .in1(N__14974),
            .in2(N__10186),
            .in3(N__14278),
            .lcout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMSO1N7_0_2_LC_6_5_4.C_ON=1'b0;
    defparam beamY_RNIMSO1N7_0_2_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIMSO1N7_0_2_LC_6_5_4.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIMSO1N7_0_2_LC_6_5_4 (
            .in0(N__12004),
            .in1(N__11167),
            .in2(N__12934),
            .in3(N__11110),
            .lcout(),
            .ltout(beamY_RNIMSO1N7_0Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJEAL7H_2_LC_6_5_5.C_ON=1'b0;
    defparam beamY_RNIJEAL7H_2_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIJEAL7H_2_LC_6_5_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 beamY_RNIJEAL7H_2_LC_6_5_5 (
            .in0(_gnd_net_),
            .in1(N__10672),
            .in2(N__10084),
            .in3(N__11864),
            .lcout(g4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_79_LC_6_5_6.C_ON=1'b0;
    defparam Pixel_RNO_79_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_79_LC_6_5_6.LUT_INIT=16'b0110100100000000;
    LogicCell40 Pixel_RNO_79_LC_6_5_6 (
            .in0(N__14279),
            .in1(N__10185),
            .in2(N__14985),
            .in3(N__10168),
            .lcout(),
            .ltout(g2_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_64_LC_6_5_7.C_ON=1'b0;
    defparam Pixel_RNO_64_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_64_LC_6_5_7.LUT_INIT=16'b0110011000110110;
    LogicCell40 Pixel_RNO_64_LC_6_5_7 (
            .in0(N__10072),
            .in1(N__15058),
            .in2(N__10066),
            .in3(N__12005),
            .lcout(chary_if_generate_plus_mult1_un68_sum_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_66_LC_6_6_0.C_ON=1'b0;
    defparam Pixel_RNO_66_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_66_LC_6_6_0.LUT_INIT=16'b0001010001000001;
    LogicCell40 Pixel_RNO_66_LC_6_6_0 (
            .in0(N__12654),
            .in1(N__12014),
            .in2(N__11127),
            .in3(N__11865),
            .lcout(Pixel_RNOZ0Z_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_2_4_LC_6_6_1.C_ON=1'b0;
    defparam beamY_RNIBFP3_2_4_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_2_4_LC_6_6_1.LUT_INIT=16'b0110011010101010;
    LogicCell40 beamY_RNIBFP3_2_4_LC_6_6_1 (
            .in0(N__12460),
            .in1(N__12652),
            .in2(_gnd_net_),
            .in3(N__12878),
            .lcout(un5_visibley_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_65_LC_6_6_2.C_ON=1'b0;
    defparam Pixel_RNO_65_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_65_LC_6_6_2.LUT_INIT=16'b0101011010101001;
    LogicCell40 Pixel_RNO_65_LC_6_6_2 (
            .in0(N__12880),
            .in1(N__10717),
            .in2(N__10741),
            .in3(N__15067),
            .lcout(g2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_87_LC_6_6_3.C_ON=1'b0;
    defparam Pixel_RNO_87_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_87_LC_6_6_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 Pixel_RNO_87_LC_6_6_3 (
            .in0(_gnd_net_),
            .in1(N__12653),
            .in2(_gnd_net_),
            .in3(N__12879),
            .lcout(un5_visibley_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_67_LC_6_6_5.C_ON=1'b0;
    defparam Pixel_RNO_67_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_67_LC_6_6_5.LUT_INIT=16'b1001011000000000;
    LogicCell40 Pixel_RNO_67_LC_6_6_5 (
            .in0(N__11866),
            .in1(N__11123),
            .in2(N__12019),
            .in3(N__12655),
            .lcout(Pixel_RNOZ0Z_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4H2_6_LC_6_7_1.C_ON=1'b0;
    defparam beamY_RNIN4H2_6_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4H2_6_LC_6_7_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIN4H2_6_LC_6_7_1 (
            .in0(N__12322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12241),
            .lcout(un8_beamy_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_1_3_LC_6_7_3.C_ON=1'b0;
    defparam beamY_RNIHUG2_1_3_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_1_3_LC_6_7_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIHUG2_1_3_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(N__12588),
            .in2(_gnd_net_),
            .in3(N__12838),
            .lcout(),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_6_LC_6_7_4.C_ON=1'b0;
    defparam beamY_RNI2KA6_6_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_6_LC_6_7_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI2KA6_6_LC_6_7_4 (
            .in0(N__12242),
            .in1(N__12441),
            .in2(N__10147),
            .in3(N__12323),
            .lcout(un4_beamylt8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_8_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_8_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_6_8_5.C_ON=1'b0;
    defparam beamY_0_LC_6_8_5.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_6_8_5.LUT_INIT=16'b0101010100100010;
    LogicCell40 beamY_0_LC_6_8_5 (
            .in0(N__13391),
            .in1(N__13531),
            .in2(_gnd_net_),
            .in3(N__13026),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13421),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_6_8_6.C_ON=1'b0;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_6_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_6_8_6 (
            .in0(N__14358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_Clock12MHz_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_6_9_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_6_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__10344),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_6_9_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_6_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_6_9_1 (
            .in0(_gnd_net_),
            .in1(N__10278),
            .in2(N__10240),
            .in3(N__10445),
            .lcout(G_383),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_6_9_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_6_9_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__10448),
            .in2(N__10198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_LC_6_9_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_LC_6_9_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_4_c_LC_6_9_3 (
            .in0(_gnd_net_),
            .in1(N__10279),
            .in2(N__10495),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_6_9_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_6_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_s_5_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__10483),
            .in2(_gnd_net_),
            .in3(N__10270),
            .lcout(un6_rowlto0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_9_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_i_LC_6_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10231),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_10_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(N__10230),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_6_10_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_6_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(N__10549),
            .in2(N__10471),
            .in3(N__10189),
            .lcout(if_generate_plus_mult1_un75_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(N__11643),
            .in2(N__10396),
            .in3(N__10486),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_6_10_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_6_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_6_10_3 (
            .in0(N__10446),
            .in1(N__10614),
            .in2(N__10603),
            .in3(N__10477),
            .lcout(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_6_10_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_6_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_s_5_LC_6_10_4 (
            .in0(_gnd_net_),
            .in1(N__10636),
            .in2(_gnd_net_),
            .in3(N__10474),
            .lcout(un6_rowlto1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_column_1_i_2_sbtinv_2_LC_6_10_5.C_ON=1'b0;
    defparam content_column_1_i_2_sbtinv_2_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam content_column_1_i_2_sbtinv_2_LC_6_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 content_column_1_i_2_sbtinv_2_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11641),
            .lcout(content_column_1_i_2_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram5__RNIKAVJ9F_0_LC_6_10_7.C_ON=1'b0;
    defparam content_content_ram5__RNIKAVJ9F_0_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam content_content_ram5__RNIKAVJ9F_0_LC_6_10_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 content_content_ram5__RNIKAVJ9F_0_LC_6_10_7 (
            .in0(N__10447),
            .in1(_gnd_net_),
            .in2(N__11056),
            .in3(N__10510),
            .lcout(content_N_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(N__10593),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__10371),
            .in2(N__10405),
            .in3(N__10387),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(N__11571),
            .in2(N__10384),
            .in3(N__10375),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3 (
            .in0(N__11642),
            .in1(N__10372),
            .in2(N__10645),
            .in3(N__10630),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(N__10627),
            .in2(_gnd_net_),
            .in3(N__10621),
            .lcout(content_column_1_i_2_2),
            .ltout(content_column_1_i_2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_6_11_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_6_11_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10618),
            .in3(N__10615),
            .lcout(if_generate_plus_mult1_un75_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_i_LC_6_11_7 (
            .in0(N__10594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram8__e_0_RNI0I9HN1_0_LC_6_12_1.C_ON=1'b0;
    defparam content_content_ram8__e_0_RNI0I9HN1_0_LC_6_12_1.SEQ_MODE=4'b0000;
    defparam content_content_ram8__e_0_RNI0I9HN1_0_LC_6_12_1.LUT_INIT=16'b0100010101100111;
    LogicCell40 content_content_ram8__e_0_RNI0I9HN1_0_LC_6_12_1 (
            .in0(N__11646),
            .in1(N__11574),
            .in2(N__11812),
            .in3(N__11365),
            .lcout(),
            .ltout(content_m7_ns_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram0__RNIEAKG02_0_LC_6_12_2.C_ON=1'b0;
    defparam content_content_ram0__RNIEAKG02_0_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam content_content_ram0__RNIEAKG02_0_LC_6_12_2.LUT_INIT=16'b0111000001111010;
    LogicCell40 content_content_ram0__RNIEAKG02_0_LC_6_12_2 (
            .in0(N__11575),
            .in1(N__11779),
            .in2(N__10543),
            .in3(N__11499),
            .lcout(content_N_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_LC_6_12_4.C_ON=1'b0;
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_LC_6_12_4.LUT_INIT=16'b1101100010101010;
    LogicCell40 content_content_ram11__e_0_RNIQ1Q3O1_0_LC_6_12_4 (
            .in0(N__11573),
            .in1(N__11526),
            .in2(N__11035),
            .in3(N__11645),
            .lcout(),
            .ltout(content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram7__RNI6B0NG3_0_LC_6_12_5.C_ON=1'b0;
    defparam content_content_ram7__RNI6B0NG3_0_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam content_content_ram7__RNI6B0NG3_0_LC_6_12_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 content_content_ram7__RNI6B0NG3_0_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(N__11721),
            .in2(N__10513),
            .in3(N__10501),
            .lcout(content_content_ram7__RNI6B0NG3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_0_LC_6_12_6.C_ON=1'b0;
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_0_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam content_content_ram11__e_0_RNIQ1Q3O1_0_0_LC_6_12_6.LUT_INIT=16'b1100100001000000;
    LogicCell40 content_content_ram11__e_0_RNIQ1Q3O1_0_0_LC_6_12_6 (
            .in0(N__11572),
            .in1(N__11644),
            .in2(N__11034),
            .in3(N__11525),
            .lcout(content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_92_LC_7_4_0.C_ON=1'b0;
    defparam Pixel_RNO_92_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_92_LC_7_4_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 Pixel_RNO_92_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__12660),
            .in2(_gnd_net_),
            .in3(N__12881),
            .lcout(un5_visibley_2_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_85_LC_7_4_1.C_ON=1'b0;
    defparam Pixel_RNO_85_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_85_LC_7_4_1.LUT_INIT=16'b1010001000101010;
    LogicCell40 Pixel_RNO_85_LC_7_4_1 (
            .in0(N__14719),
            .in1(N__10992),
            .in2(N__14984),
            .in3(N__14281),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_75_LC_7_4_2.C_ON=1'b0;
    defparam Pixel_RNO_75_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_75_LC_7_4_2.LUT_INIT=16'b0011110000110110;
    LogicCell40 Pixel_RNO_75_LC_7_4_2 (
            .in0(N__10678),
            .in1(N__15063),
            .in2(N__10693),
            .in3(N__12002),
            .lcout(chary_if_generate_plus_mult1_un68_sum_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_86_LC_7_4_3.C_ON=1'b0;
    defparam Pixel_RNO_86_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_86_LC_7_4_3.LUT_INIT=16'b0010100010000010;
    LogicCell40 Pixel_RNO_86_LC_7_4_3 (
            .in0(N__10684),
            .in1(N__10993),
            .in2(N__14983),
            .in3(N__14282),
            .lcout(g2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMSO1N7_2_LC_7_5_0.C_ON=1'b0;
    defparam beamY_RNIMSO1N7_2_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIMSO1N7_2_LC_7_5_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIMSO1N7_2_LC_7_5_0 (
            .in0(N__11994),
            .in1(N__11155),
            .in2(N__11119),
            .in3(N__12882),
            .lcout(beamY_RNIMSO1N7Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_82_LC_7_5_2.C_ON=1'b0;
    defparam Pixel_RNO_82_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_82_LC_7_5_2.LUT_INIT=16'b1000010011001100;
    LogicCell40 Pixel_RNO_82_LC_7_5_2 (
            .in0(N__14277),
            .in1(N__14703),
            .in2(N__14986),
            .in3(N__10702),
            .lcout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_91_LC_7_5_3.C_ON=1'b0;
    defparam Pixel_RNO_91_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_91_LC_7_5_3.LUT_INIT=16'b1000101000101010;
    LogicCell40 Pixel_RNO_91_LC_7_5_3 (
            .in0(N__14702),
            .in1(N__14982),
            .in2(N__11929),
            .in3(N__14275),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_84_LC_7_5_4.C_ON=1'b0;
    defparam Pixel_RNO_84_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_84_LC_7_5_4.LUT_INIT=16'b0000101111110100;
    LogicCell40 Pixel_RNO_84_LC_7_5_4 (
            .in0(N__11993),
            .in1(N__10654),
            .in2(N__10666),
            .in3(N__15056),
            .lcout(chary_if_generate_plus_mult1_un68_sum_1_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6C1MV_3_LC_7_5_5.C_ON=1'b0;
    defparam beamY_RNI6C1MV_3_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI6C1MV_3_LC_7_5_5.LUT_INIT=16'b0110000010010000;
    LogicCell40 beamY_RNI6C1MV_3_LC_7_5_5 (
            .in0(N__10701),
            .in1(N__14981),
            .in2(N__11137),
            .in3(N__14276),
            .lcout(g2_0),
            .ltout(g2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_68_LC_7_5_6.C_ON=1'b0;
    defparam Pixel_RNO_68_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_68_LC_7_5_6.LUT_INIT=16'b0010001111011100;
    LogicCell40 Pixel_RNO_68_LC_7_5_6 (
            .in0(N__11995),
            .in1(N__10774),
            .in2(N__10768),
            .in3(N__15057),
            .lcout(chary_if_generate_plus_mult1_un68_sum_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSyncZ0_LC_7_5_7.C_ON=1'b0;
    defparam VSyncZ0_LC_7_5_7.SEQ_MODE=4'b1000;
    defparam VSyncZ0_LC_7_5_7.LUT_INIT=16'b1111011101110111;
    LogicCell40 VSyncZ0_LC_7_5_7 (
            .in0(N__11074),
            .in1(N__10711),
            .in2(N__12919),
            .in3(N__13251),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13425),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_80_LC_7_6_0.C_ON=1'b0;
    defparam Pixel_RNO_80_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_80_LC_7_6_0.LUT_INIT=16'b1000101000101010;
    LogicCell40 Pixel_RNO_80_LC_7_6_0 (
            .in0(N__14717),
            .in1(N__14949),
            .in2(N__10732),
            .in3(N__14284),
            .lcout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_4_4_LC_7_6_1.C_ON=1'b0;
    defparam beamY_RNIBFP3_4_4_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_4_4_LC_7_6_1.LUT_INIT=16'b0110011010101010;
    LogicCell40 beamY_RNIBFP3_4_4_LC_7_6_1 (
            .in0(N__12458),
            .in1(N__12649),
            .in2(_gnd_net_),
            .in3(N__12875),
            .lcout(un5_visibley_3_28),
            .ltout(un5_visibley_3_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_88_LC_7_6_2.C_ON=1'b0;
    defparam Pixel_RNO_88_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_88_LC_7_6_2.LUT_INIT=16'b0011110011000011;
    LogicCell40 Pixel_RNO_88_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(N__14948),
            .in2(N__10723),
            .in3(N__14283),
            .lcout(),
            .ltout(g1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_81_LC_7_6_3.C_ON=1'b0;
    defparam Pixel_RNO_81_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_81_LC_7_6_3.LUT_INIT=16'b0001000001000000;
    LogicCell40 Pixel_RNO_81_LC_7_6_3 (
            .in0(N__11984),
            .in1(N__12651),
            .in2(N__10720),
            .in3(N__12877),
            .lcout(g2_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_RNO_1_LC_7_6_5.C_ON=1'b0;
    defparam VSync_RNO_1_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam VSync_RNO_1_LC_7_6_5.LUT_INIT=16'b0000000000100010;
    LogicCell40 VSync_RNO_1_LC_7_6_5 (
            .in0(N__10839),
            .in1(N__13485),
            .in2(_gnd_net_),
            .in3(N__12106),
            .lcout(un1_beamylto9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_1_4_LC_7_6_7.C_ON=1'b0;
    defparam beamY_RNIBFP3_1_4_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_1_4_LC_7_6_7.LUT_INIT=16'b0110011010101010;
    LogicCell40 beamY_RNIBFP3_1_4_LC_7_6_7 (
            .in0(N__12459),
            .in1(N__12650),
            .in2(_gnd_net_),
            .in3(N__12876),
            .lcout(un5_visibley_1_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_7_7_0.C_ON=1'b0;
    defparam beamY_1_LC_7_7_0.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_7_7_0.LUT_INIT=16'b0001001010101010;
    LogicCell40 beamY_1_LC_7_7_0 (
            .in0(N__13156),
            .in1(N__13520),
            .in2(N__13074),
            .in3(N__13384),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI70BUG1_LC_7_7_2.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI70BUG1_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI70BUG1_LC_7_7_2.LUT_INIT=16'b0001100010001000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI70BUG1_LC_7_7_2 (
            .in0(N__10792),
            .in1(N__10950),
            .in2(N__10816),
            .in3(N__10974),
            .lcout(),
            .ltout(chessboardpixel_un200_pixellto4_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQF0E52_1_LC_7_7_3.C_ON=1'b0;
    defparam beamY_RNIQF0E52_1_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIQF0E52_1_LC_7_7_3.LUT_INIT=16'b1000000001000000;
    LogicCell40 beamY_RNIQF0E52_1_LC_7_7_3 (
            .in0(N__10975),
            .in1(N__13155),
            .in2(N__10855),
            .in3(N__10814),
            .lcout(chessboardpixel_un200_pixellt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIID25_0_7_LC_7_7_4.C_ON=1'b0;
    defparam beamY_RNIID25_0_7_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIID25_0_7_LC_7_7_4.LUT_INIT=16'b0100010000000000;
    LogicCell40 beamY_RNIID25_0_7_LC_7_7_4 (
            .in0(N__12103),
            .in1(N__10838),
            .in2(_gnd_net_),
            .in3(N__12165),
            .lcout(un5_beamx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_7_7_5.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_7_7_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_3_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(N__12587),
            .in2(_gnd_net_),
            .in3(N__12806),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_7_7_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_7_7_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_7_7_6 (
            .in0(N__12807),
            .in1(N__15483),
            .in2(_gnd_net_),
            .in3(N__10815),
            .lcout(beamY_i_2),
            .ltout(beamY_i_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_0_LC_7_7_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_0_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_0_LC_7_7_7.LUT_INIT=16'b1111111100001111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_0_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10819),
            .in3(N__10791),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_8_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__10810),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_LC_7_8_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_LC_7_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__10927),
            .in2(N__11328),
            .in3(N__10783),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLG_LC_7_8_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLG_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLG_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLG_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__11323),
            .in2(N__11212),
            .in3(N__10780),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777J_LC_7_8_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777J_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777J_LC_7_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777J_LC_7_8_3 (
            .in0(_gnd_net_),
            .in1(N__11200),
            .in2(N__11329),
            .in3(N__10777),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_8_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__10984),
            .in2(N__11353),
            .in3(N__11319),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEK_LC_7_8_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEK_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEK_LC_7_8_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEK_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(N__11341),
            .in2(_gnd_net_),
            .in3(N__10978),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIN7I542_LC_7_8_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIN7I542_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIN7I542_LC_7_8_6.LUT_INIT=16'b1010101010011010;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIN7I542_LC_7_8_6 (
            .in0(N__10966),
            .in1(N__10960),
            .in2(N__10954),
            .in3(N__10951),
            .lcout(chessboardpixel_un178_pixel_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_7_8_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_7_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11229),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_7_9_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_7_9_1.LUT_INIT=16'b0110111000010111;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_7_9_1 (
            .in0(N__15190),
            .in1(N__15709),
            .in2(N__15295),
            .in3(N__15121),
            .lcout(if_generate_plus_mult1_un54_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_c5_LC_7_10_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_c5_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_c5_LC_7_10_0.LUT_INIT=16'b0000110111110100;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_c5_LC_7_10_0 (
            .in0(N__10886),
            .in1(N__14791),
            .in2(N__10909),
            .in3(N__15290),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_cZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_axb3_LC_7_10_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_axb3_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_axb3_LC_7_10_1.LUT_INIT=16'b1000100001100110;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_axb3_LC_7_10_1 (
            .in0(N__15191),
            .in1(N__15717),
            .in2(_gnd_net_),
            .in3(N__15122),
            .lcout(row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3),
            .ltout(row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_7_10_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_7_10_2.LUT_INIT=16'b1101001001001011;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_7_10_2 (
            .in0(N__10885),
            .in1(N__14790),
            .in2(N__10867),
            .in3(N__15289),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram9__e_0_RNIFBHPN1_0_LC_7_11_1.C_ON=1'b0;
    defparam content_content_ram9__e_0_RNIFBHPN1_0_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam content_content_ram9__e_0_RNIFBHPN1_0_LC_7_11_1.LUT_INIT=16'b1110011011000100;
    LogicCell40 content_content_ram9__e_0_RNIFBHPN1_0_LC_7_11_1 (
            .in0(N__11652),
            .in1(N__11589),
            .in2(N__13726),
            .in3(N__11043),
            .lcout(content_content_ram9__e_0_RNIFBHPN1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram9__e_0_RNIFBHPN1_0_0_LC_7_11_2.C_ON=1'b0;
    defparam content_content_ram9__e_0_RNIFBHPN1_0_0_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam content_content_ram9__e_0_RNIFBHPN1_0_0_LC_7_11_2.LUT_INIT=16'b1101100000000000;
    LogicCell40 content_content_ram9__e_0_RNIFBHPN1_0_0_LC_7_11_2 (
            .in0(N__11590),
            .in1(N__13725),
            .in2(N__11047),
            .in3(N__11653),
            .lcout(),
            .ltout(content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram5__RNIEM2QF3_0_LC_7_11_3.C_ON=1'b0;
    defparam content_content_ram5__RNIEM2QF3_0_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam content_content_ram5__RNIEM2QF3_0_LC_7_11_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 content_content_ram5__RNIEM2QF3_0_LC_7_11_3 (
            .in0(_gnd_net_),
            .in1(N__11460),
            .in2(N__11065),
            .in3(N__11062),
            .lcout(content_content_ram5__RNIEM2QF3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram9__e_0_0_LC_7_11_5.C_ON=1'b0;
    defparam content_content_ram9__e_0_0_LC_7_11_5.SEQ_MODE=4'b1000;
    defparam content_content_ram9__e_0_0_LC_7_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 content_content_ram9__e_0_0_LC_7_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14539),
            .lcout(content_ram9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14339),
            .ce(N__11506),
            .sr(_gnd_net_));
    defparam content_content_ram11__e_0_0_LC_7_12_0.C_ON=1'b0;
    defparam content_content_ram11__e_0_0_LC_7_12_0.SEQ_MODE=4'b1000;
    defparam content_content_ram11__e_0_0_LC_7_12_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 content_content_ram11__e_0_0_LC_7_12_0 (
            .in0(N__14542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(content_ram11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14340),
            .ce(N__11470),
            .sr(_gnd_net_));
    defparam nCS1_1_LC_7_14_0.C_ON=1'b0;
    defparam nCS1_1_LC_7_14_0.SEQ_MODE=4'b1001;
    defparam nCS1_1_LC_7_14_0.LUT_INIT=16'b1011111100010101;
    LogicCell40 nCS1_1_LC_7_14_0 (
            .in0(N__14436),
            .in1(N__14191),
            .in2(N__14581),
            .in3(N__11004),
            .lcout(nCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14344),
            .ce(),
            .sr(N__11701));
    defparam beamY_RNIBFP3_3_4_LC_8_4_3.C_ON=1'b0;
    defparam beamY_RNIBFP3_3_4_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_3_4_LC_8_4_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 beamY_RNIBFP3_3_4_LC_8_4_3 (
            .in0(N__12858),
            .in1(N__12438),
            .in2(_gnd_net_),
            .in3(N__12600),
            .lcout(un5_visibley_2_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4QL4A1_4_LC_8_5_1.C_ON=1'b0;
    defparam beamY_RNI4QL4A1_4_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI4QL4A1_4_LC_8_5_1.LUT_INIT=16'b1001000011110000;
    LogicCell40 beamY_RNI4QL4A1_4_LC_8_5_1 (
            .in0(N__14266),
            .in1(N__14951),
            .in2(N__14715),
            .in3(N__14827),
            .lcout(chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPAS0A1_4_LC_8_5_3.C_ON=1'b0;
    defparam beamY_RNIPAS0A1_4_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIPAS0A1_4_LC_8_5_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 beamY_RNIPAS0A1_4_LC_8_5_3 (
            .in0(N__14267),
            .in1(_gnd_net_),
            .in2(N__14716),
            .in3(N__14950),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6C1MV_1_3_LC_8_5_4.C_ON=1'b0;
    defparam beamY_RNI6C1MV_1_3_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI6C1MV_1_3_LC_8_5_4.LUT_INIT=16'b0110000010010000;
    LogicCell40 beamY_RNI6C1MV_1_3_LC_8_5_4 (
            .in0(N__14952),
            .in1(N__14828),
            .in2(N__11239),
            .in3(N__14265),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVMI9D5_3_LC_8_5_5.C_ON=1'b0;
    defparam beamY_RNIVMI9D5_3_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIVMI9D5_3_LC_8_5_5.LUT_INIT=16'b0101010110011010;
    LogicCell40 beamY_RNIVMI9D5_3_LC_8_5_5 (
            .in0(N__15052),
            .in1(N__11983),
            .in2(N__11191),
            .in3(N__11188),
            .lcout(beamY_RNIVMI9D5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_8_5_6.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_8_5_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_0_3_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(N__12636),
            .in2(_gnd_net_),
            .in3(N__12857),
            .lcout(un5_visibley_1_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6C1MV_0_3_LC_8_5_7.C_ON=1'b0;
    defparam beamY_RNI6C1MV_0_3_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI6C1MV_0_3_LC_8_5_7.LUT_INIT=16'b0110111100000110;
    LogicCell40 beamY_RNI6C1MV_0_3_LC_8_5_7 (
            .in0(N__14268),
            .in1(N__14953),
            .in2(N__14846),
            .in3(N__11238),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8325_6_LC_8_6_1.C_ON=1'b0;
    defparam beamY_RNI8325_6_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI8325_6_LC_8_6_1.LUT_INIT=16'b1111111011101110;
    LogicCell40 beamY_RNI8325_6_LC_8_6_1 (
            .in0(N__12227),
            .in1(N__12308),
            .in2(N__12586),
            .in3(N__12750),
            .lcout(),
            .ltout(beamY_RNI8325Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPOR8_6_LC_8_6_2.C_ON=1'b0;
    defparam beamY_RNIPOR8_6_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIPOR8_6_LC_8_6_2.LUT_INIT=16'b1111001111100010;
    LogicCell40 beamY_RNIPOR8_6_LC_8_6_2 (
            .in0(N__12309),
            .in1(N__12406),
            .in2(N__11080),
            .in3(N__12228),
            .lcout(un5_visibley_c5),
            .ltout(un5_visibley_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJNLC_9_LC_8_6_3.C_ON=1'b0;
    defparam beamY_RNIJNLC_9_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIJNLC_9_LC_8_6_3.LUT_INIT=16'b1001110111010101;
    LogicCell40 beamY_RNIJNLC_9_LC_8_6_3 (
            .in0(N__13467),
            .in1(N__12080),
            .in2(N__11077),
            .in3(N__12152),
            .lcout(beamY_RNIJNLCZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_RNO_0_LC_8_6_7.C_ON=1'b0;
    defparam VSync_RNO_0_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam VSync_RNO_0_LC_8_6_7.LUT_INIT=16'b0000000000010001;
    LogicCell40 VSync_RNO_0_LC_8_6_7 (
            .in0(N__12538),
            .in1(N__12433),
            .in2(_gnd_net_),
            .in3(N__12153),
            .lcout(un1_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_4_LC_8_7_0.C_ON=1'b0;
    defparam beamY_RNIBFP3_4_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_4_LC_8_7_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 beamY_RNIBFP3_4_LC_8_7_0 (
            .in0(N__12394),
            .in1(N__12529),
            .in2(_gnd_net_),
            .in3(N__12742),
            .lcout(un5_visibley_c3),
            .ltout(un5_visibley_c3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV7J7_7_LC_8_7_1.C_ON=1'b0;
    defparam beamY_RNIV7J7_7_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIV7J7_7_LC_8_7_1.LUT_INIT=16'b1010101010101001;
    LogicCell40 beamY_RNIV7J7_7_LC_8_7_1 (
            .in0(N__12149),
            .in1(N__12223),
            .in2(N__11068),
            .in3(N__12303),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8325_9_LC_8_7_2.C_ON=1'b0;
    defparam beamY_RNI8325_9_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI8325_9_LC_8_7_2.LUT_INIT=16'b0000000010000000;
    LogicCell40 beamY_RNI8325_9_LC_8_7_2 (
            .in0(N__13452),
            .in1(N__12531),
            .in2(N__12434),
            .in3(N__13101),
            .lcout(),
            .ltout(un5_beamx_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_1_LC_8_7_3.C_ON=1'b0;
    defparam beamY_RNI9DLC_1_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_1_LC_8_7_3.LUT_INIT=16'b0100000000000000;
    LogicCell40 beamY_RNI9DLC_1_LC_8_7_3 (
            .in0(N__12743),
            .in1(N__13197),
            .in2(N__11260),
            .in3(N__11257),
            .lcout(beamY_RNI9DLCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8325_0_6_LC_8_7_4.C_ON=1'b0;
    defparam beamY_RNI8325_0_6_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI8325_0_6_LC_8_7_4.LUT_INIT=16'b1100100110011001;
    LogicCell40 beamY_RNI8325_0_6_LC_8_7_4 (
            .in0(N__12304),
            .in1(N__12226),
            .in2(N__12805),
            .in3(N__12530),
            .lcout(beamY_RNI8325_0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIID25_7_LC_8_7_5.C_ON=1'b0;
    defparam beamY_RNIID25_7_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIID25_7_LC_8_7_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_RNIID25_7_LC_8_7_5 (
            .in0(N__12148),
            .in1(N__12222),
            .in2(N__12093),
            .in3(N__12302),
            .lcout(),
            .ltout(un5_visibley_ac0_11_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ7DB_9_LC_8_7_6.C_ON=1'b0;
    defparam beamY_RNIQ7DB_9_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ7DB_9_LC_8_7_6.LUT_INIT=16'b1010011010100101;
    LogicCell40 beamY_RNIQ7DB_9_LC_8_7_6 (
            .in0(N__13451),
            .in1(N__12076),
            .in2(N__11251),
            .in3(N__11895),
            .lcout(chary_if_generate_plus_mult1_un33_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPOR8_0_6_LC_8_7_7.C_ON=1'b0;
    defparam beamY_RNIPOR8_0_6_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIPOR8_0_6_LC_8_7_7.LUT_INIT=16'b1110010010110001;
    LogicCell40 beamY_RNIPOR8_0_6_LC_8_7_7 (
            .in0(N__12405),
            .in1(N__12224),
            .in2(N__11248),
            .in3(N__12305),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_8_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(N__11228),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOU4_LC_8_8_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOU4_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOU4_LC_8_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOU4_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__11426),
            .in2(N__11302),
            .in3(N__11203),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIG7_LC_8_8_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIG7_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIG7_LC_8_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIG7_LC_8_8_2 (
            .in0(_gnd_net_),
            .in1(N__11293),
            .in2(N__11431),
            .in3(N__11194),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5V28_LC_8_8_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5V28_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5V28_LC_8_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5V28_LC_8_8_3 (
            .in0(_gnd_net_),
            .in1(N__11430),
            .in2(N__11284),
            .in3(N__11344),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8PPUJ_LC_8_8_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8PPUJ_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8PPUJ_LC_8_8_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8PPUJ_LC_8_8_4 (
            .in0(N__11327),
            .in1(N__11407),
            .in2(N__11272),
            .in3(N__11335),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37B_LC_8_8_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37B_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37B_LC_8_8_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37B_LC_8_8_5 (
            .in0(_gnd_net_),
            .in1(N__11443),
            .in2(_gnd_net_),
            .in3(N__11332),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_8_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_8_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_8_6 (
            .in0(N__14835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_9_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_9_0 (
            .in0(_gnd_net_),
            .in1(N__14847),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLM2_LC_8_9_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLM2_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLM2_LC_8_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLM2_LC_8_9_1 (
            .in0(_gnd_net_),
            .in1(N__13591),
            .in2(N__11395),
            .in3(N__11287),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJ2193_LC_8_9_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJ2193_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJ2193_LC_8_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJ2193_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__13594),
            .in2(N__13675),
            .in3(N__11275),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NT3_LC_8_9_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NT3_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NT3_LC_8_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NT3_LC_8_9_3 (
            .in0(_gnd_net_),
            .in1(N__13592),
            .in2(N__13654),
            .in3(N__11263),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNITBNTA_LC_8_9_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNITBNTA_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNITBNTA_LC_8_9_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNITBNTA_LC_8_9_4 (
            .in0(N__11425),
            .in1(N__11401),
            .in2(N__13636),
            .in3(N__11437),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_LC_8_9_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_LC_8_9_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_LC_8_9_5 (
            .in0(_gnd_net_),
            .in1(N__13612),
            .in2(_gnd_net_),
            .in3(N__11434),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_0_LC_8_9_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_0_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_0_LC_8_9_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_0_LC_8_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11410),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJ54_LC_8_9_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJ54_LC_8_9_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJ54_LC_8_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJ54_LC_8_9_7 (
            .in0(_gnd_net_),
            .in1(N__13635),
            .in2(_gnd_net_),
            .in3(N__13590),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_10_0.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14769),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN49K_8_LC_8_10_1.C_ON=1'b0;
    defparam beamY_RNIN49K_8_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIN49K_8_LC_8_10_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_RNIN49K_8_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__15123),
            .in2(_gnd_net_),
            .in3(N__15188),
            .lcout(CO4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un47_sum_c5_LC_8_10_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un47_sum_c5_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un47_sum_c5_LC_8_10_4.LUT_INIT=16'b0101101000001010;
    LogicCell40 row_1_if_generate_plus_mult1_un47_sum_c5_LC_8_10_4 (
            .in0(N__15189),
            .in1(_gnd_net_),
            .in2(N__15127),
            .in3(N__15718),
            .lcout(row_1_if_generate_plus_mult1_un47_sum_cZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram8__e_0_0_LC_8_11_2.C_ON=1'b0;
    defparam content_content_ram8__e_0_0_LC_8_11_2.SEQ_MODE=4'b1000;
    defparam content_content_ram8__e_0_0_LC_8_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 content_content_ram8__e_0_0_LC_8_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14538),
            .lcout(content_ram8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14341),
            .ce(N__11482),
            .sr(_gnd_net_));
    defparam content_content_ram10__e_0_RNIOLNMN1_0_0_LC_8_11_3.C_ON=1'b0;
    defparam content_content_ram10__e_0_RNIOLNMN1_0_0_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam content_content_ram10__e_0_RNIOLNMN1_0_0_LC_8_11_3.LUT_INIT=16'b1010100000001000;
    LogicCell40 content_content_ram10__e_0_RNIOLNMN1_0_0_LC_8_11_3 (
            .in0(N__11658),
            .in1(N__13828),
            .in2(N__11599),
            .in3(N__13797),
            .lcout(),
            .ltout(content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram6__RNI1FLOF3_0_LC_8_11_4.C_ON=1'b0;
    defparam content_content_ram6__RNI1FLOF3_0_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam content_content_ram6__RNI1FLOF3_0_LC_8_11_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 content_content_ram6__RNI1FLOF3_0_LC_8_11_4 (
            .in0(_gnd_net_),
            .in1(N__11743),
            .in2(N__11695),
            .in3(N__11533),
            .lcout(content_N_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram10__e_0_RNIOLNMN1_0_LC_8_11_5.C_ON=1'b0;
    defparam content_content_ram10__e_0_RNIOLNMN1_0_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam content_content_ram10__e_0_RNIOLNMN1_0_LC_8_11_5.LUT_INIT=16'b1111100001011000;
    LogicCell40 content_content_ram10__e_0_RNIOLNMN1_0_LC_8_11_5 (
            .in0(N__11657),
            .in1(N__13827),
            .in2(N__11598),
            .in3(N__13796),
            .lcout(content_content_ram10__e_0_RNIOLNMN1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram3__0_LC_8_12_1.C_ON=1'b0;
    defparam content_content_ram3__0_LC_8_12_1.SEQ_MODE=4'b1000;
    defparam content_content_ram3__0_LC_8_12_1.LUT_INIT=16'b1111000010111000;
    LogicCell40 content_content_ram3__0_LC_8_12_1 (
            .in0(N__14541),
            .in1(N__13807),
            .in2(N__11527),
            .in3(N__14047),
            .lcout(content_ram3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14342),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram9__e_0_RNO_0_LC_8_12_2.C_ON=1'b0;
    defparam content_content_ram9__e_0_RNO_0_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam content_content_ram9__e_0_RNO_0_LC_8_12_2.LUT_INIT=16'b1000000000001000;
    LogicCell40 content_content_ram9__e_0_RNO_0_LC_8_12_2 (
            .in0(N__13782),
            .in1(N__13757),
            .in2(N__13918),
            .in3(N__14173),
            .lcout(content_awe9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram0__0_LC_8_12_4.C_ON=1'b0;
    defparam content_content_ram0__0_LC_8_12_4.SEQ_MODE=4'b1000;
    defparam content_content_ram0__0_LC_8_12_4.LUT_INIT=16'b1111100001110000;
    LogicCell40 content_content_ram0__0_LC_8_12_4 (
            .in0(N__11788),
            .in1(N__13758),
            .in2(N__11500),
            .in3(N__14540),
            .lcout(content_ram0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14342),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram8__e_0_RNO_0_LC_8_12_5.C_ON=1'b0;
    defparam content_content_ram8__e_0_RNO_0_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam content_content_ram8__e_0_RNO_0_LC_8_12_5.LUT_INIT=16'b0000000001000000;
    LogicCell40 content_content_ram8__e_0_RNO_0_LC_8_12_5 (
            .in0(N__13698),
            .in1(N__14045),
            .in2(N__13763),
            .in3(N__14111),
            .lcout(content_awe8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram11__e_0_RNO_0_LC_8_12_7.C_ON=1'b0;
    defparam content_content_ram11__e_0_RNO_0_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam content_content_ram11__e_0_RNO_0_LC_8_12_7.LUT_INIT=16'b0000000000010000;
    LogicCell40 content_content_ram11__e_0_RNO_0_LC_8_12_7 (
            .in0(N__13697),
            .in1(N__14046),
            .in2(N__13764),
            .in3(N__14112),
            .lcout(content_awe11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram5__0_LC_8_13_0.C_ON=1'b0;
    defparam content_content_ram5__0_LC_8_13_0.SEQ_MODE=4'b1000;
    defparam content_content_ram5__0_LC_8_13_0.LUT_INIT=16'b1111100001110000;
    LogicCell40 content_content_ram5__0_LC_8_13_0 (
            .in0(N__11760),
            .in1(N__13783),
            .in2(N__11461),
            .in3(N__14537),
            .lcout(content_ram5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14345),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_0_LC_8_13_1.C_ON=1'b0;
    defparam counter_0_LC_8_13_1.SEQ_MODE=4'b1000;
    defparam counter_0_LC_8_13_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 counter_0_LC_8_13_1 (
            .in0(_gnd_net_),
            .in1(N__14608),
            .in2(_gnd_net_),
            .in3(N__14044),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14345),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1_LC_8_13_3.C_ON=1'b0;
    defparam counter_1_LC_8_13_3.SEQ_MODE=4'b1000;
    defparam counter_1_LC_8_13_3.LUT_INIT=16'b0110011000000000;
    LogicCell40 counter_1_LC_8_13_3 (
            .in0(N__14116),
            .in1(N__14043),
            .in2(_gnd_net_),
            .in3(N__14609),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14345),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram12__0_LC_8_13_4.C_ON=1'b0;
    defparam content_content_ram12__0_LC_8_13_4.SEQ_MODE=4'b1000;
    defparam content_content_ram12__0_LC_8_13_4.LUT_INIT=16'b1111001011010000;
    LogicCell40 content_content_ram12__0_LC_8_13_4 (
            .in0(N__11761),
            .in1(N__13699),
            .in2(N__11808),
            .in3(N__14535),
            .lcout(content_ram12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14345),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNINMOJ_3_LC_8_13_5.C_ON=1'b0;
    defparam counter_RNINMOJ_3_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam counter_RNINMOJ_3_LC_8_13_5.LUT_INIT=16'b0001000000100000;
    LogicCell40 counter_RNINMOJ_3_LC_8_13_5 (
            .in0(N__14171),
            .in1(N__14110),
            .in2(N__14059),
            .in3(N__13903),
            .lcout(content_awe0_0_a2_0),
            .ltout(content_awe0_0_a2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram4__0_LC_8_13_6.C_ON=1'b0;
    defparam content_content_ram4__0_LC_8_13_6.SEQ_MODE=4'b1000;
    defparam content_content_ram4__0_LC_8_13_6.LUT_INIT=16'b1101111110000000;
    LogicCell40 content_content_ram4__0_LC_8_13_6 (
            .in0(N__11759),
            .in1(N__14536),
            .in2(N__11782),
            .in3(N__11775),
            .lcout(content_ram4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14345),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIHRI6_1_LC_8_13_7.C_ON=1'b0;
    defparam counter_RNIHRI6_1_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam counter_RNIHRI6_1_LC_8_13_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 counter_RNIHRI6_1_LC_8_13_7 (
            .in0(_gnd_net_),
            .in1(N__14042),
            .in2(_gnd_net_),
            .in3(N__14109),
            .lcout(content_N_40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIVRML1_2_LC_8_14_0.C_ON=1'b0;
    defparam counter_RNIVRML1_2_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam counter_RNIVRML1_2_LC_8_14_0.LUT_INIT=16'b1000000001000000;
    LogicCell40 counter_RNIVRML1_2_LC_8_14_0 (
            .in0(N__13973),
            .in1(N__14433),
            .in2(N__14395),
            .in3(N__13955),
            .lcout(content_N_36),
            .ltout(content_N_36_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIGN9S1_1_LC_8_14_1.C_ON=1'b0;
    defparam counter_RNIGN9S1_1_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam counter_RNIGN9S1_1_LC_8_14_1.LUT_INIT=16'b1100000000110000;
    LogicCell40 counter_RNIGN9S1_1_LC_8_14_1 (
            .in0(_gnd_net_),
            .in1(N__14115),
            .in2(N__11749),
            .in3(N__14053),
            .lcout(content_awe7_1),
            .ltout(content_awe7_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram6__0_LC_8_14_2.C_ON=1'b0;
    defparam content_content_ram6__0_LC_8_14_2.SEQ_MODE=4'b1000;
    defparam content_content_ram6__0_LC_8_14_2.LUT_INIT=16'b1101111110000000;
    LogicCell40 content_content_ram6__0_LC_8_14_2 (
            .in0(N__14054),
            .in1(N__14530),
            .in2(N__11746),
            .in3(N__11742),
            .lcout(content_ram6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14347),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram7__0_LC_8_14_3.C_ON=1'b0;
    defparam content_content_ram7__0_LC_8_14_3.SEQ_MODE=4'b1000;
    defparam content_content_ram7__0_LC_8_14_3.LUT_INIT=16'b1111000010111000;
    LogicCell40 content_content_ram7__0_LC_8_14_3 (
            .in0(N__14531),
            .in1(N__11728),
            .in2(N__11722),
            .in3(N__14055),
            .lcout(content_ram7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14347),
            .ce(),
            .sr(_gnd_net_));
    defparam nCS1_1_RNO_0_LC_8_14_4.C_ON=1'b0;
    defparam nCS1_1_RNO_0_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam nCS1_1_RNO_0_LC_8_14_4.LUT_INIT=16'b1110111000000000;
    LogicCell40 nCS1_1_RNO_0_LC_8_14_4 (
            .in0(N__14571),
            .in1(N__11880),
            .in2(_gnd_net_),
            .in3(N__14434),
            .lcout(nCS1_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIICFG_4_LC_8_14_5.C_ON=1'b0;
    defparam counter_RNIICFG_4_LC_8_14_5.SEQ_MODE=4'b0000;
    defparam counter_RNIICFG_4_LC_8_14_5.LUT_INIT=16'b1100100011001100;
    LogicCell40 counter_RNIICFG_4_LC_8_14_5 (
            .in0(N__13954),
            .in1(N__13851),
            .in2(N__13917),
            .in3(N__13974),
            .lcout(un19_slaveselectlt5_0),
            .ltout(un19_slaveselectlt5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI4HQB1_5_LC_8_14_6.C_ON=1'b0;
    defparam counter_RNI4HQB1_5_LC_8_14_6.SEQ_MODE=4'b0000;
    defparam counter_RNI4HQB1_5_LC_8_14_6.LUT_INIT=16'b0000010101110111;
    LogicCell40 counter_RNI4HQB1_5_LC_8_14_6 (
            .in0(N__14572),
            .in1(N__14184),
            .in2(N__11884),
            .in3(N__14435),
            .lcout(counter_RNI4HQB1Z0Z_5),
            .ltout(counter_RNI4HQB1Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_LC_8_14_7.C_ON=1'b0;
    defparam slaveselect_LC_8_14_7.SEQ_MODE=4'b1000;
    defparam slaveselect_LC_8_14_7.LUT_INIT=16'b0001000100001111;
    LogicCell40 slaveselect_LC_8_14_7 (
            .in0(N__11881),
            .in1(N__14573),
            .in2(N__11872),
            .in3(N__14440),
            .lcout(slaveselectZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14347),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4FVGV_4_LC_9_4_5.C_ON=1'b0;
    defparam beamY_RNI4FVGV_4_LC_9_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI4FVGV_4_LC_9_4_5.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI4FVGV_4_LC_9_4_5 (
            .in0(N__14967),
            .in1(N__14280),
            .in2(_gnd_net_),
            .in3(N__12437),
            .lcout(),
            .ltout(beamY_RNI4FVGVZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7LOHP1_3_LC_9_4_6.C_ON=1'b0;
    defparam beamY_RNI7LOHP1_3_LC_9_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI7LOHP1_3_LC_9_4_6.LUT_INIT=16'b0000110100111101;
    LogicCell40 beamY_RNI7LOHP1_3_LC_9_4_6 (
            .in0(N__14302),
            .in1(N__12599),
            .in2(N__11869),
            .in3(N__12856),
            .lcout(chary_if_generate_plus_mult1_un75_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_90_LC_9_5_0.C_ON=1'b0;
    defparam Pixel_RNO_90_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_90_LC_9_5_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 Pixel_RNO_90_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__12637),
            .in2(_gnd_net_),
            .in3(N__12859),
            .lcout(un5_visibley_3_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_49_LC_9_5_1.C_ON=1'b0;
    defparam Pixel_RNO_49_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_49_LC_9_5_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 Pixel_RNO_49_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__13075),
            .in2(_gnd_net_),
            .in3(N__13252),
            .lcout(N_596_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_93_LC_9_5_3.C_ON=1'b0;
    defparam Pixel_RNO_93_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_93_LC_9_5_3.LUT_INIT=16'b0101111110100000;
    LogicCell40 Pixel_RNO_93_LC_9_5_3 (
            .in0(N__12861),
            .in1(_gnd_net_),
            .in2(N__12669),
            .in3(N__12440),
            .lcout(),
            .ltout(un5_visibley_4_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_89_LC_9_5_4.C_ON=1'b0;
    defparam Pixel_RNO_89_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_89_LC_9_5_4.LUT_INIT=16'b0011010011000001;
    LogicCell40 Pixel_RNO_89_LC_9_5_4 (
            .in0(N__14704),
            .in1(N__14966),
            .in2(N__11815),
            .in3(N__14274),
            .lcout(),
            .ltout(g1_8_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_83_LC_9_5_5.C_ON=1'b0;
    defparam Pixel_RNO_83_LC_9_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_83_LC_9_5_5.LUT_INIT=16'b0000110010101100;
    LogicCell40 Pixel_RNO_83_LC_9_5_5 (
            .in0(N__12028),
            .in1(N__14705),
            .in2(N__12022),
            .in3(N__11992),
            .lcout(g1_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_94_LC_9_5_6.C_ON=1'b0;
    defparam Pixel_RNO_94_LC_9_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_94_LC_9_5_6.LUT_INIT=16'b0110011010101010;
    LogicCell40 Pixel_RNO_94_LC_9_5_6 (
            .in0(N__12439),
            .in1(N__12638),
            .in2(_gnd_net_),
            .in3(N__12860),
            .lcout(un5_visibley_1_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_0_4_LC_9_6_0.C_ON=1'b0;
    defparam beamY_RNIBFP3_0_4_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_0_4_LC_9_6_0.LUT_INIT=16'b0111100001111000;
    LogicCell40 beamY_RNIBFP3_0_4_LC_9_6_0 (
            .in0(N__12534),
            .in1(N__12746),
            .in2(N__12436),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_5_LC_9_6_2.C_ON=1'b0;
    defparam beamY_RNI6125_5_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_5_LC_9_6_2.LUT_INIT=16'b1000000001111111;
    LogicCell40 beamY_RNI6125_5_LC_9_6_2 (
            .in0(N__12533),
            .in1(N__12745),
            .in2(N__12435),
            .in3(N__12307),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0H2_4_LC_9_6_3.C_ON=1'b0;
    defparam beamY_RNIJ0H2_4_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0H2_4_LC_9_6_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_RNIJ0H2_4_LC_9_6_3 (
            .in0(_gnd_net_),
            .in1(N__12398),
            .in2(_gnd_net_),
            .in3(N__12532),
            .lcout(),
            .ltout(beamY_RNIJ0H2Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITSR8_8_LC_9_6_4.C_ON=1'b0;
    defparam beamY_RNITSR8_8_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNITSR8_8_LC_9_6_4.LUT_INIT=16'b1010101010010101;
    LogicCell40 beamY_RNITSR8_8_LC_9_6_4 (
            .in0(N__12078),
            .in1(N__12744),
            .in2(N__11917),
            .in3(N__11905),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJNLC_0_9_LC_9_6_5.C_ON=1'b0;
    defparam beamY_RNIJNLC_0_9_LC_9_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIJNLC_0_9_LC_9_6_5.LUT_INIT=16'b1001001000100101;
    LogicCell40 beamY_RNIJNLC_0_9_LC_9_6_5 (
            .in0(N__13468),
            .in1(N__12079),
            .in2(N__11914),
            .in3(N__12151),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKOP3_7_LC_9_6_6.C_ON=1'b0;
    defparam beamY_RNIKOP3_7_LC_9_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIKOP3_7_LC_9_6_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamY_RNIKOP3_7_LC_9_6_6 (
            .in0(N__12150),
            .in1(N__12225),
            .in2(_gnd_net_),
            .in3(N__12306),
            .lcout(un5_visibley_c6_0_0_0),
            .ltout(un5_visibley_c6_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_9_6_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_9_6_7.LUT_INIT=16'b1100110011000011;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_9_6_7 (
            .in0(_gnd_net_),
            .in1(N__12077),
            .in2(N__11899),
            .in3(N__11896),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_47_LC_9_7_0.C_ON=1'b1;
    defparam Pixel_RNO_47_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_47_LC_9_7_0.LUT_INIT=16'b1001100110011001;
    LogicCell40 Pixel_RNO_47_LC_9_7_0 (
            .in0(N__13076),
            .in1(N__13201),
            .in2(N__13105),
            .in3(_gnd_net_),
            .lcout(g2_1_1_0),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_9_7_1.C_ON=1'b1;
    defparam beamY_2_LC_9_7_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_9_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_2_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(N__12804),
            .in2(_gnd_net_),
            .in3(N__12676),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_3_LC_9_7_2.C_ON=1'b1;
    defparam beamY_3_LC_9_7_2.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_9_7_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_3_LC_9_7_2 (
            .in0(N__13529),
            .in1(N__12585),
            .in2(_gnd_net_),
            .in3(N__12463),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_4_LC_9_7_3.C_ON=1'b1;
    defparam beamY_4_LC_9_7_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_9_7_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_4_LC_9_7_3 (
            .in0(N__13518),
            .in1(N__12432),
            .in2(_gnd_net_),
            .in3(N__12331),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_5_LC_9_7_4.C_ON=1'b1;
    defparam beamY_5_LC_9_7_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_9_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__12256),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_6_LC_9_7_5.C_ON=1'b1;
    defparam beamY_6_LC_9_7_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_9_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(N__12240),
            .in2(_gnd_net_),
            .in3(N__12175),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_7_LC_9_7_6.C_ON=1'b1;
    defparam beamY_7_LC_9_7_6.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_9_7_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_7_LC_9_7_6 (
            .in0(N__13530),
            .in1(N__12163),
            .in2(_gnd_net_),
            .in3(N__12109),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_8_LC_9_7_7.C_ON=1'b1;
    defparam beamY_8_LC_9_7_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_9_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(N__12092),
            .in2(_gnd_net_),
            .in3(N__12031),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(N__13426),
            .ce(N__13392),
            .sr(_gnd_net_));
    defparam beamY_9_LC_9_8_0.C_ON=1'b0;
    defparam beamY_9_LC_9_8_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_9_8_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_9_8_0 (
            .in0(N__13466),
            .in1(N__13519),
            .in2(_gnd_net_),
            .in3(N__13489),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13424),
            .ce(N__13393),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_9_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(N__15273),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_9_9_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_9_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(N__13303),
            .in2(N__15417),
            .in3(N__13324),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBC41_LC_9_9_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBC41_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBC41_LC_9_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBC41_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__15412),
            .in2(N__15649),
            .in3(N__13321),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEG81_LC_9_9_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEG81_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEG81_LC_9_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEG81_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(N__15625),
            .in2(N__15418),
            .in3(N__13318),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIFFA42_LC_9_9_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIFFA42_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIFFA42_LC_9_9_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIFFA42_LC_9_9_4 (
            .in0(N__13568),
            .in1(N__13309),
            .in2(N__15451),
            .in3(N__13315),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_9_9_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_9_9_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_9_9_5 (
            .in0(N__15416),
            .in1(N__15382),
            .in2(N__15436),
            .in3(N__13312),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_9_9_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_9_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15408),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_9_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_9_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15704),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_10_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(N__14747),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_9_10_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_9_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(N__13537),
            .in2(N__13569),
            .in3(N__13666),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_9_10_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_9_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_9_10_2 (
            .in0(_gnd_net_),
            .in1(N__13564),
            .in2(N__13663),
            .in3(N__13645),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4L02_LC_9_10_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4L02_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4L02_LC_9_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4L02_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(N__13642),
            .in2(N__13570),
            .in3(N__13624),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNISRO94_LC_9_10_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNISRO94_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNISRO94_LC_9_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNISRO94_LC_9_10_4 (
            .in0(N__13593),
            .in1(N__13543),
            .in2(N__13621),
            .in3(N__13606),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IU42_LC_9_10_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IU42_LC_9_10_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IU42_LC_9_10_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IU42_LC_9_10_5 (
            .in0(_gnd_net_),
            .in1(N__13603),
            .in2(_gnd_net_),
            .in3(N__13597),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_9_10_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_9_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13560),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_10_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_10_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_10_7 (
            .in0(N__15274),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram10__e_0_0_LC_9_11_0.C_ON=1'b0;
    defparam content_content_ram10__e_0_0_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam content_content_ram10__e_0_0_LC_9_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 content_content_ram10__e_0_0_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14534),
            .lcout(content_ram10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14343),
            .ce(N__13819),
            .sr(_gnd_net_));
    defparam content_content_ram10__e_0_RNO_0_LC_9_12_0.C_ON=1'b0;
    defparam content_content_ram10__e_0_RNO_0_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam content_content_ram10__e_0_RNO_0_LC_9_12_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 content_content_ram10__e_0_RNO_0_LC_9_12_0 (
            .in0(N__14113),
            .in1(N__13696),
            .in2(N__13765),
            .in3(N__14048),
            .lcout(content_awe10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIVRML1_0_2_LC_9_12_2.C_ON=1'b0;
    defparam counter_RNIVRML1_0_2_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam counter_RNIVRML1_0_2_LC_9_12_2.LUT_INIT=16'b0100100000000000;
    LogicCell40 counter_RNIVRML1_0_2_LC_9_12_2 (
            .in0(N__13978),
            .in1(N__14442),
            .in2(N__13960),
            .in3(N__14390),
            .lcout(content_N_35),
            .ltout(content_N_35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIMIF92_1_LC_9_12_3.C_ON=1'b0;
    defparam counter_RNIMIF92_1_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam counter_RNIMIF92_1_LC_9_12_3.LUT_INIT=16'b1000000000100000;
    LogicCell40 counter_RNIMIF92_1_LC_9_12_3 (
            .in0(N__13695),
            .in1(N__14056),
            .in2(N__13810),
            .in3(N__14114),
            .lcout(content_awe3_1),
            .ltout(content_awe3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram2__0_LC_9_12_4.C_ON=1'b0;
    defparam content_content_ram2__0_LC_9_12_4.SEQ_MODE=4'b1000;
    defparam content_content_ram2__0_LC_9_12_4.LUT_INIT=16'b1011111110000000;
    LogicCell40 content_content_ram2__0_LC_9_12_4 (
            .in0(N__14533),
            .in1(N__14049),
            .in2(N__13801),
            .in3(N__13798),
            .lcout(content_ram2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14346),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram1__RNO_0_0_LC_9_12_5.C_ON=1'b0;
    defparam content_content_ram1__RNO_0_0_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam content_content_ram1__RNO_0_0_LC_9_12_5.LUT_INIT=16'b0110011000000000;
    LogicCell40 content_content_ram1__RNO_0_0_LC_9_12_5 (
            .in0(N__13915),
            .in1(N__14172),
            .in2(_gnd_net_),
            .in3(N__13781),
            .lcout(),
            .ltout(content_awe1_0_a2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam content_content_ram1__0_LC_9_12_6.C_ON=1'b0;
    defparam content_content_ram1__0_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam content_content_ram1__0_LC_9_12_6.LUT_INIT=16'b1011111110000000;
    LogicCell40 content_content_ram1__0_LC_9_12_6 (
            .in0(N__14532),
            .in1(N__13762),
            .in2(N__13729),
            .in3(N__13716),
            .lcout(content_ram1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14346),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIRAS9_2_LC_9_13_0.C_ON=1'b0;
    defparam counter_RNIRAS9_2_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam counter_RNIRAS9_2_LC_9_13_0.LUT_INIT=16'b1100100011001000;
    LogicCell40 counter_RNIRAS9_2_LC_9_13_0 (
            .in0(N__14105),
            .in1(N__13948),
            .in2(N__14058),
            .in3(_gnd_net_),
            .lcout(un7_slaveselectlt5),
            .ltout(un7_slaveselectlt5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_3_LC_9_13_1.C_ON=1'b0;
    defparam counter_RNI6R5D_3_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_3_LC_9_13_1.LUT_INIT=16'b0000111111110000;
    LogicCell40 counter_RNI6R5D_3_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13702),
            .in3(N__13908),
            .lcout(N_190_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIN1J6_4_LC_9_13_2.C_ON=1'b0;
    defparam counter_RNIN1J6_4_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam counter_RNIN1J6_4_LC_9_13_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_RNIN1J6_4_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(N__13849),
            .in2(_gnd_net_),
            .in3(N__13888),
            .lcout(slaveselect_1lto5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIAV5D_4_LC_9_13_4.C_ON=1'b0;
    defparam counter_RNIAV5D_4_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam counter_RNIAV5D_4_LC_9_13_4.LUT_INIT=16'b1111111000000000;
    LogicCell40 counter_RNIAV5D_4_LC_9_13_4 (
            .in0(N__14106),
            .in1(N__13949),
            .in2(N__13916),
            .in3(N__13850),
            .lcout(un1_counter_0_1),
            .ltout(un1_counter_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI9UU01_5_LC_9_13_5.C_ON=1'b0;
    defparam counter_RNI9UU01_5_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam counter_RNI9UU01_5_LC_9_13_5.LUT_INIT=16'b0000010000000101;
    LogicCell40 counter_RNI9UU01_5_LC_9_13_5 (
            .in0(N__14569),
            .in1(N__14170),
            .in2(N__14149),
            .in3(N__14142),
            .lcout(un5_slaveselect),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI0GS9_5_LC_9_13_6.C_ON=1'b0;
    defparam counter_RNI0GS9_5_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam counter_RNI0GS9_5_LC_9_13_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 counter_RNI0GS9_5_LC_9_13_6 (
            .in0(N__14107),
            .in1(N__13950),
            .in2(_gnd_net_),
            .in3(N__14570),
            .lcout(),
            .ltout(slaveselect_1lto5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNIK7MV_LC_9_13_7.C_ON=1'b0;
    defparam slaveselect_RNIK7MV_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam slaveselect_RNIK7MV_LC_9_13_7.LUT_INIT=16'b1111110111011101;
    LogicCell40 slaveselect_RNIK7MV_LC_9_13_7 (
            .in0(N__14441),
            .in1(N__14359),
            .in2(N__14146),
            .in3(N__14143),
            .lcout(SCLK1_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIHRI6_0_1_LC_9_14_0.C_ON=1'b1;
    defparam counter_RNIHRI6_0_1_LC_9_14_0.SEQ_MODE=4'b0000;
    defparam counter_RNIHRI6_0_1_LC_9_14_0.LUT_INIT=16'b0001000100010001;
    LogicCell40 counter_RNIHRI6_0_1_LC_9_14_0 (
            .in0(N__14035),
            .in1(N__14108),
            .in2(N__14057),
            .in3(_gnd_net_),
            .lcout(un7_slaveselectlt2_0),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_9_14_1.C_ON=1'b1;
    defparam counter_2_LC_9_14_1.SEQ_MODE=4'b1000;
    defparam counter_2_LC_9_14_1.LUT_INIT=16'b0010001010001000;
    LogicCell40 counter_2_LC_9_14_1 (
            .in0(N__14610),
            .in1(N__13956),
            .in2(_gnd_net_),
            .in3(N__13921),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(counter_cry_1),
            .carryout(counter_cry_2),
            .clk(N__14351),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_3_LC_9_14_2.C_ON=1'b1;
    defparam counter_3_LC_9_14_2.SEQ_MODE=4'b1000;
    defparam counter_3_LC_9_14_2.LUT_INIT=16'b0010001010001000;
    LogicCell40 counter_3_LC_9_14_2 (
            .in0(N__14606),
            .in1(N__13904),
            .in2(_gnd_net_),
            .in3(N__13855),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(counter_cry_2),
            .carryout(counter_cry_3),
            .clk(N__14351),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_4_LC_9_14_3.C_ON=1'b1;
    defparam counter_4_LC_9_14_3.SEQ_MODE=4'b1000;
    defparam counter_4_LC_9_14_3.LUT_INIT=16'b0010001010001000;
    LogicCell40 counter_4_LC_9_14_3 (
            .in0(N__14611),
            .in1(N__13852),
            .in2(_gnd_net_),
            .in3(N__13831),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(counter_cry_3),
            .carryout(counter_cry_4),
            .clk(N__14351),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_5_LC_9_14_4.C_ON=1'b0;
    defparam counter_5_LC_9_14_4.SEQ_MODE=4'b1000;
    defparam counter_5_LC_9_14_4.LUT_INIT=16'b0010001010001000;
    LogicCell40 counter_5_LC_9_14_4 (
            .in0(N__14607),
            .in1(N__14577),
            .in2(_gnd_net_),
            .in3(N__14584),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14351),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATAZ0Z2_LC_9_14_6.C_ON=1'b0;
    defparam SDATAZ0Z2_LC_9_14_6.SEQ_MODE=4'b1000;
    defparam SDATAZ0Z2_LC_9_14_6.LUT_INIT=16'b1100101000001010;
    LogicCell40 SDATAZ0Z2_LC_9_14_6 (
            .in0(N__14370),
            .in1(N__14521),
            .in2(N__14443),
            .in3(N__14394),
            .lcout(SDATA2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14351),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUR98A_9_LC_11_5_0.C_ON=1'b0;
    defparam beamY_RNIUR98A_9_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIUR98A_9_LC_11_5_0.LUT_INIT=16'b0110011001100110;
    LogicCell40 beamY_RNIUR98A_9_LC_11_5_0 (
            .in0(N__14650),
            .in1(N__14875),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII78UP_4_LC_11_5_1.C_ON=1'b0;
    defparam beamY_RNII78UP_4_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNII78UP_4_LC_11_5_1.LUT_INIT=16'b0110001111000110;
    LogicCell40 beamY_RNII78UP_4_LC_11_5_1 (
            .in0(N__14785),
            .in1(N__14202),
            .in2(N__14305),
            .in3(N__14850),
            .lcout(beamY_RNII78UPZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5VO45_6_LC_11_5_2.C_ON=1'b0;
    defparam beamY_RNI5VO45_6_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI5VO45_6_LC_11_5_2.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI5VO45_6_LC_11_5_2 (
            .in0(N__15342),
            .in1(N__14782),
            .in2(_gnd_net_),
            .in3(N__15293),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI3R2DF_6_LC_11_5_3.C_ON=1'b0;
    defparam beamY_RNI3R2DF_6_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI3R2DF_6_LC_11_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamY_RNI3R2DF_6_LC_11_5_3 (
            .in0(_gnd_net_),
            .in1(N__14873),
            .in2(N__14290),
            .in3(N__14646),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFC5HA_1_4_LC_11_5_4.C_ON=1'b0;
    defparam beamY_RNIFC5HA_1_4_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIFC5HA_1_4_LC_11_5_4.LUT_INIT=16'b0001010001111101;
    LogicCell40 beamY_RNIFC5HA_1_4_LC_11_5_4 (
            .in0(N__14848),
            .in1(N__14874),
            .in2(N__14653),
            .in3(N__14783),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKBULF_6_LC_11_5_5.C_ON=1'b0;
    defparam beamY_RNIKBULF_6_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIKBULF_6_LC_11_5_5.LUT_INIT=16'b0010011100011011;
    LogicCell40 beamY_RNIKBULF_6_LC_11_5_5 (
            .in0(N__15294),
            .in1(N__14786),
            .in2(N__14287),
            .in3(N__15343),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c5),
            .ltout(chary_if_generate_plus_mult1_un61_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIS5VDP1_4_LC_11_5_6.C_ON=1'b0;
    defparam beamY_RNIS5VDP1_4_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIS5VDP1_4_LC_11_5_6.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIS5VDP1_4_LC_11_5_6 (
            .in0(N__14203),
            .in1(N__15013),
            .in2(N__14194),
            .in3(N__14917),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFC5HA_0_4_LC_11_5_7.C_ON=1'b0;
    defparam beamY_RNIFC5HA_0_4_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIFC5HA_0_4_LC_11_5_7.LUT_INIT=16'b0100110111010100;
    LogicCell40 beamY_RNIFC5HA_0_4_LC_11_5_7 (
            .in0(N__14784),
            .in1(N__14849),
            .in2(N__14881),
            .in3(N__14651),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIOMEH5_0_9_LC_11_6_1.C_ON=1'b0;
    defparam beamY_RNIOMEH5_0_9_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIOMEH5_0_9_LC_11_6_1.LUT_INIT=16'b0000110111110100;
    LogicCell40 beamY_RNIOMEH5_0_9_LC_11_6_1 (
            .in0(N__15335),
            .in1(N__14787),
            .in2(N__15006),
            .in3(N__15291),
            .lcout(chary_if_generate_plus_mult1_un54_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIOMEH5_9_LC_11_6_3.C_ON=1'b0;
    defparam beamY_RNIOMEH5_9_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIOMEH5_9_LC_11_6_3.LUT_INIT=16'b1101001001001011;
    LogicCell40 beamY_RNIOMEH5_9_LC_11_6_3 (
            .in0(N__15336),
            .in1(N__14788),
            .in2(N__15007),
            .in3(N__15292),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMIOPF_9_LC_11_6_4.C_ON=1'b0;
    defparam beamY_RNIMIOPF_9_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIMIOPF_9_LC_11_6_4.LUT_INIT=16'b0011110011000011;
    LogicCell40 beamY_RNIMIOPF_9_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(N__14642),
            .in2(N__14989),
            .in3(N__14879),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFC5HA_4_LC_11_6_7.C_ON=1'b0;
    defparam beamY_RNIFC5HA_4_LC_11_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIFC5HA_4_LC_11_6_7.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIFC5HA_4_LC_11_6_7 (
            .in0(N__14880),
            .in1(N__14851),
            .in2(N__14652),
            .in3(N__14789),
            .lcout(beamY_RNIFC5HAZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI94I81_9_LC_11_7_0.C_ON=1'b0;
    defparam beamY_RNI94I81_9_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI94I81_9_LC_11_7_0.LUT_INIT=16'b1001011011000011;
    LogicCell40 beamY_RNI94I81_9_LC_11_7_0 (
            .in0(N__15180),
            .in1(N__15706),
            .in2(N__15322),
            .in3(N__15114),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axb4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI94I81_0_9_LC_11_7_1.C_ON=1'b0;
    defparam beamY_RNI94I81_0_9_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI94I81_0_9_LC_11_7_1.LUT_INIT=16'b1010011101011000;
    LogicCell40 beamY_RNI94I81_0_9_LC_11_7_1 (
            .in0(N__15115),
            .in1(N__15708),
            .in2(N__15192),
            .in3(N__15319),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axbxc5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI65RM4_9_LC_11_7_3.C_ON=1'b0;
    defparam beamY_RNI65RM4_9_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI65RM4_9_LC_11_7_3.LUT_INIT=16'b1001110001101001;
    LogicCell40 beamY_RNI65RM4_9_LC_11_7_3 (
            .in0(N__15223),
            .in1(N__15364),
            .in2(N__14620),
            .in3(N__15352),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI94I81_1_9_LC_11_7_4.C_ON=1'b0;
    defparam beamY_RNI94I81_1_9_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI94I81_1_9_LC_11_7_4.LUT_INIT=16'b0000100100001100;
    LogicCell40 beamY_RNI94I81_1_9_LC_11_7_4 (
            .in0(N__15181),
            .in1(N__15705),
            .in2(N__15321),
            .in3(N__15113),
            .lcout(chary_if_generate_plus_mult1_un47_sum_ac0_8),
            .ltout(chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI65RM4_0_9_LC_11_7_5.C_ON=1'b0;
    defparam beamY_RNI65RM4_0_9_LC_11_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI65RM4_0_9_LC_11_7_5.LUT_INIT=16'b0011011000111100;
    LogicCell40 beamY_RNI65RM4_0_9_LC_11_7_5 (
            .in0(N__15222),
            .in1(N__15363),
            .in2(N__15355),
            .in3(N__15351),
            .lcout(beamY_RNI65RM4_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBO4T_9_LC_11_7_6.C_ON=1'b0;
    defparam beamY_RNIBO4T_9_LC_11_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIBO4T_9_LC_11_7_6.LUT_INIT=16'b1000100011101110;
    LogicCell40 beamY_RNIBO4T_9_LC_11_7_6 (
            .in0(N__15320),
            .in1(N__15280),
            .in2(_gnd_net_),
            .in3(N__15707),
            .lcout(chary_if_generate_plus_mult1_un47_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ7DB_0_9_LC_11_7_7.C_ON=1'b0;
    defparam beamY_RNIQ7DB_0_9_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ7DB_0_9_LC_11_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNIQ7DB_0_9_LC_11_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15179),
            .lcout(beamY_RNIQ7DB_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_11_8_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_11_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(N__15214),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STC_LC_11_8_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STC_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STC_LC_11_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STC_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(N__15202),
            .in2(N__15550),
            .in3(N__15196),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUC_LC_11_8_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUC_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUC_LC_11_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUC_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__15193),
            .in2(N__15551),
            .in3(N__15133),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_11_8_3.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_11_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_11_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15130),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITSR8_0_8_LC_11_8_6.C_ON=1'b0;
    defparam beamY_RNITSR8_0_8_LC_11_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNITSR8_0_8_LC_11_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNITSR8_0_8_LC_11_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15112),
            .lcout(beamY_RNITSR8_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_11_9_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_11_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(N__15716),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJG_LC_11_9_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJG_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJG_LC_11_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJG_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__15655),
            .in2(N__15598),
            .in3(N__15637),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMK_LC_11_9_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMK_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMK_LC_11_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMK_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__15575),
            .in2(N__15634),
            .in3(N__15616),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOK_LC_11_9_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOK_LC_11_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOK_LC_11_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOK_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(N__15613),
            .in2(N__15599),
            .in3(N__15439),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_9_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__15377),
            .in2(_gnd_net_),
            .in3(N__15424),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_11_9_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_11_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_11_9_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_11_9_5 (
            .in0(N__15391),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15421),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_11_9_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_11_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_11_9_6.LUT_INIT=16'b0011001100110011;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_11_9_6 (
            .in0(_gnd_net_),
            .in1(N__15390),
            .in2(_gnd_net_),
            .in3(N__15378),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
