-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 23 2015 17:44:13

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__14780\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_\ : std_logic;
signal \beamY_RNIQ8RJCCZ0Z_3_cascade_\ : std_logic;
signal \beamY_RNIQ8RJCC_0Z0Z_3\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_\ : std_logic;
signal \beamY_RNI03RTE5Z0Z_4\ : std_logic;
signal \beamY_RNI03RTE5_0Z0Z_4\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1 : std_logic;
signal \Pixel_1_RNOZ0Z_34_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un68_sum_c4 : std_logic;
signal \beamY_RNIUAN5CR1Z0Z_3\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i : std_logic;
signal \beamY_fast_RNIEGGAZ0Z_6\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0 : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_\ : std_logic;
signal \beamY_RNIGBU92Z0Z_9_cascade_\ : std_logic;
signal \beamY_RNIIDGN6_0Z0Z_7\ : std_logic;
signal \beamY_RNIIDGN6Z0Z_7_cascade_\ : std_logic;
signal \beamY_RNIPM0M5Z0Z_9_cascade_\ : std_logic;
signal \beamY_RNIPM0M5_0Z0Z_9\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_c5 : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0 : std_logic;
signal \beamY_RNI1G0FH2Z0Z_3_cascade_\ : std_logic;
signal \beamY_RNI1G0FH2_0Z0Z_3_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cascade_\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_\ : std_logic;
signal \beamY_RNICCIKUQ_0Z0Z_3\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un61_sum_c4 : std_logic;
signal \beamY_RNICCIKUQZ0Z_3\ : std_logic;
signal un4_beamylt6 : std_logic;
signal \un4_beamylt8_0_cascade_\ : std_logic;
signal un1_beamylto9_0 : std_logic;
signal \un1_beamylto9_3_cascade_\ : std_logic;
signal \un5_beamx_4_cascade_\ : std_logic;
signal \un117_pixel_6_ns_1_3_cascade_\ : std_logic;
signal \N_192_0\ : std_logic;
signal \N_192_0_cascade_\ : std_logic;
signal \N_215_0\ : std_logic;
signal \Pixel_1_RNOZ0Z_66_cascade_\ : std_logic;
signal un117_pixel_3_1_3 : std_logic;
signal \N_234_0\ : std_logic;
signal \m3_0_cascade_\ : std_logic;
signal \un115_pixel_2_0_5__N_9_cascade_\ : std_logic;
signal \g0_3_1_cascade_\ : std_logic;
signal \un115_pixel_0_a2_0_cascade_\ : std_logic;
signal \N_281\ : std_logic;
signal \N_231\ : std_logic;
signal \Pixel_1_RNOZ0Z_62\ : std_logic;
signal \N_275_0\ : std_logic;
signal \un115_pixel_13_15__m3_a0Z0Z_0\ : std_logic;
signal \un115_pixel_13_15__m3_a0Z0Z_0_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_88\ : std_logic;
signal \Pixel_1_RNOZ0Z_63\ : std_logic;
signal \un115_pixel_2_0_5__N_14\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un82_sum_cry_1 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal \G_370\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal \un4_pixel_N_3_cascade_\ : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un75_sum_iZ0\ : std_logic;
signal \N_208_0_0_1\ : std_logic;
signal \N_1260_0_0_1_cascade_\ : std_logic;
signal \Z_decfrac2_1_0_0_0_cascade_\ : std_logic;
signal \un115_pixel_3_0_3__N_8_0_0_0_cascade_\ : std_logic;
signal un117_pixel_3_1_0_1_4 : std_logic;
signal \m4_cascade_\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1 : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_\ : std_logic;
signal \beamY_fastZ0Z_4\ : std_logic;
signal \beamY_fastZ0Z_9\ : std_logic;
signal \beamY_fast_RNICEGAZ0Z_4\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2 : std_logic;
signal \beamY_RNI9I1Q6Z0Z_9_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3 : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_\ : std_logic;
signal \beamY_RNIQQREO1Z0Z_3\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un47_sum_c5 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0 : std_logic;
signal \beamY_4_rep1_RNI9H1FZ0Z1\ : std_logic;
signal \beamY_RNIHS041Z0Z_6\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0 : std_logic;
signal \beamY_RNIF8TM3Z0Z_9\ : std_logic;
signal \beamY_RNIVD444Z0Z_9_cascade_\ : std_logic;
signal \beamY_RNIGBU92Z0Z_9\ : std_logic;
signal \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1 : std_logic;
signal \N_7_0_0_0_cascade_\ : std_logic;
signal \un8_beamy_3_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_43\ : std_logic;
signal \Pixel_1_RNOZ0Z_42\ : std_logic;
signal \N_282\ : std_logic;
signal \font_un127_pixel_1_1_cascade_\ : std_logic;
signal \N_336_0\ : std_logic;
signal un5_beamx_6 : std_logic;
signal un8_beamy_3 : std_logic;
signal g1_1 : std_logic;
signal \N_283_cascade_\ : std_logic;
signal \N_285\ : std_logic;
signal font_un13_pixel_23 : std_logic;
signal font_un73_pixellt7_0 : std_logic;
signal \font_un13_pixel_23_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_60\ : std_logic;
signal \Pixel_1_RNOZ0Z_39_cascade_\ : std_logic;
signal \d_N_6_0\ : std_logic;
signal \N_6\ : std_logic;
signal \N_5_i_0\ : std_logic;
signal \g1_0_0_cascade_\ : std_logic;
signal \N_250_0_cascade_\ : std_logic;
signal \N_266_0\ : std_logic;
signal \N_242_0_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_61\ : std_logic;
signal m3_0 : std_logic;
signal \Pixel_1_RNOZ0Z_69_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_70\ : std_logic;
signal \g0_35_1_cascade_\ : std_logic;
signal \un115_pixel_13_15___m1_e_0Z0Z_1\ : std_logic;
signal \un115_pixel_13_15__i2_mux\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_2_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \un7_pixel_1_axb1_cascade_\ : std_logic;
signal \N_203_0_cascade_\ : std_logic;
signal \N_268_0\ : std_logic;
signal g0_40_1 : std_logic;
signal \N_206\ : std_logic;
signal \g0_6_1_1_cascade_\ : std_logic;
signal \g0_6_1_cascade_\ : std_logic;
signal \N_192_0_0\ : std_logic;
signal \g1_3_1_cascade_\ : std_logic;
signal g1_3 : std_logic;
signal \g0_10_1_cascade_\ : std_logic;
signal \N_309_0_cascade_\ : std_logic;
signal \N_316_0\ : std_logic;
signal \N_323_0_cascade_\ : std_logic;
signal \N_302_0_0_0\ : std_logic;
signal \N_5_0_0_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal \un21_beamy_cry_7_c_RNIM7EZ0Z3\ : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \un21_beamy_cry_8_c_RNIOAFZ0Z3\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal un11_visibleylto9_1 : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0 : std_logic;
signal \beamY_fastZ0Z_7\ : std_logic;
signal \beamY_fastZ0Z_6\ : std_logic;
signal \beamY_fastZ0Z_5\ : std_logic;
signal un11_visibleylto9_4 : std_logic;
signal \beamY_fast_RNI198KZ0Z_2_cascade_\ : std_logic;
signal font_un127_pixel_m_1 : std_logic;
signal \un21_beamy_cry_1_c_RNIALZ0Z73\ : std_logic;
signal \beamY_fastZ0Z_8\ : std_logic;
signal \beamY_fast_RNIG57DZ0Z_8\ : std_logic;
signal \beamY_fast_RNIG57DZ0Z_8_cascade_\ : std_logic;
signal un5_visibley_c6_0_1 : std_logic;
signal \un21_beamy_cry_6_c_RNIK4DZ0Z3\ : std_logic;
signal \un21_beamy_cry_2_c_RNICOZ0Z83\ : std_logic;
signal \un21_beamy_cry_5_c_RNII1CZ0Z3\ : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \beamY_RNI9DLCZ0Z_0\ : std_logic;
signal \un21_beamy_cry_3_c_RNIERZ0Z93\ : std_logic;
signal \un21_beamy_cry_4_c_RNIGUAZ0Z3\ : std_logic;
signal \N_338_0_0_0\ : std_logic;
signal \font_un127_pixel_m_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal font_un127_pixel_m_4 : std_logic;
signal \g0_0_1_cascade_\ : std_logic;
signal font_un69_pixellto3 : std_logic;
signal g0_0_2 : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_82\ : std_logic;
signal \font_un127_pixel_m_4_1_1_cascade_\ : std_logic;
signal font_un127_pixel_m_4_1 : std_logic;
signal \un7_pixel_1_c4_cascade_\ : std_logic;
signal font_un127_pixel_m_7_1_0 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\ : std_logic;
signal \N_307_0_0_1\ : std_logic;
signal \font_un13_pixel_0_1_0_0_22_cascade_\ : std_logic;
signal \beamY_RNIVV787O2Z0Z_2\ : std_logic;
signal \Pixel_1_RNOZ0Z_47\ : std_logic;
signal \N_1482_0_cascade_\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un7_pixel_1_axb2_cascade_\ : std_logic;
signal un7_pixel_1_axb2_i : std_logic;
signal \Pixel_1_RNOZ0Z_44\ : std_logic;
signal \N_305_0_cascade_\ : std_logic;
signal \N_326_0_0\ : std_logic;
signal g0_18_1 : std_logic;
signal \N_321_0_cascade_\ : std_logic;
signal \N_314_0_0_0\ : std_logic;
signal \N_328_0_0_0\ : std_logic;
signal \g1_2_0_0_cascade_\ : std_logic;
signal \N_192_0_1\ : std_logic;
signal \un117_pixel_6_1_0_1_4_cascade_\ : std_logic;
signal \N_219_0_0_1\ : std_logic;
signal un7_pixel_1_axb3_i : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal un7_pixel_1_axb3 : std_logic;
signal \un7_pixel_1_axb3_cascade_\ : std_logic;
signal un7_pixel_1_axb1 : std_logic;
signal \N_532_i\ : std_logic;
signal un117_pixel_2_6_i3_mux : std_logic;
signal un7_pixel_1_axb2 : std_logic;
signal \un4_pixel_N_3\ : std_logic;
signal \Pixel_1_RNOZ0Z_73_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_72\ : std_logic;
signal font_un36_pixel_23 : std_logic;
signal \Pixel_1_RNOZ0Z_48_cascade_\ : std_logic;
signal \N_234_0_0\ : std_logic;
signal \d_N_3_0_0\ : std_logic;
signal un7_pixel_0_axb3_i : std_logic;
signal \bfn_7_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \Pixel_1_RNOZ0Z_18\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0\ : std_logic;
signal un43lto1 : std_logic;
signal \un43lto4_1_cascade_\ : std_logic;
signal \un43lt10_cascade_\ : std_logic;
signal \un1_beamY_26\ : std_logic;
signal un42lt10 : std_logic;
signal un5_visibley_c7 : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_19\ : std_logic;
signal un1_visiblex_27 : std_logic;
signal un5_visibley_ac0_7 : std_logic;
signal \un5_visibley_ac0_7_cascade_\ : std_logic;
signal font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0 : std_logic;
signal \beamY_4_rep1_RNICDQEZ0_cascade_\ : std_logic;
signal \beamY_fastZ0Z_3\ : std_logic;
signal un5_visibley_c2 : std_logic;
signal un11_visibley : std_logic;
signal un44 : std_logic;
signal \Pixel_1_e_1\ : std_logic;
signal \beamY_fastZ0Z_2\ : std_logic;
signal \beamY_4_repZ0Z1\ : std_logic;
signal \beamY_fast_RNIK8HHZ0Z_2\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \beamY_RNIKOP3Z0Z_7\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal un8_beamylto9_1 : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1\ : std_logic;
signal un14_visibleylt9_0 : std_logic;
signal un14_visibleylt4_0 : std_logic;
signal \un3_beamx_5_cascade_\ : std_logic;
signal \N_324_0_0_0\ : std_logic;
signal \N_303_0_0_0\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal g1_0_0_0_1 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\ : std_logic;
signal \g3_0_0_0_cascade_\ : std_logic;
signal g1_4_0_0_0 : std_logic;
signal \N_1869_0_0\ : std_logic;
signal \N_1870_0_0\ : std_logic;
signal \font_un127_pixel_6_ns_1_0_0_cascade_\ : std_logic;
signal font_un13_pixel_0_1_0_0_22 : std_logic;
signal \N_520\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal \beamY_RNIJ0DBZ0Z_8\ : std_logic;
signal \VSync_c\ : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4 : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum0_2 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4 : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum1_4 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum0_4 : std_logic;
signal \un7_pixel_0_axb4_cascade_\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum1_5 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum0_5 : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal un7_pixel_0_axb4 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal un4_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal un7_pixel_0_axb4_i : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal un4_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal un7_pixel_0_axb3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum1_3 : std_logic;
signal un4_pixel_if_generate_plus_mult1_un47_sum0_3 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_3 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \beamY_RNIALEQZ0Z_9\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\ : std_logic;
signal \beamY_RNIALEQ_1Z0Z_9\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum\ : std_logic;
signal \beamY_RNIQNF11_0Z0Z_8\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16\ : std_logic;
signal \HSync_c\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx : std_logic;
signal un5_visiblex_i_25 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i : std_logic;
signal if_generate_plus_mult1_un47_sum_m_1 : std_logic;
signal un5_visiblex_i_0_25 : std_logic;
signal \N_32\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx : std_logic;
signal if_generate_plus_mult1_un47_sum_0_cry_3_ma : std_logic;
signal \N_158_0_i\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7 : std_logic;
signal \N_20_i\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal un18_beamylt4 : std_logic;
signal \un18_beamylto9_2_cascade_\ : std_logic;
signal un4_beamy_0 : std_logic;
signal \un18_beamylt10_0_cascade_\ : std_logic;
signal un8_beamy : std_logic;
signal un13_beamylt7 : std_logic;
signal \un15_beamy_2_cascade_\ : std_logic;
signal un15_beamy : std_logic;
signal \un1_beamx_2_cascade_\ : std_logic;
signal un1_beamx : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un3_beamx_7 : std_logic;
signal un1_beamx_2 : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0\ : std_logic;
signal un3_beamx_g : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un33_sum_i : std_logic;
signal \PixelClock_g\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un75_sum : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un1_visiblex_24 : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\ : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\ : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum : std_logic;
signal font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \PixelDebug_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    PixelDebug <= \PixelDebug_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__6190\,
            RESETB => \N__14610\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14780\,
            DIN => \N__14779\,
            DOUT => \N__14778\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14780\,
            PADOUT => \N__14779\,
            PADIN => \N__14778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11317\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14771\,
            DIN => \N__14770\,
            DOUT => \N__14769\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14771\,
            PADOUT => \N__14770\,
            PADIN => \N__14769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12366\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14762\,
            DIN => \N__14761\,
            DOUT => \N__14760\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14762\,
            PADOUT => \N__14761\,
            PADIN => \N__14760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14753\,
            DIN => \N__14752\,
            DOUT => \N__14751\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14753\,
            PADOUT => \N__14752\,
            PADIN => \N__14751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14744\,
            DIN => \N__14743\,
            DOUT => \N__14742\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14744\,
            PADOUT => \N__14743\,
            PADIN => \N__14742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14735\,
            DIN => \N__14734\,
            DOUT => \N__14733\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14735\,
            PADOUT => \N__14734\,
            PADIN => \N__14733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12373\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14726\,
            DIN => \N__14725\,
            DOUT => \N__14724\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14726\,
            PADOUT => \N__14725\,
            PADIN => \N__14724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8116\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__14707\,
            I => \N__14704\
        );

    \I__3379\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14701\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14691\
        );

    \I__3377\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14688\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14685\
        );

    \I__3375\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14682\
        );

    \I__3374\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14679\
        );

    \I__3373\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14676\
        );

    \I__3372\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14671\
        );

    \I__3371\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14671\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__14691\,
            I => \N__14666\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__14688\,
            I => \N__14666\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__14685\,
            I => \N__14663\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__14682\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__14679\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14676\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__14671\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__14666\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__14663\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__3360\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14644\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__14644\,
            I => \N__14641\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__14638\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0\
        );

    \I__3356\ : InMux
    port map (
            O => \N__14635\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__3355\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14627\
        );

    \I__3354\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14624\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__14630\,
            I => \N__14620\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14614\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__14624\,
            I => \N__14614\
        );

    \I__3350\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14611\
        );

    \I__3349\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14601\
        );

    \I__3348\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14601\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__14614\,
            I => \N__14596\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14596\
        );

    \I__3345\ : IoInMux
    port map (
            O => \N__14610\,
            I => \N__14589\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__14609\,
            I => \N__14586\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__14608\,
            I => \N__14583\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__14607\,
            I => \N__14580\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__14606\,
            I => \N__14577\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__14601\,
            I => \N__14572\
        );

    \I__3339\ : Span4Mux_s3_h
    port map (
            O => \N__14596\,
            I => \N__14572\
        );

    \I__3338\ : InMux
    port map (
            O => \N__14595\,
            I => \N__14569\
        );

    \I__3337\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14566\
        );

    \I__3336\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14563\
        );

    \I__3335\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14560\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__14589\,
            I => \N__14557\
        );

    \I__3333\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14553\
        );

    \I__3332\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14550\
        );

    \I__3331\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14545\
        );

    \I__3330\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14545\
        );

    \I__3329\ : Sp12to4
    port map (
            O => \N__14572\,
            I => \N__14536\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14536\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__14566\,
            I => \N__14536\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__14563\,
            I => \N__14536\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__14560\,
            I => \N__14533\
        );

    \I__3324\ : IoSpan4Mux
    port map (
            O => \N__14557\,
            I => \N__14530\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__14556\,
            I => \N__14527\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14520\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__14550\,
            I => \N__14520\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__14545\,
            I => \N__14520\
        );

    \I__3319\ : Span12Mux_v
    port map (
            O => \N__14536\,
            I => \N__14517\
        );

    \I__3318\ : Span4Mux_v
    port map (
            O => \N__14533\,
            I => \N__14514\
        );

    \I__3317\ : IoSpan4Mux
    port map (
            O => \N__14530\,
            I => \N__14511\
        );

    \I__3316\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14508\
        );

    \I__3315\ : Span4Mux_v
    port map (
            O => \N__14520\,
            I => \N__14505\
        );

    \I__3314\ : Odrv12
    port map (
            O => \N__14517\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__14514\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__14511\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__14508\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__14505\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3309\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14490\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14487\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__14490\,
            I => \N__14484\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__14487\,
            I => \N__14481\
        );

    \I__3305\ : Span4Mux_v
    port map (
            O => \N__14484\,
            I => \N__14478\
        );

    \I__3304\ : Span4Mux_v
    port map (
            O => \N__14481\,
            I => \N__14475\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__14478\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__14475\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0\
        );

    \I__3301\ : InMux
    port map (
            O => \N__14470\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__3300\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14464\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__14464\,
            I => \N__14461\
        );

    \I__3298\ : Span4Mux_v
    port map (
            O => \N__14461\,
            I => \N__14458\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__14458\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\
        );

    \I__3296\ : InMux
    port map (
            O => \N__14455\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__3295\ : InMux
    port map (
            O => \N__14452\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__3294\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14445\
        );

    \I__3293\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14442\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__14445\,
            I => \N__14437\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14437\
        );

    \I__3290\ : Span4Mux_h
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__14434\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__14431\,
            I => \N__14428\
        );

    \I__3287\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14425\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__14425\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\
        );

    \I__3285\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14418\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__14421\,
            I => \N__14415\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__14418\,
            I => \N__14403\
        );

    \I__3282\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14400\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__14414\,
            I => \N__14397\
        );

    \I__3280\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14394\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14391\
        );

    \I__3278\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14384\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14384\
        );

    \I__3276\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14384\
        );

    \I__3275\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14377\
        );

    \I__3274\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14377\
        );

    \I__3273\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14377\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__14403\,
            I => \N__14371\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14367\
        );

    \I__3270\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14364\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14352\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__14391\,
            I => \N__14347\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14347\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14344\
        );

    \I__3265\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14337\
        );

    \I__3264\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14337\
        );

    \I__3263\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14337\
        );

    \I__3262\ : Span4Mux_v
    port map (
            O => \N__14371\,
            I => \N__14334\
        );

    \I__3261\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14331\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__14367\,
            I => \N__14326\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__14364\,
            I => \N__14326\
        );

    \I__3258\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14321\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14321\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14316\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14316\
        );

    \I__3254\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14305\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14305\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14305\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14305\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14355\,
            I => \N__14305\
        );

    \I__3249\ : Span4Mux_v
    port map (
            O => \N__14352\,
            I => \N__14296\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__14347\,
            I => \N__14296\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__14344\,
            I => \N__14296\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__14337\,
            I => \N__14296\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__14334\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14331\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__14326\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__14321\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__14316\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14305\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__14296\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__14281\,
            I => \N__14278\
        );

    \I__3237\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__14275\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__14272\,
            I => \N__14269\
        );

    \I__3234\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__14266\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_i
        );

    \I__3232\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__3231\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14257\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__14257\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__14254\,
            I => \N__14251\
        );

    \I__3228\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14245\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__14245\,
            I => \N__14242\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__14242\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11\
        );

    \I__3224\ : InMux
    port map (
            O => \N__14239\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__14236\,
            I => \N__14233\
        );

    \I__3222\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__14230\,
            I => \N__14227\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__14227\,
            I => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__14224\,
            I => \N__14221\
        );

    \I__3218\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14218\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__14218\,
            I => \N__14215\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__14215\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1\
        );

    \I__3215\ : InMux
    port map (
            O => \N__14212\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__14209\,
            I => \N__14206\
        );

    \I__3213\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14203\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__14203\,
            I => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0\
        );

    \I__3211\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14197\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__14197\,
            I => \N__14194\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__14194\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__3208\ : InMux
    port map (
            O => \N__14191\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__3207\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14185\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14185\,
            I => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__3205\ : InMux
    port map (
            O => \N__14182\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__3204\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14176\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14171\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14168\
        );

    \I__3201\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14165\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__14171\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__14168\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14165\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__14152\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_i
        );

    \I__3194\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14140\
        );

    \I__3193\ : InMux
    port map (
            O => \N__14148\,
            I => \N__14140\
        );

    \I__3192\ : InMux
    port map (
            O => \N__14147\,
            I => \N__14140\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__14140\,
            I => \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0\
        );

    \I__3190\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14131\
        );

    \I__3189\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14131\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__14131\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_i_8
        );

    \I__3187\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14124\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__14127\,
            I => \N__14120\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__14124\,
            I => \N__14116\
        );

    \I__3184\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14113\
        );

    \I__3183\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14110\
        );

    \I__3182\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14107\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__14116\,
            I => \N__14102\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__14113\,
            I => \N__14102\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__14110\,
            I => \N__14099\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__14107\,
            I => \beamXZ0Z_2\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__14102\,
            I => \beamXZ0Z_2\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__14099\,
            I => \beamXZ0Z_2\
        );

    \I__3175\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14087\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14080\
        );

    \I__3173\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14080\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__14087\,
            I => \N__14077\
        );

    \I__3171\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14074\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14071\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__14080\,
            I => \N__14068\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__14077\,
            I => \N__14065\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14074\,
            I => \N__14062\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__14071\,
            I => \N__14059\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__14068\,
            I => \N__14056\
        );

    \I__3164\ : Span4Mux_h
    port map (
            O => \N__14065\,
            I => \N__14053\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__14062\,
            I => \N__14048\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__14059\,
            I => \N__14048\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__14056\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__14053\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__14048\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__3158\ : InMux
    port map (
            O => \N__14041\,
            I => un5_visiblex_cry_1
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__14038\,
            I => \N__14033\
        );

    \I__3156\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14029\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__14036\,
            I => \N__14026\
        );

    \I__3154\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14022\
        );

    \I__3153\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14019\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__14029\,
            I => \N__14016\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14026\,
            I => \N__14013\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14010\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__14022\,
            I => \N__14007\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__14019\,
            I => \N__14002\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__14016\,
            I => \N__14002\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__14013\,
            I => \N__13999\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__14010\,
            I => \beamXZ0Z_3\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__14007\,
            I => \beamXZ0Z_3\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__14002\,
            I => \beamXZ0Z_3\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__13999\,
            I => \beamXZ0Z_3\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__13990\,
            I => \N__13987\
        );

    \I__3140\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13984\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__13984\,
            I => \N__13979\
        );

    \I__3138\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13976\
        );

    \I__3137\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13972\
        );

    \I__3136\ : Span4Mux_v
    port map (
            O => \N__13979\,
            I => \N__13965\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__13976\,
            I => \N__13965\
        );

    \I__3134\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13962\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__13972\,
            I => \N__13959\
        );

    \I__3132\ : InMux
    port map (
            O => \N__13971\,
            I => \N__13956\
        );

    \I__3131\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13953\
        );

    \I__3130\ : Span4Mux_v
    port map (
            O => \N__13965\,
            I => \N__13950\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__13962\,
            I => \N__13947\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__13959\,
            I => \N__13944\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13939\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__13953\,
            I => \N__13939\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__13950\,
            I => un1_visiblex_24
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__13947\,
            I => un1_visiblex_24
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__13944\,
            I => un1_visiblex_24
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__13939\,
            I => un1_visiblex_24
        );

    \I__3121\ : InMux
    port map (
            O => \N__13930\,
            I => un5_visiblex_cry_2
        );

    \I__3120\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13920\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__13926\,
            I => \N__13917\
        );

    \I__3118\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13913\
        );

    \I__3117\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13908\
        );

    \I__3116\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13908\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__13920\,
            I => \N__13905\
        );

    \I__3114\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13902\
        );

    \I__3113\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13899\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__13913\,
            I => \N__13892\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__13908\,
            I => \N__13892\
        );

    \I__3110\ : Span4Mux_h
    port map (
            O => \N__13905\,
            I => \N__13892\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__13902\,
            I => \N__13889\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__13899\,
            I => \beamXZ0Z_4\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__13892\,
            I => \beamXZ0Z_4\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__13889\,
            I => \beamXZ0Z_4\
        );

    \I__3105\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13876\
        );

    \I__3104\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13871\
        );

    \I__3103\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13871\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__13879\,
            I => \N__13865\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__13876\,
            I => \N__13860\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__13871\,
            I => \N__13860\
        );

    \I__3099\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13857\
        );

    \I__3098\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13853\
        );

    \I__3097\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13850\
        );

    \I__3096\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13847\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__13860\,
            I => \N__13842\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__13857\,
            I => \N__13842\
        );

    \I__3093\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13839\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__13853\,
            I => \N__13836\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__13850\,
            I => \N__13833\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13830\
        );

    \I__3089\ : Span4Mux_v
    port map (
            O => \N__13842\,
            I => \N__13825\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__13839\,
            I => \N__13825\
        );

    \I__3087\ : Span4Mux_h
    port map (
            O => \N__13836\,
            I => \N__13820\
        );

    \I__3086\ : Span4Mux_h
    port map (
            O => \N__13833\,
            I => \N__13820\
        );

    \I__3085\ : Odrv4
    port map (
            O => \N__13830\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__13825\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__13820\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__3082\ : InMux
    port map (
            O => \N__13813\,
            I => un5_visiblex_cry_3
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \N__13805\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__13809\,
            I => \N__13801\
        );

    \I__3079\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13796\
        );

    \I__3078\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13791\
        );

    \I__3077\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13791\
        );

    \I__3076\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13788\
        );

    \I__3075\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13785\
        );

    \I__3074\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13782\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__13796\,
            I => \N__13777\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__13791\,
            I => \N__13777\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13788\,
            I => \N__13774\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__13785\,
            I => \beamXZ0Z_5\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__13782\,
            I => \beamXZ0Z_5\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__13777\,
            I => \beamXZ0Z_5\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__13774\,
            I => \beamXZ0Z_5\
        );

    \I__3066\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13756\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13753\
        );

    \I__3064\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13750\
        );

    \I__3063\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13747\
        );

    \I__3062\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13744\
        );

    \I__3061\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13741\
        );

    \I__3060\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13738\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13735\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13732\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13750\,
            I => \N__13729\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__13747\,
            I => \N__13726\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13723\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13720\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__13738\,
            I => \N__13717\
        );

    \I__3052\ : Span4Mux_h
    port map (
            O => \N__13735\,
            I => \N__13710\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__13732\,
            I => \N__13710\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__13729\,
            I => \N__13710\
        );

    \I__3049\ : Span4Mux_h
    port map (
            O => \N__13726\,
            I => \N__13703\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__13723\,
            I => \N__13703\
        );

    \I__3047\ : Span4Mux_h
    port map (
            O => \N__13720\,
            I => \N__13703\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__13717\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__13710\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__13703\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__3043\ : InMux
    port map (
            O => \N__13696\,
            I => un5_visiblex_cry_4
        );

    \I__3042\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__13690\,
            I => \N__13683\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__13689\,
            I => \N__13680\
        );

    \I__3039\ : InMux
    port map (
            O => \N__13688\,
            I => \N__13674\
        );

    \I__3038\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13674\
        );

    \I__3037\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13671\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__13683\,
            I => \N__13668\
        );

    \I__3035\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13665\
        );

    \I__3034\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13662\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__13674\,
            I => \N__13657\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__13671\,
            I => \N__13657\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__13668\,
            I => \N__13654\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__13665\,
            I => \N__13651\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__13662\,
            I => \beamXZ0Z_6\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__13657\,
            I => \beamXZ0Z_6\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__13654\,
            I => \beamXZ0Z_6\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__13651\,
            I => \beamXZ0Z_6\
        );

    \I__3025\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13638\
        );

    \I__3024\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13629\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__13638\,
            I => \N__13626\
        );

    \I__3022\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13623\
        );

    \I__3021\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13620\
        );

    \I__3020\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13617\
        );

    \I__3019\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13614\
        );

    \I__3018\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13611\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__13632\,
            I => \N__13608\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13629\,
            I => \N__13604\
        );

    \I__3015\ : Span4Mux_h
    port map (
            O => \N__13626\,
            I => \N__13597\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13597\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__13620\,
            I => \N__13597\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__13617\,
            I => \N__13594\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__13614\,
            I => \N__13591\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__13611\,
            I => \N__13588\
        );

    \I__3009\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13585\
        );

    \I__3008\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13582\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__13604\,
            I => \N__13579\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__13597\,
            I => \N__13572\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__13594\,
            I => \N__13572\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__13591\,
            I => \N__13572\
        );

    \I__3003\ : Odrv12
    port map (
            O => \N__13588\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__13585\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__13582\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__13579\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__13572\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2998\ : InMux
    port map (
            O => \N__13561\,
            I => un5_visiblex_cry_5
        );

    \I__2997\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13547\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13547\
        );

    \I__2995\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13547\
        );

    \I__2994\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13543\
        );

    \I__2993\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13540\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13537\
        );

    \I__2991\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13534\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__13543\,
            I => \N__13531\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__13540\,
            I => \beamXZ0Z_7\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__13537\,
            I => \beamXZ0Z_7\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__13534\,
            I => \beamXZ0Z_7\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__13531\,
            I => \beamXZ0Z_7\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__13522\,
            I => \N__13518\
        );

    \I__2984\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13515\
        );

    \I__2983\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13512\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13507\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__13512\,
            I => \N__13504\
        );

    \I__2980\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13496\
        );

    \I__2979\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13493\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__13507\,
            I => \N__13490\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__13504\,
            I => \N__13487\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13482\
        );

    \I__2975\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13482\
        );

    \I__2974\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13479\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13474\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13474\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__13496\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__13493\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__13490\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__13487\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__13482\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__13479\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__13474\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__2964\ : InMux
    port map (
            O => \N__13459\,
            I => un5_visiblex_cry_6
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__13456\,
            I => \N__13451\
        );

    \I__2962\ : InMux
    port map (
            O => \N__13455\,
            I => \N__13445\
        );

    \I__2961\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13445\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13442\
        );

    \I__2959\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13439\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13436\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__13442\,
            I => \N__13433\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__13439\,
            I => \beamXZ0Z_8\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__13436\,
            I => \beamXZ0Z_8\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__13433\,
            I => \beamXZ0Z_8\
        );

    \I__2953\ : InMux
    port map (
            O => \N__13426\,
            I => \bfn_9_12_0_\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__13423\,
            I => \N__13419\
        );

    \I__2951\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13412\
        );

    \I__2950\ : InMux
    port map (
            O => \N__13419\,
            I => \N__13412\
        );

    \I__2949\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13409\
        );

    \I__2948\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13406\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__13412\,
            I => \N__13403\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__13409\,
            I => \N__13400\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__13406\,
            I => \beamXZ0Z_9\
        );

    \I__2944\ : Odrv12
    port map (
            O => \N__13403\,
            I => \beamXZ0Z_9\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__13400\,
            I => \beamXZ0Z_9\
        );

    \I__2942\ : InMux
    port map (
            O => \N__13393\,
            I => un5_visiblex_cry_8
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__13390\,
            I => \N__13385\
        );

    \I__2940\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13379\
        );

    \I__2939\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13379\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13376\
        );

    \I__2937\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13373\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__13379\,
            I => \N__13370\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__13376\,
            I => \N__13367\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__13373\,
            I => \beamXZ0Z_10\
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__13370\,
            I => \beamXZ0Z_10\
        );

    \I__2932\ : Odrv12
    port map (
            O => \N__13367\,
            I => \beamXZ0Z_10\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13357\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__13357\,
            I => \N__13354\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__13354\,
            I => un3_beamx_7
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__13351\,
            I => \N__13348\
        );

    \I__2927\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13344\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13341\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__13344\,
            I => \N__13338\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13341\,
            I => un1_beamx_2
        );

    \I__2923\ : Odrv12
    port map (
            O => \N__13338\,
            I => un1_beamx_2
        );

    \I__2922\ : IoInMux
    port map (
            O => \N__13333\,
            I => \N__13330\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13327\
        );

    \I__2920\ : Span4Mux_s0_h
    port map (
            O => \N__13327\,
            I => \N__13324\
        );

    \I__2919\ : Span4Mux_h
    port map (
            O => \N__13324\,
            I => \N__13321\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__13321\,
            I => \N__13318\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__13318\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__2916\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13309\
        );

    \I__2915\ : InMux
    port map (
            O => \N__13314\,
            I => \N__13309\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__13309\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__13306\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__2911\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13297\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__13297\,
            I => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13287\
        );

    \I__2908\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13284\
        );

    \I__2907\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13281\
        );

    \I__2906\ : InMux
    port map (
            O => \N__13291\,
            I => \N__13276\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13276\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13287\,
            I => \N__13267\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__13284\,
            I => \N__13264\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__13281\,
            I => \N__13261\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__13276\,
            I => \N__13258\
        );

    \I__2900\ : CEMux
    port map (
            O => \N__13275\,
            I => \N__13237\
        );

    \I__2899\ : CEMux
    port map (
            O => \N__13274\,
            I => \N__13237\
        );

    \I__2898\ : CEMux
    port map (
            O => \N__13273\,
            I => \N__13237\
        );

    \I__2897\ : CEMux
    port map (
            O => \N__13272\,
            I => \N__13237\
        );

    \I__2896\ : CEMux
    port map (
            O => \N__13271\,
            I => \N__13237\
        );

    \I__2895\ : CEMux
    port map (
            O => \N__13270\,
            I => \N__13237\
        );

    \I__2894\ : Glb2LocalMux
    port map (
            O => \N__13267\,
            I => \N__13237\
        );

    \I__2893\ : Glb2LocalMux
    port map (
            O => \N__13264\,
            I => \N__13237\
        );

    \I__2892\ : Glb2LocalMux
    port map (
            O => \N__13261\,
            I => \N__13237\
        );

    \I__2891\ : Glb2LocalMux
    port map (
            O => \N__13258\,
            I => \N__13237\
        );

    \I__2890\ : GlobalMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__2889\ : gio2CtrlBuf
    port map (
            O => \N__13234\,
            I => un3_beamx_g
        );

    \I__2888\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__13228\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_i
        );

    \I__2886\ : ClkMux
    port map (
            O => \N__13225\,
            I => \N__13186\
        );

    \I__2885\ : ClkMux
    port map (
            O => \N__13224\,
            I => \N__13186\
        );

    \I__2884\ : ClkMux
    port map (
            O => \N__13223\,
            I => \N__13186\
        );

    \I__2883\ : ClkMux
    port map (
            O => \N__13222\,
            I => \N__13186\
        );

    \I__2882\ : ClkMux
    port map (
            O => \N__13221\,
            I => \N__13186\
        );

    \I__2881\ : ClkMux
    port map (
            O => \N__13220\,
            I => \N__13186\
        );

    \I__2880\ : ClkMux
    port map (
            O => \N__13219\,
            I => \N__13186\
        );

    \I__2879\ : ClkMux
    port map (
            O => \N__13218\,
            I => \N__13186\
        );

    \I__2878\ : ClkMux
    port map (
            O => \N__13217\,
            I => \N__13186\
        );

    \I__2877\ : ClkMux
    port map (
            O => \N__13216\,
            I => \N__13186\
        );

    \I__2876\ : ClkMux
    port map (
            O => \N__13215\,
            I => \N__13186\
        );

    \I__2875\ : ClkMux
    port map (
            O => \N__13214\,
            I => \N__13186\
        );

    \I__2874\ : ClkMux
    port map (
            O => \N__13213\,
            I => \N__13186\
        );

    \I__2873\ : GlobalMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__2872\ : gio2CtrlBuf
    port map (
            O => \N__13183\,
            I => \PixelClock_g\
        );

    \I__2871\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13175\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13172\
        );

    \I__2869\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13169\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13161\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__13172\,
            I => \N__13156\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__13169\,
            I => \N__13156\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13153\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__13167\,
            I => \N__13150\
        );

    \I__2863\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13145\
        );

    \I__2862\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13145\
        );

    \I__2861\ : InMux
    port map (
            O => \N__13164\,
            I => \N__13142\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__13161\,
            I => \N__13139\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__13156\,
            I => \N__13134\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__13153\,
            I => \N__13134\
        );

    \I__2857\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13131\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__13145\,
            I => \beamXZ0Z_0\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__13142\,
            I => \beamXZ0Z_0\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__13139\,
            I => \beamXZ0Z_0\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__13134\,
            I => \beamXZ0Z_0\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__13131\,
            I => \beamXZ0Z_0\
        );

    \I__2851\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13115\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \N__13110\
        );

    \I__2849\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13107\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__13115\,
            I => \N__13104\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \N__13101\
        );

    \I__2846\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13098\
        );

    \I__2845\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13095\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__13107\,
            I => \N__13092\
        );

    \I__2843\ : Span4Mux_h
    port map (
            O => \N__13104\,
            I => \N__13089\
        );

    \I__2842\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13086\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__13098\,
            I => \beamXZ0Z_1\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__13095\,
            I => \beamXZ0Z_1\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__13092\,
            I => \beamXZ0Z_1\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__13089\,
            I => \beamXZ0Z_1\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__13086\,
            I => \beamXZ0Z_1\
        );

    \I__2836\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13061\
        );

    \I__2835\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13061\
        );

    \I__2834\ : InMux
    port map (
            O => \N__13073\,
            I => \N__13058\
        );

    \I__2833\ : InMux
    port map (
            O => \N__13072\,
            I => \N__13052\
        );

    \I__2832\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13052\
        );

    \I__2831\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13049\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13040\
        );

    \I__2829\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13040\
        );

    \I__2828\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13040\
        );

    \I__2827\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13040\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13037\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__13058\,
            I => \N__13034\
        );

    \I__2824\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13031\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13024\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13024\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13040\,
            I => \N__13024\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__13037\,
            I => \N__13019\
        );

    \I__2819\ : Span4Mux_v
    port map (
            O => \N__13034\,
            I => \N__13019\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__13031\,
            I => \N__13016\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__13024\,
            I => \N__13013\
        );

    \I__2816\ : Sp12to4
    port map (
            O => \N__13019\,
            I => \N__13008\
        );

    \I__2815\ : Span12Mux_s5_v
    port map (
            O => \N__13016\,
            I => \N__13008\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__13013\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__13008\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2812\ : InMux
    port map (
            O => \N__13003\,
            I => un5_visiblex_cry_0
        );

    \I__2811\ : InMux
    port map (
            O => \N__13000\,
            I => un8_beamx_cry_1
        );

    \I__2810\ : InMux
    port map (
            O => \N__12997\,
            I => un8_beamx_cry_2
        );

    \I__2809\ : InMux
    port map (
            O => \N__12994\,
            I => un8_beamx_cry_3
        );

    \I__2808\ : InMux
    port map (
            O => \N__12991\,
            I => un8_beamx_cry_4
        );

    \I__2807\ : InMux
    port map (
            O => \N__12988\,
            I => un8_beamx_cry_5
        );

    \I__2806\ : InMux
    port map (
            O => \N__12985\,
            I => un8_beamx_cry_6
        );

    \I__2805\ : InMux
    port map (
            O => \N__12982\,
            I => un8_beamx_cry_7
        );

    \I__2804\ : InMux
    port map (
            O => \N__12979\,
            I => \bfn_9_10_0_\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12976\,
            I => un8_beamx_cry_9
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__12973\,
            I => \N__12970\
        );

    \I__2801\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12967\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__12967\,
            I => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12964\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__12961\,
            I => \N__12958\
        );

    \I__2797\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12955\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__12955\,
            I => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1\
        );

    \I__2795\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12949\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__12949\,
            I => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12946\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__2792\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12940\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__12940\,
            I => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62\
        );

    \I__2790\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12934\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__12934\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__2788\ : InMux
    port map (
            O => \N__12931\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__2787\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12925\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__12925\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__2785\ : InMux
    port map (
            O => \N__12922\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__2784\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12915\
        );

    \I__2783\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12912\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__12915\,
            I => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__12912\,
            I => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__12907\,
            I => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__12904\,
            I => \N__12900\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12892\
        );

    \I__2776\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12892\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__12892\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__2774\ : InMux
    port map (
            O => \N__12889\,
            I => \N__12884\
        );

    \I__2773\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12879\
        );

    \I__2772\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12879\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__12884\,
            I => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__12879\,
            I => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__12874\,
            I => \N__12870\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__12873\,
            I => \N__12867\
        );

    \I__2767\ : InMux
    port map (
            O => \N__12870\,
            I => \N__12862\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12862\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__12862\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__2764\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12856\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__12856\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__2762\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12850\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__12850\,
            I => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12847\,
            I => un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__12844\,
            I => \N__12841\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12841\,
            I => \N__12837\
        );

    \I__2757\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12837\,
            I => \N__12829\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__12834\,
            I => \N__12829\
        );

    \I__2754\ : Span4Mux_h
    port map (
            O => \N__12829\,
            I => \N__12826\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__12826\,
            I => un18_beamylt4
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__12823\,
            I => \un18_beamylto9_2_cascade_\
        );

    \I__2751\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12817\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__12817\,
            I => \N__12814\
        );

    \I__2749\ : Odrv12
    port map (
            O => \N__12814\,
            I => un4_beamy_0
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__12811\,
            I => \un18_beamylt10_0_cascade_\
        );

    \I__2747\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12805\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__12805\,
            I => \N__12802\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__12802\,
            I => \N__12799\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__12799\,
            I => un8_beamy
        );

    \I__2743\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12793\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12793\,
            I => un13_beamylt7
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__12790\,
            I => \un15_beamy_2_cascade_\
        );

    \I__2740\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12784\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12784\,
            I => \N__12780\
        );

    \I__2738\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12777\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__12780\,
            I => \N__12774\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__12777\,
            I => \N__12771\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__12774\,
            I => un15_beamy
        );

    \I__2734\ : Odrv12
    port map (
            O => \N__12771\,
            I => un15_beamy
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__12766\,
            I => \un1_beamx_2_cascade_\
        );

    \I__2732\ : InMux
    port map (
            O => \N__12763\,
            I => \N__12759\
        );

    \I__2731\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12756\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__12759\,
            I => \N__12751\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__12756\,
            I => \N__12751\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__12751\,
            I => un1_beamx
        );

    \I__2727\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12745\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__12745\,
            I => un1_beamxlt10_0
        );

    \I__2725\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12739\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12734\
        );

    \I__2723\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12729\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12729\
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__12734\,
            I => \N_32\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__12729\,
            I => \N_32\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12721\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__12721\,
            I => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__12718\,
            I => \N__12715\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12712\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__12712\,
            I => if_generate_plus_mult1_un47_sum_0_cry_3_ma
        );

    \I__2714\ : InMux
    port map (
            O => \N__12709\,
            I => \N__12706\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__12706\,
            I => \N_158_0_i\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12703\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__2711\ : InMux
    port map (
            O => \N__12700\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__2710\ : InMux
    port map (
            O => \N__12697\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__2709\ : InMux
    port map (
            O => \N__12694\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7
        );

    \I__2708\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12687\
        );

    \I__2707\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12683\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__12687\,
            I => \N__12680\
        );

    \I__2705\ : InMux
    port map (
            O => \N__12686\,
            I => \N__12674\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__12683\,
            I => \N__12669\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__12680\,
            I => \N__12669\
        );

    \I__2702\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12666\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__12678\,
            I => \N__12663\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12658\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12653\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__12669\,
            I => \N__12650\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__12666\,
            I => \N__12647\
        );

    \I__2696\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12642\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12642\
        );

    \I__2694\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12637\
        );

    \I__2693\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12637\
        );

    \I__2692\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12632\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12632\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__12653\,
            I => \N_20_i\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__12650\,
            I => \N_20_i\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__12647\,
            I => \N_20_i\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__12642\,
            I => \N_20_i\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12637\,
            I => \N_20_i\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N_20_i\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__12619\,
            I => \N__12616\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12613\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__12613\,
            I => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx
        );

    \I__2681\ : InMux
    port map (
            O => \N__12610\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__2680\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12603\
        );

    \I__2679\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12600\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__12600\,
            I => \N__12594\
        );

    \I__2676\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12591\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__12594\,
            I => \N__12588\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12591\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__12588\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__12583\,
            I => \N__12580\
        );

    \I__2671\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__12577\,
            I => un5_visiblex_i_24
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__12574\,
            I => \N__12571\
        );

    \I__2668\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__12568\,
            I => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx
        );

    \I__2666\ : InMux
    port map (
            O => \N__12565\,
            I => \N__12562\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__12562\,
            I => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__12559\,
            I => \N__12556\
        );

    \I__2663\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12553\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__12553\,
            I => un5_visiblex_i_25
        );

    \I__2661\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__12547\,
            I => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__2658\ : InMux
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__12538\,
            I => font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i
        );

    \I__2656\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12532\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__12532\,
            I => \N__12529\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__12529\,
            I => \N__12526\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__12526\,
            I => if_generate_plus_mult1_un47_sum_m_1
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__2651\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12517\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__12517\,
            I => un5_visiblex_i_0_25
        );

    \I__2649\ : InMux
    port map (
            O => \N__12514\,
            I => \N__12511\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__12511\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__2647\ : InMux
    port map (
            O => \N__12508\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__2646\ : InMux
    port map (
            O => \N__12505\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__2645\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12498\
        );

    \I__2644\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12495\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__12498\,
            I => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__12495\,
            I => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__12490\,
            I => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__12487\,
            I => \N__12483\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__12486\,
            I => \N__12480\
        );

    \I__2638\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12475\
        );

    \I__2637\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12475\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__12475\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__12472\,
            I => \N__12469\
        );

    \I__2634\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12466\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__12466\,
            I => \N__12463\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__12463\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__12460\,
            I => \N__12457\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12454\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__12454\,
            I => \N__12451\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__12451\,
            I => \N__12448\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__12448\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1\
        );

    \I__2626\ : InMux
    port map (
            O => \N__12445\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__12442\,
            I => \N__12439\
        );

    \I__2624\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12436\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12433\
        );

    \I__2622\ : Odrv12
    port map (
            O => \N__12433\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2\
        );

    \I__2621\ : InMux
    port map (
            O => \N__12430\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__2620\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12424\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12421\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__12421\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__2617\ : InMux
    port map (
            O => \N__12418\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__2616\ : InMux
    port map (
            O => \N__12415\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__2615\ : InMux
    port map (
            O => \N__12412\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__2614\ : InMux
    port map (
            O => \N__12409\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__2613\ : InMux
    port map (
            O => \N__12406\,
            I => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__2612\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12400\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__12400\,
            I => \N__12397\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__12397\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__12394\,
            I => \N__12391\
        );

    \I__2608\ : InMux
    port map (
            O => \N__12391\,
            I => \N__12388\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12388\,
            I => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0\
        );

    \I__2606\ : InMux
    port map (
            O => \N__12385\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__2605\ : InMux
    port map (
            O => \N__12382\,
            I => \N__12379\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12379\,
            I => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12376\,
            I => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__2602\ : IoInMux
    port map (
            O => \N__12373\,
            I => \N__12370\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12370\,
            I => \N__12367\
        );

    \I__2600\ : Span4Mux_s2_v
    port map (
            O => \N__12367\,
            I => \N__12363\
        );

    \I__2599\ : IoInMux
    port map (
            O => \N__12366\,
            I => \N__12360\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__12363\,
            I => \N__12357\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__12360\,
            I => \N__12354\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__2595\ : Span4Mux_s3_v
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__12351\,
            I => \HSync_c\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__12348\,
            I => \HSync_c\
        );

    \I__2592\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__2591\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12337\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__12337\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__12334\,
            I => \N__12331\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__12328\,
            I => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156\
        );

    \I__2586\ : InMux
    port map (
            O => \N__12325\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__2585\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12319\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__12319\,
            I => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12316\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2582\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12310\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__12310\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__2580\ : InMux
    port map (
            O => \N__12307\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2579\ : InMux
    port map (
            O => \N__12304\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2578\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12298\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12298\,
            I => font_un13_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__2576\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12290\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12287\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12284\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__12290\,
            I => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__12287\,
            I => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__12284\,
            I => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__12277\,
            I => \N__12273\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__12276\,
            I => \N__12270\
        );

    \I__2568\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12265\
        );

    \I__2567\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12265\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__12265\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__2565\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12259\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__12259\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \N__12253\
        );

    \I__2562\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__12250\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i
        );

    \I__2560\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12244\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12244\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__2558\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12238\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__12238\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983\
        );

    \I__2556\ : InMux
    port map (
            O => \N__12235\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__12232\,
            I => \N__12228\
        );

    \I__2554\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12223\
        );

    \I__2553\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12223\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__12223\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4\
        );

    \I__2551\ : InMux
    port map (
            O => \N__12220\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__2550\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12214\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__12214\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__2548\ : InMux
    port map (
            O => \N__12211\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__2547\ : InMux
    port map (
            O => \N__12208\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__12205\,
            I => \N__12201\
        );

    \I__2545\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12196\
        );

    \I__2544\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12189\
        );

    \I__2543\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12189\
        );

    \I__2542\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12189\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__12196\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__12189\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12184\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\
        );

    \I__2538\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12178\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__12178\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__12175\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__2534\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12165\
        );

    \I__2533\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12161\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__12165\,
            I => \N__12158\
        );

    \I__2531\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12155\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__12161\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__12158\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__12155\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__2527\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12139\
        );

    \I__2526\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12139\
        );

    \I__2525\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12136\
        );

    \I__2524\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12126\
        );

    \I__2523\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12126\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__12139\,
            I => \N__12123\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__12136\,
            I => \N__12120\
        );

    \I__2520\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12115\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12115\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12112\
        );

    \I__2517\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12107\
        );

    \I__2516\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12107\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__12126\,
            I => \N__12102\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__12123\,
            I => \N__12102\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__12120\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__12115\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__12112\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__12107\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__12102\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__2508\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__12088\,
            I => \beamY_RNIQNF11_0Z0Z_8\
        );

    \I__2506\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12081\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__12084\,
            I => \N__12076\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__12081\,
            I => \N__12073\
        );

    \I__2503\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12069\
        );

    \I__2502\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12064\
        );

    \I__2501\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12064\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__12073\,
            I => \N__12061\
        );

    \I__2499\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12058\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__12069\,
            I => \beamY_i_2\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__12064\,
            I => \beamY_i_2\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__12061\,
            I => \beamY_i_2\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__12058\,
            I => \beamY_i_2\
        );

    \I__2494\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12045\
        );

    \I__2493\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__12045\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__12042\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12034\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12034\,
            I => \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4\
        );

    \I__2488\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12028\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__12028\,
            I => \N__12025\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__12025\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6\
        );

    \I__2485\ : InMux
    port map (
            O => \N__12022\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__2483\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12013\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__12013\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9\
        );

    \I__2481\ : InMux
    port map (
            O => \N__12010\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__2480\ : InMux
    port map (
            O => \N__12007\,
            I => \N__12004\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__12004\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__2478\ : InMux
    port map (
            O => \N__12001\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__2477\ : InMux
    port map (
            O => \N__11998\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__11995\,
            I => \N__11991\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11987\
        );

    \I__2474\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11982\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11982\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11987\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11982\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__11977\,
            I => \N__11974\
        );

    \I__2469\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11971\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__11971\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\
        );

    \I__2467\ : InMux
    port map (
            O => \N__11968\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11962\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__11962\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11959\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11956\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__11953\,
            I => \N__11948\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11938\
        );

    \I__2460\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11938\
        );

    \I__2459\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11938\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11938\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__11938\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11929\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__11929\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \N__11921\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11908\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11908\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11908\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11901\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11901\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11901\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11893\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11916\,
            I => \N__11893\
        );

    \I__2444\ : InMux
    port map (
            O => \N__11915\,
            I => \N__11890\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__11908\,
            I => \N__11887\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__11901\,
            I => \N__11884\
        );

    \I__2441\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11881\
        );

    \I__2440\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11876\
        );

    \I__2439\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11876\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11873\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__11890\,
            I => \N__11870\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__11887\,
            I => \N__11861\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__11884\,
            I => \N__11861\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__11881\,
            I => \N__11861\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__11876\,
            I => \N__11861\
        );

    \I__2432\ : Span4Mux_s2_v
    port map (
            O => \N__11873\,
            I => \N__11858\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__11870\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__11861\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__11858\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__11851\,
            I => \N__11848\
        );

    \I__2427\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__11845\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\
        );

    \I__2425\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11839\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__11839\,
            I => \beamY_RNIALEQZ0Z_9\
        );

    \I__2423\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11833\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__11833\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\
        );

    \I__2421\ : InMux
    port map (
            O => \N__11830\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\
        );

    \I__2420\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__11824\,
            I => \beamY_RNIALEQ_1Z0Z_9\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__11818\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\
        );

    \I__2416\ : InMux
    port map (
            O => \N__11815\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11807\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11804\
        );

    \I__2413\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11801\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__11807\,
            I => \N__11798\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__11804\,
            I => \N__11788\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__11801\,
            I => \N__11781\
        );

    \I__2409\ : Span4Mux_s2_v
    port map (
            O => \N__11798\,
            I => \N__11781\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11797\,
            I => \N__11774\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11774\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11774\
        );

    \I__2405\ : InMux
    port map (
            O => \N__11794\,
            I => \N__11765\
        );

    \I__2404\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11765\
        );

    \I__2403\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11765\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11765\
        );

    \I__2401\ : Span4Mux_s2_v
    port map (
            O => \N__11788\,
            I => \N__11762\
        );

    \I__2400\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11759\
        );

    \I__2399\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11756\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__11781\,
            I => \N__11753\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11746\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11746\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__11762\,
            I => \N__11746\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__11759\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__11756\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__11753\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__11746\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__2390\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11734\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__11734\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\
        );

    \I__2388\ : InMux
    port map (
            O => \N__11731\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__11728\,
            I => \N__11725\
        );

    \I__2386\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11722\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__11722\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11719\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__11716\,
            I => \N__11713\
        );

    \I__2382\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11710\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\
        );

    \I__2380\ : InMux
    port map (
            O => \N__11707\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__2379\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__11701\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\
        );

    \I__2377\ : InMux
    port map (
            O => \N__11698\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__2376\ : InMux
    port map (
            O => \N__11695\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__11692\,
            I => \N__11688\
        );

    \I__2374\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11678\
        );

    \I__2373\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11678\
        );

    \I__2372\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11678\
        );

    \I__2371\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11675\
        );

    \I__2370\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11672\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__11678\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__11675\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__11672\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__2366\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__11662\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921\
        );

    \I__2364\ : InMux
    port map (
            O => \N__11659\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__2362\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11650\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__11650\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\
        );

    \I__2360\ : InMux
    port map (
            O => \N__11647\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\
        );

    \I__2359\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11641\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__11641\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum1_4
        );

    \I__2357\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11635\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__11635\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum0_4
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__11632\,
            I => \un7_pixel_0_axb4_cascade_\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11625\
        );

    \I__2353\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11620\
        );

    \I__2352\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11620\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__11620\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum1_5
        );

    \I__2350\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11614\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__11614\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \N__11608\
        );

    \I__2347\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11605\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__11605\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__2345\ : InMux
    port map (
            O => \N__11602\,
            I => un4_pixel_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__2344\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__11593\,
            I => \N__11589\
        );

    \I__2341\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11586\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__11589\,
            I => un7_pixel_0_axb4
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__11586\,
            I => un7_pixel_0_axb4
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__2337\ : InMux
    port map (
            O => \N__11578\,
            I => \N__11575\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__11575\,
            I => \N__11572\
        );

    \I__2335\ : Odrv12
    port map (
            O => \N__11572\,
            I => if_generate_plus_mult1_un47_sum_m_2
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11563\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__11563\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__2331\ : InMux
    port map (
            O => \N__11560\,
            I => un4_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__11557\,
            I => \N__11553\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__11556\,
            I => \N__11550\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11545\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11545\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__11545\,
            I => un7_pixel_0_axb4_i
        );

    \I__2325\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__11539\,
            I => \un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__11536\,
            I => un4_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2322\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__11530\,
            I => \un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__2320\ : InMux
    port map (
            O => \N__11527\,
            I => un4_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2319\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11518\
        );

    \I__2317\ : Span4Mux_h
    port map (
            O => \N__11518\,
            I => \N__11512\
        );

    \I__2316\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11509\
        );

    \I__2315\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11506\
        );

    \I__2314\ : InMux
    port map (
            O => \N__11515\,
            I => \N__11503\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__11512\,
            I => un7_pixel_0_axb3
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__11509\,
            I => un7_pixel_0_axb3
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__11506\,
            I => un7_pixel_0_axb3
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__11503\,
            I => un7_pixel_0_axb3
        );

    \I__2309\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11488\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__11488\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum1_3
        );

    \I__2306\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__11482\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum0_3
        );

    \I__2304\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11476\,
            I => if_generate_plus_mult1_un47_sum_m_3
        );

    \I__2302\ : InMux
    port map (
            O => \N__11473\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2
        );

    \I__2301\ : InMux
    port map (
            O => \N__11470\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3
        );

    \I__2300\ : InMux
    port map (
            O => \N__11467\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4
        );

    \I__2299\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__11461\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum0_2
        );

    \I__2297\ : InMux
    port map (
            O => \N__11458\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1
        );

    \I__2296\ : InMux
    port map (
            O => \N__11455\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2
        );

    \I__2295\ : InMux
    port map (
            O => \N__11452\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3
        );

    \I__2294\ : InMux
    port map (
            O => \N__11449\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__11446\,
            I => \un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_\
        );

    \I__2292\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__11440\,
            I => g1_0_0_0_1
        );

    \I__2290\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11430\
        );

    \I__2289\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11427\
        );

    \I__2288\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11422\
        );

    \I__2287\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11422\
        );

    \I__2286\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11419\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__11430\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__11427\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__11422\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__11419\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__11410\,
            I => \g3_0_0_0_cascade_\
        );

    \I__2280\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11404\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__11404\,
            I => g1_4_0_0_0
        );

    \I__2278\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__11398\,
            I => \N_1869_0_0\
        );

    \I__2276\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N_1870_0_0\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__11389\,
            I => \font_un127_pixel_6_ns_1_0_0_cascade_\
        );

    \I__2273\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11380\
        );

    \I__2272\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11380\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__11380\,
            I => font_un13_pixel_0_1_0_0_22
        );

    \I__2270\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11374\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__11374\,
            I => \N__11371\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__11371\,
            I => \N_520\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__11368\,
            I => \N__11365\
        );

    \I__2266\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__11356\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__2261\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__11347\,
            I => \N__11344\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__11344\,
            I => \N__11341\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__11341\,
            I => \un4_pixel_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__2257\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11334\
        );

    \I__2256\ : SRMux
    port map (
            O => \N__11337\,
            I => \N__11331\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__11334\,
            I => \N__11328\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__11331\,
            I => \N__11325\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__11328\,
            I => \N__11322\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__11325\,
            I => \beamY_RNIJ0DBZ0Z_8\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__11322\,
            I => \beamY_RNIJ0DBZ0Z_8\
        );

    \I__2250\ : IoInMux
    port map (
            O => \N__11317\,
            I => \N__11314\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__11314\,
            I => \N__11310\
        );

    \I__2248\ : IoInMux
    port map (
            O => \N__11313\,
            I => \N__11307\
        );

    \I__2247\ : Span4Mux_s2_v
    port map (
            O => \N__11310\,
            I => \N__11304\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__11307\,
            I => \N__11301\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__11304\,
            I => \N__11298\
        );

    \I__2244\ : Span4Mux_s1_v
    port map (
            O => \N__11301\,
            I => \N__11295\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__11298\,
            I => \N__11292\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__11295\,
            I => \N__11289\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__11292\,
            I => \VSync_c\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__11289\,
            I => \VSync_c\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__2238\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11275\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__11275\,
            I => \un4_pixel_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11272\,
            I => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1
        );

    \I__2234\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__11266\,
            I => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__11263\,
            I => \N__11260\
        );

    \I__2231\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11256\
        );

    \I__2230\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11253\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__11256\,
            I => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__11253\,
            I => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0\
        );

    \I__2227\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11245\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__11245\,
            I => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321\
        );

    \I__2225\ : InMux
    port map (
            O => \N__11242\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__2224\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__11236\,
            I => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__11233\,
            I => \N__11229\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__11232\,
            I => \N__11226\
        );

    \I__2220\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11221\
        );

    \I__2219\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11221\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__11221\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__2217\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__11215\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__2215\ : InMux
    port map (
            O => \N__11212\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__2214\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11206\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__11206\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__2212\ : InMux
    port map (
            O => \N__11203\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \N__11196\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11192\
        );

    \I__2209\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11187\
        );

    \I__2208\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11187\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11192\,
            I => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__11187\,
            I => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11179\
        );

    \I__2204\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11176\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__11176\,
            I => \N__11173\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__11170\,
            I => un14_visibleylt9_0
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11161\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__11161\,
            I => un14_visibleylt4_0
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \un3_beamx_5_cascade_\
        );

    \I__2196\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11152\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11149\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__11146\,
            I => \N_324_0_0_0\
        );

    \I__2192\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11140\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__11140\,
            I => \N__11137\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__11137\,
            I => \N__11134\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__11134\,
            I => \N_303_0_0_0\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__11131\,
            I => \N__11125\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__11130\,
            I => \N__11120\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__11129\,
            I => \N__11116\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11113\
        );

    \I__2184\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11109\
        );

    \I__2183\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11106\
        );

    \I__2182\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11103\
        );

    \I__2181\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11100\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11095\
        );

    \I__2179\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11095\
        );

    \I__2178\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11092\
        );

    \I__2177\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11085\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__11109\,
            I => \N__11078\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__11106\,
            I => \N__11078\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__11103\,
            I => \N__11078\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11073\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__11095\,
            I => \N__11073\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__11092\,
            I => \N__11070\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11067\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11064\
        );

    \I__2168\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11061\
        );

    \I__2167\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11058\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11055\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__11078\,
            I => \N__11052\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__11073\,
            I => \N__11049\
        );

    \I__2163\ : Span12Mux_s7_h
    port map (
            O => \N__11070\,
            I => \N__11044\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__11067\,
            I => \N__11044\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__11064\,
            I => \beamYZ0Z_0\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__11061\,
            I => \beamYZ0Z_0\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__11058\,
            I => \beamYZ0Z_0\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__11055\,
            I => \beamYZ0Z_0\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__11052\,
            I => \beamYZ0Z_0\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__11049\,
            I => \beamYZ0Z_0\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__11044\,
            I => \beamYZ0Z_0\
        );

    \I__2154\ : InMux
    port map (
            O => \N__11029\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__2153\ : InMux
    port map (
            O => \N__11026\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__2152\ : InMux
    port map (
            O => \N__11023\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__2151\ : InMux
    port map (
            O => \N__11020\,
            I => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__11017\,
            I => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_\
        );

    \I__2149\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11011\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__11011\,
            I => font_un13_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__2147\ : InMux
    port map (
            O => \N__11008\,
            I => \N__11001\
        );

    \I__2146\ : InMux
    port map (
            O => \N__11007\,
            I => \N__10998\
        );

    \I__2145\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10993\
        );

    \I__2144\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10993\
        );

    \I__2143\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10988\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__11001\,
            I => \N__10982\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10979\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__10993\,
            I => \N__10976\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10973\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__10991\,
            I => \N__10970\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__10988\,
            I => \N__10966\
        );

    \I__2136\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10963\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10960\
        );

    \I__2134\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10957\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__10982\,
            I => \N__10952\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__10979\,
            I => \N__10952\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__10976\,
            I => \N__10947\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__10973\,
            I => \N__10947\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10942\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10942\
        );

    \I__2127\ : Odrv12
    port map (
            O => \N__10966\,
            I => \beamYZ0Z_7\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10963\,
            I => \beamYZ0Z_7\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10960\,
            I => \beamYZ0Z_7\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__10957\,
            I => \beamYZ0Z_7\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__10952\,
            I => \beamYZ0Z_7\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__10947\,
            I => \beamYZ0Z_7\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10942\,
            I => \beamYZ0Z_7\
        );

    \I__2120\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10919\
        );

    \I__2119\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10919\
        );

    \I__2118\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10916\
        );

    \I__2117\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10908\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__10919\,
            I => \N__10905\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__10916\,
            I => \N__10902\
        );

    \I__2114\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10899\
        );

    \I__2113\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10896\
        );

    \I__2112\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10893\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10888\
        );

    \I__2110\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10888\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__10908\,
            I => \N__10881\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__10905\,
            I => \N__10874\
        );

    \I__2107\ : Span4Mux_v
    port map (
            O => \N__10902\,
            I => \N__10874\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__10899\,
            I => \N__10871\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10864\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10864\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10864\
        );

    \I__2102\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10861\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10854\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10854\
        );

    \I__2099\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10854\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__10881\,
            I => \N__10851\
        );

    \I__2097\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10846\
        );

    \I__2096\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10846\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__10874\,
            I => \beamYZ0Z_9\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__10871\,
            I => \beamYZ0Z_9\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__10864\,
            I => \beamYZ0Z_9\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__10861\,
            I => \beamYZ0Z_9\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10854\,
            I => \beamYZ0Z_9\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__10851\,
            I => \beamYZ0Z_9\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__10846\,
            I => \beamYZ0Z_9\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__10831\,
            I => \N__10828\
        );

    \I__2087\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10825\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10822\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__10822\,
            I => un8_beamylto9_1
        );

    \I__2084\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10814\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10806\
        );

    \I__2082\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10806\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10803\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10800\
        );

    \I__2079\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10794\
        );

    \I__2078\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10794\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__10806\,
            I => \N__10788\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__10803\,
            I => \N__10788\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10800\,
            I => \N__10785\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10782\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10794\,
            I => \N__10778\
        );

    \I__2072\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10775\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__10788\,
            I => \N__10772\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__10785\,
            I => \N__10767\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__10782\,
            I => \N__10767\
        );

    \I__2068\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10764\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__10778\,
            I => \N__10761\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__10775\,
            I => \beamYZ0Z_8\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__10772\,
            I => \beamYZ0Z_8\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__10767\,
            I => \beamYZ0Z_8\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__10764\,
            I => \beamYZ0Z_8\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__10761\,
            I => \beamYZ0Z_8\
        );

    \I__2061\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10747\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__10744\,
            I => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0\
        );

    \I__2058\ : InMux
    port map (
            O => \N__10741\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__10738\,
            I => \un5_visibley_ac0_7_cascade_\
        );

    \I__2056\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10726\
        );

    \I__2055\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10726\
        );

    \I__2054\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10726\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__10723\,
            I => \N__10720\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__10720\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__10717\,
            I => \beamY_4_rep1_RNICDQEZ0_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10708\
        );

    \I__2048\ : InMux
    port map (
            O => \N__10713\,
            I => \N__10705\
        );

    \I__2047\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10700\
        );

    \I__2046\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10700\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__10708\,
            I => \beamY_fastZ0Z_3\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__10705\,
            I => \beamY_fastZ0Z_3\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__10700\,
            I => \beamY_fastZ0Z_3\
        );

    \I__2042\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10688\
        );

    \I__2041\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10685\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10682\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__10688\,
            I => \N__10677\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__10685\,
            I => \N__10674\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__10682\,
            I => \N__10671\
        );

    \I__2036\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10666\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10666\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__10677\,
            I => \N__10660\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__10674\,
            I => \N__10660\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__10671\,
            I => \N__10655\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10655\
        );

    \I__2030\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10652\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__10660\,
            I => un5_visibley_c2
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__10655\,
            I => un5_visibley_c2
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__10652\,
            I => un5_visibley_c2
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__10645\,
            I => \N__10642\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10638\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10635\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__10638\,
            I => un11_visibley
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__10635\,
            I => un11_visibley
        );

    \I__2021\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__10627\,
            I => \N__10624\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__10624\,
            I => un44
        );

    \I__2018\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10618\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__10618\,
            I => \Pixel_1_e_1\
        );

    \I__2016\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10607\
        );

    \I__2015\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10607\
        );

    \I__2014\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10602\
        );

    \I__2013\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10602\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__10607\,
            I => \beamY_fastZ0Z_2\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__10602\,
            I => \beamY_fastZ0Z_2\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__10597\,
            I => \N__10590\
        );

    \I__2009\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10587\
        );

    \I__2008\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10584\
        );

    \I__2007\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10579\
        );

    \I__2006\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10579\
        );

    \I__2005\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10576\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10587\,
            I => \beamY_4_repZ0Z1\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__10584\,
            I => \beamY_4_repZ0Z1\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__10579\,
            I => \beamY_4_repZ0Z1\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__10576\,
            I => \beamY_4_repZ0Z1\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10564\
        );

    \I__1999\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10561\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__10561\,
            I => \beamY_fast_RNIK8HHZ0Z_2\
        );

    \I__1997\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10549\
        );

    \I__1996\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10546\
        );

    \I__1995\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10540\
        );

    \I__1994\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10540\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__10554\,
            I => \N__10537\
        );

    \I__1992\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10534\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__10552\,
            I => \N__10529\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__10549\,
            I => \N__10523\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10520\
        );

    \I__1988\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10517\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10514\
        );

    \I__1986\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10511\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10508\
        );

    \I__1984\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10505\
        );

    \I__1983\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10500\
        );

    \I__1982\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10500\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10493\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10493\
        );

    \I__1979\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10493\
        );

    \I__1978\ : Odrv12
    port map (
            O => \N__10523\,
            I => \beamYZ0Z_6\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__10520\,
            I => \beamYZ0Z_6\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__10517\,
            I => \beamYZ0Z_6\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__10514\,
            I => \beamYZ0Z_6\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__10511\,
            I => \beamYZ0Z_6\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__10508\,
            I => \beamYZ0Z_6\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__10505\,
            I => \beamYZ0Z_6\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__10500\,
            I => \beamYZ0Z_6\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__10493\,
            I => \beamYZ0Z_6\
        );

    \I__1969\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10469\
        );

    \I__1968\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10466\
        );

    \I__1967\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10459\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__10469\,
            I => \N__10455\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10448\
        );

    \I__1964\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10445\
        );

    \I__1963\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10440\
        );

    \I__1962\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10440\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__10462\,
            I => \N__10436\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10432\
        );

    \I__1959\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10429\
        );

    \I__1958\ : Span12Mux_s6_v
    port map (
            O => \N__10455\,
            I => \N__10426\
        );

    \I__1957\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10423\
        );

    \I__1956\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10420\
        );

    \I__1955\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10417\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10414\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__10448\,
            I => \N__10411\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__10445\,
            I => \N__10406\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__10440\,
            I => \N__10406\
        );

    \I__1950\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10399\
        );

    \I__1949\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10399\
        );

    \I__1948\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10399\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__10432\,
            I => \beamYZ0Z_5\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__10429\,
            I => \beamYZ0Z_5\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__10426\,
            I => \beamYZ0Z_5\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__10423\,
            I => \beamYZ0Z_5\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__10420\,
            I => \beamYZ0Z_5\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__10417\,
            I => \beamYZ0Z_5\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__10414\,
            I => \beamYZ0Z_5\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__10411\,
            I => \beamYZ0Z_5\
        );

    \I__1939\ : Odrv12
    port map (
            O => \N__10406\,
            I => \beamYZ0Z_5\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__10399\,
            I => \beamYZ0Z_5\
        );

    \I__1937\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10375\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__10375\,
            I => \beamY_RNIKOP3Z0Z_7\
        );

    \I__1935\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10369\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__10369\,
            I => un42lt10
        );

    \I__1933\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10358\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10355\
        );

    \I__1931\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10348\
        );

    \I__1930\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10348\
        );

    \I__1929\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10348\
        );

    \I__1928\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10345\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__10358\,
            I => un5_visibley_c7
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10355\,
            I => un5_visibley_c7
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__10348\,
            I => un5_visibley_c7
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10345\,
            I => un5_visibley_c7
        );

    \I__1923\ : InMux
    port map (
            O => \N__10336\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1922\ : InMux
    port map (
            O => \N__10333\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__1921\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10324\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__10324\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__1918\ : InMux
    port map (
            O => \N__10321\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__1917\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__10315\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0\
        );

    \I__1915\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10308\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10305\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__10308\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__10305\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__10300\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_\
        );

    \I__1910\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__10294\,
            I => \Pixel_1_RNOZ0Z_19\
        );

    \I__1908\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10288\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__10288\,
            I => un1_visiblex_27
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__1905\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10279\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__10276\,
            I => \N__10273\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__10273\,
            I => un5_visibley_ac0_7
        );

    \I__1901\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10267\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__10267\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8\
        );

    \I__1899\ : InMux
    port map (
            O => \N__10264\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__10261\,
            I => \N__10258\
        );

    \I__1897\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10255\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__10255\,
            I => \N__10252\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__10252\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__10249\,
            I => \N__10244\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__10248\,
            I => \N__10240\
        );

    \I__1892\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10236\
        );

    \I__1891\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10227\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10227\
        );

    \I__1889\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10227\
        );

    \I__1888\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10227\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__10236\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__10227\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0\
        );

    \I__1885\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10219\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__10219\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\
        );

    \I__1883\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10213\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__10213\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\
        );

    \I__1881\ : InMux
    port map (
            O => \N__10210\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\
        );

    \I__1880\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__10204\,
            I => \Pixel_1_RNOZ0Z_18\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__10201\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__10195\,
            I => \N__10191\
        );

    \I__1875\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10188\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__10191\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10188\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf\
        );

    \I__1872\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10179\
        );

    \I__1871\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10176\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__10179\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__10176\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0\
        );

    \I__1868\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1867\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10165\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__10165\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0\
        );

    \I__1865\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10157\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__10161\,
            I => \N__10154\
        );

    \I__1863\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10141\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__10157\,
            I => \N__10130\
        );

    \I__1861\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10120\
        );

    \I__1860\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10117\
        );

    \I__1859\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10110\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10110\
        );

    \I__1857\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10110\
        );

    \I__1856\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10105\
        );

    \I__1855\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10105\
        );

    \I__1854\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10100\
        );

    \I__1853\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10100\
        );

    \I__1852\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10097\
        );

    \I__1851\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10092\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__10141\,
            I => \N__10089\
        );

    \I__1849\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10076\
        );

    \I__1848\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10076\
        );

    \I__1847\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10076\
        );

    \I__1846\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10071\
        );

    \I__1845\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10071\
        );

    \I__1844\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10068\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__10134\,
            I => \N__10065\
        );

    \I__1842\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10061\
        );

    \I__1841\ : Span4Mux_h
    port map (
            O => \N__10130\,
            I => \N__10058\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10053\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10053\
        );

    \I__1838\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10042\
        );

    \I__1837\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10042\
        );

    \I__1836\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10042\
        );

    \I__1835\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10042\
        );

    \I__1834\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10042\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10029\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10029\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10029\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__10105\,
            I => \N__10029\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10029\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__10097\,
            I => \N__10029\
        );

    \I__1827\ : InMux
    port map (
            O => \N__10096\,
            I => \N__10026\
        );

    \I__1826\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10023\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__10092\,
            I => \N__10018\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__10089\,
            I => \N__10018\
        );

    \I__1823\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10013\
        );

    \I__1822\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10013\
        );

    \I__1821\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10010\
        );

    \I__1820\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10007\
        );

    \I__1819\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10002\
        );

    \I__1818\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10002\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__9995\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__9995\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__10068\,
            I => \N__9995\
        );

    \I__1814\ : InMux
    port map (
            O => \N__10065\,
            I => \N__9992\
        );

    \I__1813\ : InMux
    port map (
            O => \N__10064\,
            I => \N__9989\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__9986\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__10058\,
            I => \N__9979\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__10053\,
            I => \N__9979\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__10042\,
            I => \N__9979\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__10029\,
            I => \N__9976\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__10026\,
            I => un43lto1
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10023\,
            I => un43lto1
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__10018\,
            I => un43lto1
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__10013\,
            I => un43lto1
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__10010\,
            I => un43lto1
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10007\,
            I => un43lto1
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__10002\,
            I => un43lto1
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__9995\,
            I => un43lto1
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__9992\,
            I => un43lto1
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__9989\,
            I => un43lto1
        );

    \I__1797\ : Odrv12
    port map (
            O => \N__9986\,
            I => un43lto1
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__9979\,
            I => un43lto1
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__9976\,
            I => un43lto1
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__9949\,
            I => \un43lto4_1_cascade_\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__9946\,
            I => \un43lt10_cascade_\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9940\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__9940\,
            I => \un1_beamY_26\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \N__9934\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__9931\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9928\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__9922\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9919\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__9916\,
            I => \N__9913\
        );

    \I__1782\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__9910\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3\
        );

    \I__1780\ : InMux
    port map (
            O => \N__9907\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__9904\,
            I => \N__9901\
        );

    \I__1778\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__9898\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9895\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9889\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__9889\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9886\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \N__9878\
        );

    \I__1771\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9873\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9864\
        );

    \I__1769\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9864\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9864\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9876\,
            I => \N__9864\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__9873\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9864\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5\
        );

    \I__1764\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__9856\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\
        );

    \I__1762\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9850\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__9850\,
            I => \N__9847\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__9847\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9844\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__9841\,
            I => \N__9838\
        );

    \I__1757\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9835\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__9835\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5\
        );

    \I__1755\ : InMux
    port map (
            O => \N__9832\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9829\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\
        );

    \I__1753\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9823\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__9823\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\
        );

    \I__1751\ : InMux
    port map (
            O => \N__9820\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__9817\,
            I => \N__9813\
        );

    \I__1749\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9804\
        );

    \I__1748\ : InMux
    port map (
            O => \N__9813\,
            I => \N__9804\
        );

    \I__1747\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9804\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9801\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__9804\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__9801\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__9796\,
            I => \N__9793\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9790\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9790\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9787\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__1739\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__9781\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__1736\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9772\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__9772\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9769\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__1733\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9763\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__9763\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\
        );

    \I__1731\ : InMux
    port map (
            O => \N__9760\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__9754\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__9751\,
            I => \N__9743\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__9750\,
            I => \N__9737\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__9749\,
            I => \N__9733\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__9748\,
            I => \N__9729\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__9747\,
            I => \N__9726\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__9746\,
            I => \N__9723\
        );

    \I__1722\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9718\
        );

    \I__1721\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9718\
        );

    \I__1720\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9715\
        );

    \I__1719\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9712\
        );

    \I__1718\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9709\
        );

    \I__1717\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9696\
        );

    \I__1716\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9696\
        );

    \I__1715\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9696\
        );

    \I__1714\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9696\
        );

    \I__1713\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9696\
        );

    \I__1712\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9696\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9718\,
            I => \N__9693\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__9715\,
            I => \N__9688\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__9712\,
            I => \N__9688\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9681\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__9696\,
            I => \N__9681\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__9693\,
            I => \N__9681\
        );

    \I__1705\ : Span4Mux_s2_v
    port map (
            O => \N__9688\,
            I => \N__9678\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__9681\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__9678\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \N__9670\
        );

    \I__1701\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__9667\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9657\
        );

    \I__1697\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9653\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9649\
        );

    \I__1695\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9646\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9643\
        );

    \I__1693\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9640\
        );

    \I__1692\ : Span4Mux_s3_h
    port map (
            O => \N__9649\,
            I => \N__9635\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__9646\,
            I => \N__9635\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__9643\,
            I => \N__9632\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__9640\,
            I => \N__9627\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__9635\,
            I => \N__9627\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__9632\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__9627\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1685\ : InMux
    port map (
            O => \N__9622\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\
        );

    \I__1684\ : InMux
    port map (
            O => \N__9619\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\
        );

    \I__1683\ : InMux
    port map (
            O => \N__9616\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__1682\ : InMux
    port map (
            O => \N__9613\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__1681\ : InMux
    port map (
            O => \N__9610\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__9607\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__1678\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__9598\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9591\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__9594\,
            I => \N__9587\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9583\
        );

    \I__1673\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9578\
        );

    \I__1672\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9578\
        );

    \I__1671\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9574\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__9583\,
            I => \N__9569\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9569\
        );

    \I__1668\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9566\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9574\,
            I => \N__9561\
        );

    \I__1666\ : Span4Mux_h
    port map (
            O => \N__9569\,
            I => \N__9556\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__9566\,
            I => \N__9556\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__9565\,
            I => \N__9553\
        );

    \I__1663\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9550\
        );

    \I__1662\ : Span4Mux_s2_v
    port map (
            O => \N__9561\,
            I => \N__9547\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__9556\,
            I => \N__9544\
        );

    \I__1660\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9541\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__9550\,
            I => \N__9538\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__9547\,
            I => \N__9535\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__9544\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__9541\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__9538\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__9535\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__1652\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9520\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__9520\,
            I => \N__9517\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__9517\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__1649\ : InMux
    port map (
            O => \N__9514\,
            I => un4_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__1648\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9508\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9505\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__9505\,
            I => \un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9502\,
            I => un4_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__1644\ : InMux
    port map (
            O => \N__9499\,
            I => un4_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1643\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9468\
        );

    \I__1642\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9468\
        );

    \I__1641\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9468\
        );

    \I__1640\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9468\
        );

    \I__1639\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9465\
        );

    \I__1638\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9460\
        );

    \I__1637\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9460\
        );

    \I__1636\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9447\
        );

    \I__1635\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9447\
        );

    \I__1634\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9447\
        );

    \I__1633\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9447\
        );

    \I__1632\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9447\
        );

    \I__1631\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9447\
        );

    \I__1630\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9434\
        );

    \I__1629\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9434\
        );

    \I__1628\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9434\
        );

    \I__1627\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9434\
        );

    \I__1626\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9415\
        );

    \I__1625\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9415\
        );

    \I__1624\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9415\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9412\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9403\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__9460\,
            I => \N__9400\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__9447\,
            I => \N__9397\
        );

    \I__1619\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9388\
        );

    \I__1618\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9388\
        );

    \I__1617\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9388\
        );

    \I__1616\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9388\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9385\
        );

    \I__1614\ : InMux
    port map (
            O => \N__9433\,
            I => \N__9372\
        );

    \I__1613\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9372\
        );

    \I__1612\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9372\
        );

    \I__1611\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9372\
        );

    \I__1610\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9372\
        );

    \I__1609\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9372\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9369\
        );

    \I__1607\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9361\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9361\
        );

    \I__1605\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9354\
        );

    \I__1604\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9354\
        );

    \I__1603\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9354\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__9415\,
            I => \N__9349\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__9412\,
            I => \N__9349\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9336\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9336\
        );

    \I__1598\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9336\
        );

    \I__1597\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9336\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9336\
        );

    \I__1595\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9336\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__9403\,
            I => \N__9331\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__9400\,
            I => \N__9331\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__9397\,
            I => \N__9328\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__9388\,
            I => \N__9319\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__9385\,
            I => \N__9319\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9319\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__9369\,
            I => \N__9319\
        );

    \I__1587\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9316\
        );

    \I__1586\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9311\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9311\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__9361\,
            I => un7_pixel_1_axb3
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__9354\,
            I => un7_pixel_1_axb3
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__9349\,
            I => un7_pixel_1_axb3
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__9336\,
            I => un7_pixel_1_axb3
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__9331\,
            I => un7_pixel_1_axb3
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__9328\,
            I => un7_pixel_1_axb3
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__9319\,
            I => un7_pixel_1_axb3
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__9316\,
            I => un7_pixel_1_axb3
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__9311\,
            I => un7_pixel_1_axb3
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__9292\,
            I => \un7_pixel_1_axb3_cascade_\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__9289\,
            I => \N__9280\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__9288\,
            I => \N__9273\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9256\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__9286\,
            I => \N__9248\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9238\
        );

    \I__1569\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9238\
        );

    \I__1568\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9238\
        );

    \I__1567\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9238\
        );

    \I__1566\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9229\
        );

    \I__1565\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9229\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9229\
        );

    \I__1563\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9229\
        );

    \I__1562\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9220\
        );

    \I__1561\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9220\
        );

    \I__1560\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9220\
        );

    \I__1559\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9220\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__9269\,
            I => \N__9213\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__9268\,
            I => \N__9208\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__9267\,
            I => \N__9205\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__9266\,
            I => \N__9201\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__9265\,
            I => \N__9198\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__9264\,
            I => \N__9194\
        );

    \I__1552\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9189\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9189\
        );

    \I__1550\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9184\
        );

    \I__1549\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9184\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__9259\,
            I => \N__9177\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__9256\,
            I => \N__9173\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9170\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9157\
        );

    \I__1544\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9157\
        );

    \I__1543\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9157\
        );

    \I__1542\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9157\
        );

    \I__1541\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9157\
        );

    \I__1540\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9157\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9150\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__9229\,
            I => \N__9150\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9150\
        );

    \I__1536\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9137\
        );

    \I__1535\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9137\
        );

    \I__1534\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9137\
        );

    \I__1533\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9137\
        );

    \I__1532\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9137\
        );

    \I__1531\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9137\
        );

    \I__1530\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9134\
        );

    \I__1529\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9129\
        );

    \I__1528\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9129\
        );

    \I__1527\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9118\
        );

    \I__1526\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9118\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9118\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9118\
        );

    \I__1523\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9118\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9113\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9113\
        );

    \I__1520\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9110\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9105\
        );

    \I__1518\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9105\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9098\
        );

    \I__1516\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9098\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9098\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__9173\,
            I => un7_pixel_1_axb1
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__9170\,
            I => un7_pixel_1_axb1
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__9157\,
            I => un7_pixel_1_axb1
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__9150\,
            I => un7_pixel_1_axb1
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__9137\,
            I => un7_pixel_1_axb1
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__9134\,
            I => un7_pixel_1_axb1
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__9129\,
            I => un7_pixel_1_axb1
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__9118\,
            I => un7_pixel_1_axb1
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__9113\,
            I => un7_pixel_1_axb1
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__9110\,
            I => un7_pixel_1_axb1
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__9105\,
            I => un7_pixel_1_axb1
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__9098\,
            I => un7_pixel_1_axb1
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__9073\,
            I => \N__9070\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9067\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__9067\,
            I => \N_532_i\
        );

    \I__1499\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__9061\,
            I => un117_pixel_2_6_i3_mux
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__9058\,
            I => \N__9047\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9044\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__9056\,
            I => \N__9041\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__9055\,
            I => \N__9036\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__9054\,
            I => \N__9033\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \N__9021\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__9052\,
            I => \N__9013\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__9051\,
            I => \N__9007\
        );

    \I__1489\ : InMux
    port map (
            O => \N__9050\,
            I => \N__8998\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9047\,
            I => \N__8998\
        );

    \I__1487\ : InMux
    port map (
            O => \N__9044\,
            I => \N__8998\
        );

    \I__1486\ : InMux
    port map (
            O => \N__9041\,
            I => \N__8998\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__9040\,
            I => \N__8992\
        );

    \I__1484\ : InMux
    port map (
            O => \N__9039\,
            I => \N__8980\
        );

    \I__1483\ : InMux
    port map (
            O => \N__9036\,
            I => \N__8980\
        );

    \I__1482\ : InMux
    port map (
            O => \N__9033\,
            I => \N__8980\
        );

    \I__1481\ : InMux
    port map (
            O => \N__9032\,
            I => \N__8980\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__9031\,
            I => \N__8977\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__9030\,
            I => \N__8973\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__9029\,
            I => \N__8970\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9028\,
            I => \N__8958\
        );

    \I__1476\ : InMux
    port map (
            O => \N__9027\,
            I => \N__8958\
        );

    \I__1475\ : InMux
    port map (
            O => \N__9026\,
            I => \N__8958\
        );

    \I__1474\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8958\
        );

    \I__1473\ : InMux
    port map (
            O => \N__9024\,
            I => \N__8953\
        );

    \I__1472\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8953\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__8947\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__9019\,
            I => \N__8944\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__9018\,
            I => \N__8939\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \N__8933\
        );

    \I__1467\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8928\
        );

    \I__1466\ : InMux
    port map (
            O => \N__9013\,
            I => \N__8928\
        );

    \I__1465\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8925\
        );

    \I__1464\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8918\
        );

    \I__1463\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8918\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8918\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__8998\,
            I => \N__8915\
        );

    \I__1460\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8902\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8902\
        );

    \I__1458\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8902\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8902\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8902\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8902\
        );

    \I__1454\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8899\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8980\,
            I => \N__8896\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8881\
        );

    \I__1451\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8881\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8881\
        );

    \I__1449\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8881\
        );

    \I__1448\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8881\
        );

    \I__1447\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8881\
        );

    \I__1446\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8881\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8876\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8876\
        );

    \I__1443\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8873\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__8951\,
            I => \N__8869\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8864\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8855\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8855\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8855\
        );

    \I__1437\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8855\
        );

    \I__1436\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8844\
        );

    \I__1435\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8844\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8844\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8844\
        );

    \I__1432\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8844\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__8928\,
            I => \N__8831\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__8925\,
            I => \N__8831\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8831\
        );

    \I__1428\ : Span4Mux_h
    port map (
            O => \N__8915\,
            I => \N__8831\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8831\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__8899\,
            I => \N__8831\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__8896\,
            I => \N__8822\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__8881\,
            I => \N__8822\
        );

    \I__1423\ : Span4Mux_v
    port map (
            O => \N__8876\,
            I => \N__8822\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8822\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8815\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8815\
        );

    \I__1419\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8815\
        );

    \I__1418\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8812\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8864\,
            I => un7_pixel_1_axb2
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__8855\,
            I => un7_pixel_1_axb2
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__8844\,
            I => un7_pixel_1_axb2
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__8831\,
            I => un7_pixel_1_axb2
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__8822\,
            I => un7_pixel_1_axb2
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8815\,
            I => un7_pixel_1_axb2
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__8812\,
            I => un7_pixel_1_axb2
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__8797\,
            I => \N__8793\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8779\
        );

    \I__1408\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8776\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__8792\,
            I => \N__8771\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__8791\,
            I => \N__8767\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8755\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8755\
        );

    \I__1403\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8746\
        );

    \I__1402\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8746\
        );

    \I__1401\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8746\
        );

    \I__1400\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8746\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \N__8743\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__8783\,
            I => \N__8740\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__8782\,
            I => \N__8736\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__8779\,
            I => \N__8731\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__8776\,
            I => \N__8728\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__8775\,
            I => \N__8723\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__8774\,
            I => \N__8720\
        );

    \I__1392\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8710\
        );

    \I__1391\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8710\
        );

    \I__1390\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8710\
        );

    \I__1389\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8710\
        );

    \I__1388\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8701\
        );

    \I__1387\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8701\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8701\
        );

    \I__1385\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8701\
        );

    \I__1384\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8683\
        );

    \I__1383\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8683\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__8755\,
            I => \N__8680\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8677\
        );

    \I__1380\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8668\
        );

    \I__1379\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8668\
        );

    \I__1378\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8668\
        );

    \I__1377\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8668\
        );

    \I__1376\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8663\
        );

    \I__1375\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8663\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__8731\,
            I => \N__8658\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__8728\,
            I => \N__8658\
        );

    \I__1372\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8647\
        );

    \I__1371\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8647\
        );

    \I__1370\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8647\
        );

    \I__1369\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8647\
        );

    \I__1368\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8647\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__8710\,
            I => \N__8642\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__8701\,
            I => \N__8642\
        );

    \I__1365\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8639\
        );

    \I__1364\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8624\
        );

    \I__1363\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8624\
        );

    \I__1362\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8624\
        );

    \I__1361\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8624\
        );

    \I__1360\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8624\
        );

    \I__1359\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8624\
        );

    \I__1358\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8624\
        );

    \I__1357\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8613\
        );

    \I__1356\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8613\
        );

    \I__1355\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8613\
        );

    \I__1354\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8613\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8613\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8610\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__8680\,
            I => \un4_pixel_N_3\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__8677\,
            I => \un4_pixel_N_3\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__8668\,
            I => \un4_pixel_N_3\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__8663\,
            I => \un4_pixel_N_3\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__8658\,
            I => \un4_pixel_N_3\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__8647\,
            I => \un4_pixel_N_3\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__8642\,
            I => \un4_pixel_N_3\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__8639\,
            I => \un4_pixel_N_3\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__8624\,
            I => \un4_pixel_N_3\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__8613\,
            I => \un4_pixel_N_3\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__8610\,
            I => \un4_pixel_N_3\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__8587\,
            I => \Pixel_1_RNOZ0Z_73_cascade_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__8581\,
            I => \Pixel_1_RNOZ0Z_72\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__8578\,
            I => \N__8564\
        );

    \I__1336\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8556\
        );

    \I__1335\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8556\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__8575\,
            I => \N__8553\
        );

    \I__1333\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8549\
        );

    \I__1332\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8544\
        );

    \I__1331\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8544\
        );

    \I__1330\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8541\
        );

    \I__1329\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8536\
        );

    \I__1328\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8536\
        );

    \I__1327\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8533\
        );

    \I__1326\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8528\
        );

    \I__1325\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8528\
        );

    \I__1324\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8523\
        );

    \I__1323\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8518\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8518\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8511\
        );

    \I__1320\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8505\
        );

    \I__1319\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8505\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__8549\,
            I => \N__8502\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__8544\,
            I => \N__8491\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8491\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8491\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8491\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8491\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8486\
        );

    \I__1311\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8486\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__8523\,
            I => \N__8481\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8481\
        );

    \I__1308\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8476\
        );

    \I__1307\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8476\
        );

    \I__1306\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8471\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8471\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__8511\,
            I => \N__8468\
        );

    \I__1303\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8465\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8462\
        );

    \I__1301\ : Span4Mux_h
    port map (
            O => \N__8502\,
            I => \N__8455\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__8491\,
            I => \N__8455\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__8486\,
            I => \N__8455\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__8481\,
            I => \N__8448\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__8476\,
            I => \N__8448\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__8471\,
            I => \N__8448\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__8468\,
            I => \N__8443\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8443\
        );

    \I__1293\ : Span4Mux_h
    port map (
            O => \N__8462\,
            I => \N__8440\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__8455\,
            I => \N__8437\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__8448\,
            I => \N__8434\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__8443\,
            I => font_un36_pixel_23
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__8440\,
            I => font_un36_pixel_23
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__8437\,
            I => font_un36_pixel_23
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__8434\,
            I => font_un36_pixel_23
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__8425\,
            I => \Pixel_1_RNOZ0Z_48_cascade_\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__8419\,
            I => \N_234_0_0\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1281\ : Span4Mux_h
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__8407\,
            I => \d_N_3_0_0\
        );

    \I__1279\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8398\
        );

    \I__1278\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8398\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__8398\,
            I => un7_pixel_0_axb3_i
        );

    \I__1276\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__8392\,
            I => \N_326_0_0\
        );

    \I__1274\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__8386\,
            I => g0_18_1
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N_321_0_cascade_\
        );

    \I__1271\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__8377\,
            I => \N_314_0_0_0\
        );

    \I__1269\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__8368\,
            I => \N_328_0_0_0\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__8365\,
            I => \g1_2_0_0_cascade_\
        );

    \I__1265\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8359\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8354\
        );

    \I__1263\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8351\
        );

    \I__1262\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8348\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__8354\,
            I => \N_192_0_1\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__8351\,
            I => \N_192_0_1\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__8348\,
            I => \N_192_0_1\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__8341\,
            I => \un117_pixel_6_1_0_1_4_cascade_\
        );

    \I__1257\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N_219_0_0_1\
        );

    \I__1255\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8326\
        );

    \I__1254\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8326\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__8326\,
            I => un7_pixel_1_axb3_i
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__8323\,
            I => \N__8320\
        );

    \I__1251\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8314\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__8314\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__1248\ : InMux
    port map (
            O => \N__8311\,
            I => un4_pixel_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__8308\,
            I => \N_1482_0_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__1245\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__8299\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__1243\ : InMux
    port map (
            O => \N__8296\,
            I => un4_pixel_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1241\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__8284\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__1238\ : InMux
    port map (
            O => \N__8281\,
            I => un4_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__1237\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__8275\,
            I => \un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8272\,
            I => un4_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__1234\ : InMux
    port map (
            O => \N__8269\,
            I => un4_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__8266\,
            I => \un7_pixel_1_axb2_cascade_\
        );

    \I__1232\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8257\
        );

    \I__1231\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8257\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__8257\,
            I => un7_pixel_1_axb2_i
        );

    \I__1229\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__8251\,
            I => \Pixel_1_RNOZ0Z_44\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__8248\,
            I => \N_305_0_cascade_\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__8245\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_\
        );

    \I__1225\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__8239\,
            I => \Pixel_1_RNOZ0Z_82\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__8236\,
            I => \font_un127_pixel_m_4_1_1_cascade_\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__8230\,
            I => font_un127_pixel_m_4_1
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__8227\,
            I => \un7_pixel_1_c4_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__8218\,
            I => font_un127_pixel_m_7_1_0
        );

    \I__1216\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__8209\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__1213\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8202\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__8205\,
            I => \N__8199\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8192\
        );

    \I__1210\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8189\
        );

    \I__1209\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8186\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8183\
        );

    \I__1207\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8178\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8178\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__8192\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__8189\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__8186\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__8183\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__8178\,
            I => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__8158\,
            I => \N_307_0_0_1\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__8155\,
            I => \font_un13_pixel_0_1_0_0_22_cascade_\
        );

    \I__1195\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8148\
        );

    \I__1194\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8145\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__8148\,
            I => \N__8142\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__8145\,
            I => \beamY_RNIVV787O2Z0Z_2\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__8142\,
            I => \beamY_RNIVV787O2Z0Z_2\
        );

    \I__1190\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8134\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8131\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__8131\,
            I => \Pixel_1_RNOZ0Z_47\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__8128\,
            I => \N__8125\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N_338_0_0_0\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \font_un127_pixel_m_cascade_\
        );

    \I__1183\ : IoInMux
    port map (
            O => \N__8116\,
            I => \N__8113\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__8113\,
            I => \N__8110\
        );

    \I__1181\ : IoSpan4Mux
    port map (
            O => \N__8110\,
            I => \N__8106\
        );

    \I__1180\ : IoInMux
    port map (
            O => \N__8109\,
            I => \N__8103\
        );

    \I__1179\ : Span4Mux_s0_v
    port map (
            O => \N__8106\,
            I => \N__8100\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8097\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__1176\ : Span4Mux_s3_v
    port map (
            O => \N__8097\,
            I => \N__8091\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__8094\,
            I => \N__8085\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__8091\,
            I => \N__8085\
        );

    \I__1173\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8082\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__8085\,
            I => \Pixel_c\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__8082\,
            I => \Pixel_c\
        );

    \I__1170\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__8074\,
            I => font_un127_pixel_m_4
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \g0_0_1_cascade_\
        );

    \I__1167\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1165\ : Span4Mux_h
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__8059\,
            I => font_un69_pixellto3
        );

    \I__1163\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__8053\,
            I => g0_0_2
        );

    \I__1161\ : InMux
    port map (
            O => \N__8050\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__1160\ : InMux
    port map (
            O => \N__8047\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__8044\,
            I => \N__8040\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__8043\,
            I => \N__8037\
        );

    \I__1157\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8032\
        );

    \I__1156\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8032\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__8032\,
            I => font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__1154\ : InMux
    port map (
            O => \N__8029\,
            I => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1153\ : InMux
    port map (
            O => \N__8026\,
            I => \N__8023\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__8023\,
            I => \N__8019\
        );

    \I__1151\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8016\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__8019\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__8016\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1147\ : InMux
    port map (
            O => \N__8008\,
            I => \N__8005\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__8002\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__7999\,
            I => \beamY_fastZ0Z_8\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7992\
        );

    \I__1142\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7989\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__7992\,
            I => \N__7986\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7989\,
            I => \beamY_fast_RNIG57DZ0Z_8\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__7986\,
            I => \beamY_fast_RNIG57DZ0Z_8\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__7981\,
            I => \beamY_fast_RNIG57DZ0Z_8_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__7975\,
            I => \N__7969\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7966\
        );

    \I__1134\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7961\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7961\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__7969\,
            I => un5_visibley_c6_0_1
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7966\,
            I => un5_visibley_c6_0_1
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__7961\,
            I => un5_visibley_c6_0_1
        );

    \I__1129\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7950\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7947\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7944\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__7947\,
            I => \N__7941\
        );

    \I__1125\ : Odrv12
    port map (
            O => \N__7944\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__7941\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7933\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__7933\,
            I => \N__7930\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__7930\,
            I => \N__7926\
        );

    \I__1120\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7923\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__7926\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__7923\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7914\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7911\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7914\,
            I => \N__7908\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7911\,
            I => \N__7905\
        );

    \I__1113\ : Odrv12
    port map (
            O => \N__7908\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__7905\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__7900\,
            I => \N__7895\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__7899\,
            I => \N__7892\
        );

    \I__1109\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7885\
        );

    \I__1108\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7885\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7882\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7876\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7873\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__7885\,
            I => \N__7868\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7882\,
            I => \N__7865\
        );

    \I__1102\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7860\
        );

    \I__1101\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7860\
        );

    \I__1100\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7857\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__7876\,
            I => \N__7854\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__7873\,
            I => \N__7850\
        );

    \I__1097\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7845\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7845\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__7868\,
            I => \N__7842\
        );

    \I__1094\ : Span4Mux_v
    port map (
            O => \N__7865\,
            I => \N__7837\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__7860\,
            I => \N__7837\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7832\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__7854\,
            I => \N__7832\
        );

    \I__1090\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7829\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__7850\,
            I => \beamYZ0Z_4\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__7845\,
            I => \beamYZ0Z_4\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__7842\,
            I => \beamYZ0Z_4\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__7837\,
            I => \beamYZ0Z_4\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__7832\,
            I => \beamYZ0Z_4\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__7829\,
            I => \beamYZ0Z_4\
        );

    \I__1083\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7812\
        );

    \I__1082\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7804\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__7812\,
            I => \N__7801\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7798\
        );

    \I__1079\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7795\
        );

    \I__1078\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7788\
        );

    \I__1077\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7788\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7788\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__7804\,
            I => \N__7779\
        );

    \I__1074\ : Span4Mux_h
    port map (
            O => \N__7801\,
            I => \N__7779\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__7798\,
            I => \N__7772\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__7795\,
            I => \N__7772\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__7788\,
            I => \N__7772\
        );

    \I__1070\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7763\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7763\
        );

    \I__1068\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7763\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7763\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__7779\,
            I => \beamY_RNI9DLCZ0Z_0\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__7772\,
            I => \beamY_RNI9DLCZ0Z_0\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__7763\,
            I => \beamY_RNI9DLCZ0Z_0\
        );

    \I__1063\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7749\
        );

    \I__1062\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7749\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__7754\,
            I => \N__7746\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__7749\,
            I => \N__7743\
        );

    \I__1059\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7740\
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__7743\,
            I => \un21_beamy_cry_3_c_RNIERZ0Z93\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7740\,
            I => \un21_beamy_cry_3_c_RNIERZ0Z93\
        );

    \I__1056\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7732\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__7732\,
            I => \N__7728\
        );

    \I__1054\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7725\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__7728\,
            I => \N__7720\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__7725\,
            I => \N__7720\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__7720\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__1050\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7714\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__7714\,
            I => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0
        );

    \I__1048\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7707\
        );

    \I__1047\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7704\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__7707\,
            I => \beamY_fastZ0Z_7\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__7704\,
            I => \beamY_fastZ0Z_7\
        );

    \I__1044\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7691\
        );

    \I__1042\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7687\
        );

    \I__1041\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7684\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__7691\,
            I => \N__7681\
        );

    \I__1039\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7678\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__7687\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__7684\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__7681\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__7678\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1034\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7666\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__7663\,
            I => \N__7658\
        );

    \I__1031\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7655\
        );

    \I__1030\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7652\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__7658\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__7655\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7652\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1026\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__7642\,
            I => \N__7639\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__7639\,
            I => un11_visibleylto9_4
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__7636\,
            I => \beamY_fast_RNI198KZ0Z_2_cascade_\
        );

    \I__1022\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__7630\,
            I => \N__7627\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__7627\,
            I => font_un127_pixel_m_1
        );

    \I__1019\ : InMux
    port map (
            O => \N__7624\,
            I => un21_beamy_cry_6
        );

    \I__1018\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7615\
        );

    \I__1017\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7615\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__7615\,
            I => \un21_beamy_cry_7_c_RNIM7EZ0Z3\
        );

    \I__1015\ : InMux
    port map (
            O => \N__7612\,
            I => un21_beamy_cry_7
        );

    \I__1014\ : InMux
    port map (
            O => \N__7609\,
            I => \bfn_6_4_0_\
        );

    \I__1013\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1012\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7600\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__7600\,
            I => \un21_beamy_cry_8_c_RNIOAFZ0Z3\
        );

    \I__1010\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7593\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__7596\,
            I => \N__7589\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7582\
        );

    \I__1007\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7579\
        );

    \I__1006\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7576\
        );

    \I__1005\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7573\
        );

    \I__1004\ : InMux
    port map (
            O => \N__7587\,
            I => \N__7568\
        );

    \I__1003\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7568\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7563\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__7582\,
            I => \N__7558\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7558\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7555\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7550\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7550\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__7567\,
            I => \N__7546\
        );

    \I__995\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7543\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__7563\,
            I => \N__7540\
        );

    \I__993\ : Span4Mux_v
    port map (
            O => \N__7558\,
            I => \N__7537\
        );

    \I__992\ : Span4Mux_h
    port map (
            O => \N__7555\,
            I => \N__7532\
        );

    \I__991\ : Span4Mux_v
    port map (
            O => \N__7550\,
            I => \N__7532\
        );

    \I__990\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7527\
        );

    \I__989\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7527\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__7543\,
            I => \beamYZ0Z_3\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__7540\,
            I => \beamYZ0Z_3\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__7537\,
            I => \beamYZ0Z_3\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__7532\,
            I => \beamYZ0Z_3\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__7527\,
            I => \beamYZ0Z_3\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__7516\,
            I => \N__7512\
        );

    \I__982\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7505\
        );

    \I__981\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7505\
        );

    \I__980\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7498\
        );

    \I__979\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7498\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7494\
        );

    \I__977\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7491\
        );

    \I__976\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7488\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__7498\,
            I => \N__7483\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__7497\,
            I => \N__7479\
        );

    \I__973\ : Span4Mux_v
    port map (
            O => \N__7494\,
            I => \N__7472\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__7491\,
            I => \N__7472\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__7488\,
            I => \N__7472\
        );

    \I__970\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7467\
        );

    \I__969\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7467\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__7483\,
            I => \N__7463\
        );

    \I__967\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7458\
        );

    \I__966\ : InMux
    port map (
            O => \N__7479\,
            I => \N__7458\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__7472\,
            I => \N__7455\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__7467\,
            I => \N__7452\
        );

    \I__963\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7449\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__7463\,
            I => \N__7446\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__7458\,
            I => \N__7443\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__7455\,
            I => \N__7438\
        );

    \I__959\ : Span4Mux_h
    port map (
            O => \N__7452\,
            I => \N__7438\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__7449\,
            I => \beamYZ0Z_2\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__7446\,
            I => \beamYZ0Z_2\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__7443\,
            I => \beamYZ0Z_2\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__7438\,
            I => \beamYZ0Z_2\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__953\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__7423\,
            I => un11_visibleylto9_1
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__7420\,
            I => \N_309_0_cascade_\
        );

    \I__950\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7414\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N_316_0\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__7411\,
            I => \N_323_0_cascade_\
        );

    \I__947\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__7405\,
            I => \N_302_0_0_0\
        );

    \I__945\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__7396\,
            I => \N__7393\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__7393\,
            I => \N_5_0_0_0\
        );

    \I__941\ : InMux
    port map (
            O => \N__7390\,
            I => un21_beamy_cry_1
        );

    \I__940\ : InMux
    port map (
            O => \N__7387\,
            I => un21_beamy_cry_2
        );

    \I__939\ : InMux
    port map (
            O => \N__7384\,
            I => un21_beamy_cry_3
        );

    \I__938\ : InMux
    port map (
            O => \N__7381\,
            I => un21_beamy_cry_4
        );

    \I__937\ : InMux
    port map (
            O => \N__7378\,
            I => un21_beamy_cry_5
        );

    \I__936\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7372\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__7372\,
            I => g0_40_1
        );

    \I__934\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__932\ : Odrv12
    port map (
            O => \N__7363\,
            I => \N_206\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__7360\,
            I => \g0_6_1_1_cascade_\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__7357\,
            I => \g0_6_1_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7350\
        );

    \I__928\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7347\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N_192_0_0\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__7347\,
            I => \N_192_0_0\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__7342\,
            I => \g1_3_1_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__7333\,
            I => \N__7330\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__7330\,
            I => g1_3
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__7327\,
            I => \g0_10_1_cascade_\
        );

    \I__919\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7321\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__7321\,
            I => if_generate_plus_mult1_un75_sum_cry_2_s
        );

    \I__917\ : InMux
    port map (
            O => \N__7318\,
            I => un4_pixel_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__7315\,
            I => \N__7312\
        );

    \I__915\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7309\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7309\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__913\ : InMux
    port map (
            O => \N__7306\,
            I => un4_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__912\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__7300\,
            I => \un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__910\ : InMux
    port map (
            O => \N__7297\,
            I => un4_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__909\ : InMux
    port map (
            O => \N__7294\,
            I => un4_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__7291\,
            I => \un7_pixel_1_axb1_cascade_\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__7288\,
            I => \N_203_0_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7282\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N_268_0\
        );

    \I__904\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__7276\,
            I => m3_0
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__7273\,
            I => \Pixel_1_RNOZ0Z_69_cascade_\
        );

    \I__901\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7267\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__7267\,
            I => \Pixel_1_RNOZ0Z_70\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__7264\,
            I => \g0_35_1_cascade_\
        );

    \I__898\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7258\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__7258\,
            I => \un115_pixel_13_15___m1_e_0Z0Z_1\
        );

    \I__896\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7252\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7252\,
            I => \un115_pixel_13_15__i2_mux\
        );

    \I__894\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__7246\,
            I => \d_N_6_0\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__7243\,
            I => \N__7240\
        );

    \I__891\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N_6\
        );

    \I__889\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7231\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__7231\,
            I => \N_5_i_0\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__7228\,
            I => \g1_0_0_cascade_\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__7225\,
            I => \N_250_0_cascade_\
        );

    \I__885\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__7219\,
            I => \N_266_0\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__7216\,
            I => \N_242_0_cascade_\
        );

    \I__882\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7210\,
            I => \Pixel_1_RNOZ0Z_61\
        );

    \I__880\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7204\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N_282\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__7201\,
            I => \font_un127_pixel_1_1_cascade_\
        );

    \I__877\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7195\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N_336_0\
        );

    \I__875\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__7189\,
            I => un5_beamx_6
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__7186\,
            I => \N__7183\
        );

    \I__872\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7179\
        );

    \I__871\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7176\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7179\,
            I => un8_beamy_3
        );

    \I__869\ : LocalMux
    port map (
            O => \N__7176\,
            I => un8_beamy_3
        );

    \I__868\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__7168\,
            I => g1_1
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__7165\,
            I => \N_283_cascade_\
        );

    \I__865\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7159\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__7159\,
            I => \N_285\
        );

    \I__863\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__7153\,
            I => font_un13_pixel_23
        );

    \I__861\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__7147\,
            I => font_un73_pixellt7_0
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__7144\,
            I => \font_un13_pixel_23_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__7138\,
            I => \Pixel_1_RNOZ0Z_60\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__7135\,
            I => \Pixel_1_RNOZ0Z_39_cascade_\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__7132\,
            I => \N__7128\
        );

    \I__854\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7123\
        );

    \I__853\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7123\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7123\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0
        );

    \I__851\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7117\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__7117\,
            I => \beamY_RNIF8TM3Z0Z_9\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__7114\,
            I => \beamY_RNIVD444Z0Z_9_cascade_\
        );

    \I__848\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__7110\,
            I => \N__7100\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__7109\,
            I => \N__7096\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__7108\,
            I => \N__7093\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7090\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__7104\,
            I => \N__7087\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__7103\,
            I => \N__7083\
        );

    \I__841\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7080\
        );

    \I__840\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7073\
        );

    \I__839\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7073\
        );

    \I__838\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7073\
        );

    \I__837\ : Span4Mux_h
    port map (
            O => \N__7090\,
            I => \N__7070\
        );

    \I__836\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7063\
        );

    \I__835\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7063\
        );

    \I__834\ : InMux
    port map (
            O => \N__7083\,
            I => \N__7063\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__7080\,
            I => \beamY_RNIGBU92Z0Z_9\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__7073\,
            I => \beamY_RNIGBU92Z0Z_9\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__7070\,
            I => \beamY_RNIGBU92Z0Z_9\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__7063\,
            I => \beamY_RNIGBU92Z0Z_9\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__7054\,
            I => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_\
        );

    \I__828\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__7048\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \N_7_0_0_0_cascade_\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__7042\,
            I => \un8_beamy_3_cascade_\
        );

    \I__824\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7036\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__7036\,
            I => \Pixel_1_RNOZ0Z_43\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__7033\,
            I => \N__7030\
        );

    \I__821\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__7027\,
            I => \Pixel_1_RNOZ0Z_42\
        );

    \I__819\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__7018\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__7015\,
            I => \beamY_RNI9I1Q6Z0Z_9_cascade_\
        );

    \I__815\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7000\
        );

    \I__814\ : InMux
    port map (
            O => \N__7011\,
            I => \N__7000\
        );

    \I__813\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7000\
        );

    \I__812\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7000\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__7000\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3
        );

    \I__810\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__6994\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0
        );

    \I__808\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6982\
        );

    \I__807\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6982\
        );

    \I__806\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6982\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6974\
        );

    \I__804\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6963\
        );

    \I__803\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6963\
        );

    \I__802\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6963\
        );

    \I__801\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6963\
        );

    \I__800\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6963\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__6974\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6963\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__797\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6941\
        );

    \I__796\ : InMux
    port map (
            O => \N__6957\,
            I => \N__6941\
        );

    \I__795\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6941\
        );

    \I__794\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6941\
        );

    \I__793\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6941\
        );

    \I__792\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6936\
        );

    \I__791\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6936\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__6941\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6936\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_\
        );

    \I__787\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__6925\,
            I => \beamY_RNIQQREO1Z0Z_3\
        );

    \I__785\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6914\
        );

    \I__784\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6914\
        );

    \I__783\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6909\
        );

    \I__782\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6909\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__6914\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_c5
        );

    \I__780\ : LocalMux
    port map (
            O => \N__6909\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_c5
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__778\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6893\
        );

    \I__777\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6893\
        );

    \I__776\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6888\
        );

    \I__775\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6888\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__6893\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2
        );

    \I__773\ : LocalMux
    port map (
            O => \N__6888\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__6883\,
            I => \N__6878\
        );

    \I__771\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6875\
        );

    \I__770\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6870\
        );

    \I__769\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6870\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6867\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6870\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1
        );

    \I__766\ : Odrv4
    port map (
            O => \N__6867\,
            I => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1
        );

    \I__765\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6858\
        );

    \I__764\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6855\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__6858\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6
        );

    \I__762\ : LocalMux
    port map (
            O => \N__6855\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6
        );

    \I__761\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6847\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__6847\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0
        );

    \I__759\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6841\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6841\,
            I => \beamY_4_rep1_RNI9H1FZ0Z1\
        );

    \I__757\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6835\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__6832\,
            I => \beamY_RNIHS041Z0Z_6\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__6829\,
            I => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_\
        );

    \I__753\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6822\
        );

    \I__752\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6819\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__6822\,
            I => \beamY_fastZ0Z_4\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__6819\,
            I => \beamY_fastZ0Z_4\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__6814\,
            I => \N__6809\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__6813\,
            I => \N__6806\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__6812\,
            I => \N__6803\
        );

    \I__746\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6800\
        );

    \I__745\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6796\
        );

    \I__744\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6793\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__6800\,
            I => \N__6790\
        );

    \I__742\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6787\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__6796\,
            I => \beamY_fastZ0Z_9\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__6793\,
            I => \beamY_fastZ0Z_9\
        );

    \I__739\ : Odrv4
    port map (
            O => \N__6790\,
            I => \beamY_fastZ0Z_9\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__6787\,
            I => \beamY_fastZ0Z_9\
        );

    \I__737\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6775\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__6775\,
            I => \beamY_fast_RNICEGAZ0Z_4\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__6772\,
            I => \N__6768\
        );

    \I__734\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6757\
        );

    \I__733\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6757\
        );

    \I__732\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6757\
        );

    \I__731\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6757\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__6757\,
            I => font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_\
        );

    \I__728\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6748\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__6748\,
            I => \N__6741\
        );

    \I__726\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6736\
        );

    \I__725\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6736\
        );

    \I__724\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6731\
        );

    \I__723\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6731\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__6741\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i
        );

    \I__721\ : LocalMux
    port map (
            O => \N__6736\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i
        );

    \I__720\ : LocalMux
    port map (
            O => \N__6731\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i
        );

    \I__719\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6721\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__6721\,
            I => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__6718\,
            I => \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_\
        );

    \I__716\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__6712\,
            I => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__6709\,
            I => \font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_\
        );

    \I__713\ : InMux
    port map (
            O => \N__6706\,
            I => \N__6703\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N_208_0_0_1\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__6700\,
            I => \N_1260_0_0_1_cascade_\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__6697\,
            I => \Z_decfrac2_1_0_0_0_cascade_\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__6694\,
            I => \un115_pixel_3_0_3__N_8_0_0_0_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__6688\,
            I => un117_pixel_3_1_0_1_4
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__6685\,
            I => \m4_cascade_\
        );

    \I__705\ : InMux
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__6676\,
            I => \Pixel_1_RNOZ0Z_88\
        );

    \I__702\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6670\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__6670\,
            I => \Pixel_1_RNOZ0Z_63\
        );

    \I__700\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6664\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__6664\,
            I => \un115_pixel_2_0_5__N_14\
        );

    \I__698\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6655\
        );

    \I__697\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6655\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__6655\,
            I => \G_370\
        );

    \I__695\ : InMux
    port map (
            O => \N__6652\,
            I => un4_pixel_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \un4_pixel_N_3_cascade_\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__692\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__6640\,
            I => \un4_pixel_if_generate_plus_mult1_un75_sum_iZ0\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__6637\,
            I => \g0_3_1_cascade_\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__6634\,
            I => \un115_pixel_0_a2_0_cascade_\
        );

    \I__688\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N_281\
        );

    \I__686\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__6622\,
            I => \N_231\
        );

    \I__684\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__6616\,
            I => \Pixel_1_RNOZ0Z_62\
        );

    \I__682\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__6610\,
            I => \N_275_0\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__679\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__6601\,
            I => \un115_pixel_13_15__m3_a0Z0Z_0\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__6598\,
            I => \un115_pixel_13_15__m3_a0Z0Z_0_cascade_\
        );

    \I__676\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N_215_0\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__6589\,
            I => \Pixel_1_RNOZ0Z_66_cascade_\
        );

    \I__673\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__6583\,
            I => un117_pixel_3_1_3
        );

    \I__671\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6576\
        );

    \I__670\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6573\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N_234_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__6573\,
            I => \N_234_0\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \m3_0_cascade_\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__6565\,
            I => \un115_pixel_2_0_5__N_9_cascade_\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__664\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__662\ : Span4Mux_h
    port map (
            O => \N__6553\,
            I => \N__6549\
        );

    \I__661\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6546\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__6549\,
            I => un4_beamylt6
        );

    \I__659\ : LocalMux
    port map (
            O => \N__6546\,
            I => un4_beamylt6
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__6541\,
            I => \un4_beamylt8_0_cascade_\
        );

    \I__657\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__6535\,
            I => un1_beamylto9_0
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__6532\,
            I => \un1_beamylto9_3_cascade_\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \un5_beamx_4_cascade_\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__6526\,
            I => \un117_pixel_6_ns_1_3_cascade_\
        );

    \I__652\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N_192_0\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__6517\,
            I => \N_192_0_cascade_\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__6514\,
            I => \beamY_RNI1G0FH2_0Z0Z_3_cascade_\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cascade_\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__6508\,
            I => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_\
        );

    \I__646\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__6502\,
            I => \N__6499\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__6499\,
            I => \beamY_RNICCIKUQ_0Z0Z_3\
        );

    \I__643\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6488\
        );

    \I__641\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6483\
        );

    \I__640\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6483\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__6488\,
            I => \N__6476\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6476\
        );

    \I__637\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6473\
        );

    \I__636\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6470\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__6476\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__634\ : LocalMux
    port map (
            O => \N__6473\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6470\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__632\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6456\
        );

    \I__630\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6453\
        );

    \I__629\ : Span4Mux_s3_h
    port map (
            O => \N__6456\,
            I => \N__6449\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6446\
        );

    \I__627\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6443\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__6449\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__625\ : Odrv4
    port map (
            O => \N__6446\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__624\ : LocalMux
    port map (
            O => \N__6443\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__623\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__622\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6430\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6426\
        );

    \I__620\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6423\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__6426\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_c5
        );

    \I__618\ : LocalMux
    port map (
            O => \N__6423\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_c5
        );

    \I__617\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6414\
        );

    \I__616\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6411\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__6414\,
            I => \N__6408\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__6411\,
            I => \N__6402\
        );

    \I__613\ : Span4Mux_s3_h
    port map (
            O => \N__6408\,
            I => \N__6399\
        );

    \I__612\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6392\
        );

    \I__611\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6392\
        );

    \I__610\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6392\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__6402\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__608\ : Odrv4
    port map (
            O => \N__6399\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__607\ : LocalMux
    port map (
            O => \N__6392\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__606\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6382\,
            I => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__6379\,
            I => \font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_\
        );

    \I__603\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__6373\,
            I => \N__6368\
        );

    \I__601\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6363\
        );

    \I__600\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6363\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__6368\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__598\ : LocalMux
    port map (
            O => \N__6363\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__597\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__6352\,
            I => \beamY_RNICCIKUQZ0Z_3\
        );

    \I__594\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__6346\,
            I => \beamY_RNIIDGN6_0Z0Z_7\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__6343\,
            I => \beamY_RNIIDGN6Z0Z_7_cascade_\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__6340\,
            I => \beamY_RNIPM0M5Z0Z_9_cascade_\
        );

    \I__590\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__6334\,
            I => \beamY_RNIPM0M5_0Z0Z_9\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__587\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6319\
        );

    \I__586\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6319\
        );

    \I__585\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6319\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__6316\,
            I => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__6313\,
            I => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_\
        );

    \I__581\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6301\
        );

    \I__580\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6301\
        );

    \I__579\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6301\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__6298\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__6295\,
            I => \beamY_RNI1G0FH2Z0Z_3_cascade_\
        );

    \I__575\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6286\
        );

    \I__574\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6286\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__6286\,
            I => font_un36_pixel_if_generate_plus_mult1_un68_sum_c4
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__6283\,
            I => \N__6279\
        );

    \I__571\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6271\
        );

    \I__570\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6271\
        );

    \I__569\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6271\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__6271\,
            I => \beamY_RNIUAN5CR1Z0Z_3\
        );

    \I__567\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__566\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6262\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__6262\,
            I => font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i
        );

    \I__564\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__6256\,
            I => \beamY_fast_RNIEGGAZ0Z_6\
        );

    \I__562\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__6250\,
            I => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__6247\,
            I => \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__6244\,
            I => \beamY_RNIGBU92Z0Z_9_cascade_\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__6241\,
            I => \beamY_RNIQ8RJCCZ0Z_3_cascade_\
        );

    \I__557\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__6235\,
            I => \beamY_RNIQ8RJCC_0Z0Z_3\
        );

    \I__555\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6229\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__6229\,
            I => \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__6226\,
            I => \font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6220\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__6220\,
            I => \beamY_RNI03RTE5Z0Z_4\
        );

    \I__550\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__6214\,
            I => \beamY_RNI03RTE5_0Z0Z_4\
        );

    \I__548\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__6208\,
            I => \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i\
        );

    \I__546\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6196\
        );

    \I__545\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6196\
        );

    \I__544\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6196\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__6196\,
            I => font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__6193\,
            I => \Pixel_1_RNOZ0Z_34_cascade_\
        );

    \I__541\ : IoInMux
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6184\
        );

    \I__539\ : IoSpan4Mux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__6181\,
            I => \Clock12MHz_c\
        );

    \I__537\ : IoInMux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__535\ : Span4Mux_s1_h
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__534\ : Span4Mux_h
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__6166\,
            I => \N__6163\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__6163\,
            I => \Clock50MHz.PixelClock\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__6160\,
            I => \font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_7_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6178\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \beamX_RNI5457_0_5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__13333\,
            GLOBALBUFFEROUTPUT => un3_beamx_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \beamY_RNI03RTE5_4_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6990\,
            in1 => \N__6327\,
            in2 => \N__7900\,
            in3 => \N__6309\,
            lcout => \beamY_RNI03RTE5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILAPCPC_3_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__6492\,
            in1 => \N__6376\,
            in2 => \N__7596\,
            in3 => \N__6417\,
            lcout => \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6IISE5_3_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__6989\,
            in1 => \N__6308\,
            in2 => \_gnd_net_\,
            in3 => \N__6326\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ8RJCC_0_3_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100011110"
        )
    port map (
            in0 => \N__6491\,
            in1 => \N__9577\,
            in2 => \N__6160\,
            in3 => \N__6459\,
            lcout => \beamY_RNIQ8RJCC_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI03RTE5_0_4_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6310\,
            in1 => \N__7898\,
            in2 => \N__6331\,
            in3 => \N__6991\,
            lcout => \beamY_RNI03RTE5_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ8RJCC_3_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6496\,
            in1 => \N__6463\,
            in2 => \N__9594\,
            in3 => \N__6203\,
            lcout => OPEN,
            ltout => \beamY_RNIQ8RJCCZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFVNMRT_3_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6418\,
            in2 => \N__6241\,
            in3 => \N__6238\,
            lcout => OPEN,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4J28J12_3_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__6552\,
            in1 => \N__6232\,
            in2 => \N__6226\,
            in3 => \N__6211\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFA02UM_4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6223\,
            in1 => \N__6217\,
            in2 => \_gnd_net_\,
            in3 => \N__6435\,
            lcout => \font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7592\,
            lcout => un4_beamylt6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIH479FH_3_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111010100"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__6436\,
            in2 => \N__9664\,
            in3 => \N__6205\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un68_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUAN5CR1_3_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__6358\,
            in2 => \_gnd_net_\,
            in3 => \N__6505\,
            lcout => \beamY_RNIUAN5CR1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_34_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6268\,
            in1 => \_gnd_net_\,
            in2 => \N__6283\,
            in3 => \N__6292\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_15_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__7515\,
            in1 => \N__7597\,
            in2 => \N__6193\,
            in3 => \N__6282\,
            lcout => font_un69_pixellto3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBH9OEE_2_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6291\,
            in1 => \N__6278\,
            in2 => \N__7516\,
            in3 => \N__6267\,
            lcout => font_un36_pixel_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7549\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_3_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101010101"
        )
    port map (
            in0 => \N__10474\,
            in1 => \N__7486\,
            in2 => \N__7567\,
            in3 => \N__7891\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIEGGA_6_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__10473\,
            in1 => \N__10781\,
            in2 => \N__6814\,
            in3 => \N__7699\,
            lcout => \beamY_fast_RNIEGGAZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNITAOJ_5_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__6778\,
            in1 => \N__11007\,
            in2 => \N__6813\,
            in3 => \N__7669\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4OJ_8_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10799\,
            in1 => \N__6259\,
            in2 => \_gnd_net_\,
            in3 => \N__10691\,
            lcout => OPEN,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGBU92_9_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111110"
        )
    port map (
            in0 => \N__6253\,
            in1 => \N__6715\,
            in2 => \N__6247\,
            in3 => \N__10887\,
            lcout => \beamY_RNIGBU92Z0Z_9\,
            ltout => \beamY_RNIGBU92Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIDGN6_0_7_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100001001"
        )
    port map (
            in0 => \N__10733\,
            in1 => \N__6766\,
            in2 => \N__6244\,
            in3 => \N__11791\,
            lcout => \beamY_RNIIDGN6_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPM0M5_0_9_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__11793\,
            in1 => \N__7086\,
            in2 => \N__6772\,
            in3 => \N__11918\,
            lcout => \beamY_RNIPM0M5_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIDGN6_7_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__10734\,
            in1 => \N__6767\,
            in2 => \N__7103\,
            in3 => \N__11792\,
            lcout => OPEN,
            ltout => \beamY_RNIIDGN6Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIF0K9E_7_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6349\,
            in2 => \N__6343\,
            in3 => \N__11920\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un47_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPM0M5_9_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100101101100"
        )
    port map (
            in0 => \N__11919\,
            in1 => \N__6771\,
            in2 => \N__7104\,
            in3 => \N__11794\,
            lcout => OPEN,
            ltout => \beamY_RNIPM0M5Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM948D_7_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10735\,
            in2 => \N__6340\,
            in3 => \N__6337\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPTUH72_3_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__6746\,
            in1 => \N__6955\,
            in2 => \N__9746\,
            in3 => \N__7009\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII319A3_3_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101110110010"
        )
    port map (
            in0 => \N__9564\,
            in1 => \N__9736\,
            in2 => \N__6313\,
            in3 => \N__6981\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQT00H2_3_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000011100"
        )
    port map (
            in0 => \N__6980\,
            in1 => \N__6958\,
            in2 => \N__9749\,
            in3 => \N__7010\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5VCS42_3_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010011"
        )
    port map (
            in0 => \N__6957\,
            in1 => \N__6747\,
            in2 => \N__9750\,
            in3 => \N__6861\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1G0FH2_3_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101100101"
        )
    port map (
            in0 => \N__6978\,
            in1 => \N__6956\,
            in2 => \N__9748\,
            in3 => \N__6745\,
            lcout => OPEN,
            ltout => \beamY_RNI1G0FH2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIF9EJC4_3_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__7012\,
            in1 => \N__9732\,
            in2 => \N__6295\,
            in3 => \N__6979\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1G0FH2_0_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001010110"
        )
    port map (
            in0 => \N__6977\,
            in1 => \N__6954\,
            in2 => \N__9747\,
            in3 => \N__6744\,
            lcout => OPEN,
            ltout => \beamY_RNI1G0FH2_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRD1F25_3_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__7011\,
            in1 => \_gnd_net_\,
            in2 => \N__6514\,
            in3 => \N__6928\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM3H2_3_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11006\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7587\,
            lcout => un1_beamylto9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_3_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__7586\,
            in1 => \N__7880\,
            in2 => \_gnd_net_\,
            in3 => \N__7503\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum\,
            ltout => \un1_beamY_if_generate_plus_mult1_un61_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGM5MH6_3_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001001101"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__6724\,
            in2 => \N__6511\,
            in3 => \N__6481\,
            lcout => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11\,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICCIKUQ_0_3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6407\,
            in1 => \N__6372\,
            in2 => \N__6508\,
            in3 => \N__6429\,
            lcout => \beamY_RNICCIKUQ_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIF4A60C_3_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__6482\,
            in1 => \N__6405\,
            in2 => \N__9565\,
            in3 => \N__6452\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un61_sum_c5,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICCIKUQ_3_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6406\,
            in1 => \N__6385\,
            in2 => \N__6379\,
            in3 => \N__6371\,
            lcout => \beamY_RNICCIKUQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_4_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7881\,
            in1 => \N__10557\,
            in2 => \N__6562\,
            in3 => \N__10472\,
            lcout => OPEN,
            ltout => \un4_beamylt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_8_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__10914\,
            in1 => \N__11005\,
            in2 => \N__6541\,
            in3 => \N__10813\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVGA6_2_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__10140\,
            in1 => \N__6538\,
            in2 => \N__7899\,
            in3 => \N__7511\,
            lcout => OPEN,
            ltout => \un1_beamylto9_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0DB_8_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10818\,
            in1 => \N__7182\,
            in2 => \N__6532\,
            in3 => \N__10927\,
            lcout => \beamY_RNIJ0DBZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEIP3_8_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10139\,
            in1 => \N__7588\,
            in2 => \_gnd_net_\,
            in3 => \N__10817\,
            lcout => OPEN,
            ltout => \un5_beamx_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2BJ7_2_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7510\,
            in1 => \N__11008\,
            in2 => \N__6529\,
            in3 => \N__10926\,
            lcout => un5_beamx_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_68_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__10135\,
            in1 => \N__6579\,
            in2 => \_gnd_net_\,
            in3 => \N__6523\,
            lcout => OPEN,
            ltout => \un117_pixel_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_43_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101001010011"
        )
    port map (
            in0 => \N__10138\,
            in1 => \N__8510\,
            in2 => \N__6526\,
            in3 => \N__6595\,
            lcout => \Pixel_1_RNOZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_i_11_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000000000"
        )
    port map (
            in0 => \N__9276\,
            in1 => \N__8766\,
            in2 => \N__9054\,
            in3 => \N__9481\,
            lcout => \N_192_0\,
            ltout => \N_192_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_67_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__10064\,
            in1 => \_gnd_net_\,
            in2 => \N__6517\,
            in3 => \N__6682\,
            lcout => un117_pixel_3_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_i_9_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010000000"
        )
    port map (
            in0 => \N__9278\,
            in1 => \N__8770\,
            in2 => \N__9055\,
            in3 => \N__9482\,
            lcout => \N_215_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_66_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001000"
        )
    port map (
            in0 => \N__9483\,
            in1 => \N__9039\,
            in2 => \N__8792\,
            in3 => \N__9279\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_66_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_42_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011100110"
        )
    port map (
            in0 => \N__10136\,
            in1 => \N__8552\,
            in2 => \N__6589\,
            in3 => \N__6586\,
            lcout => \Pixel_1_RNOZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un117_pixel_3_7_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100011101011"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__10137\,
            in2 => \N__8575\,
            in3 => \N__6580\,
            lcout => \N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_0_5_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010001000"
        )
    port map (
            in0 => \N__9480\,
            in1 => \N__9032\,
            in2 => \N__8791\,
            in3 => \N__9277\,
            lcout => \N_234_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__m3_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000000100"
        )
    port map (
            in0 => \N__8762\,
            in1 => \N__9270\,
            in2 => \N__9056\,
            in3 => \N__9493\,
            lcout => m3_0,
            ltout => \m3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_60_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10083\,
            in2 => \N__6568\,
            in3 => \N__6613\,
            lcout => \Pixel_1_RNOZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_2_0_5__m8_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011100000111"
        )
    port map (
            in0 => \N__8764\,
            in1 => \N__9272\,
            in2 => \N__9058\,
            in3 => \N__9495\,
            lcout => OPEN,
            ltout => \un115_pixel_2_0_5__N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_64_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__10085\,
            in1 => \N__6625\,
            in2 => \N__6565\,
            in3 => \N__8514\,
            lcout => OPEN,
            ltout => \g0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_40_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__10084\,
            in1 => \N__6619\,
            in2 => \N__6637\,
            in3 => \N__6673\,
            lcout => \d_N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_53_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000100010101"
        )
    port map (
            in0 => \N__9496\,
            in1 => \N__9050\,
            in2 => \N__9288\,
            in3 => \N__8765\,
            lcout => font_un73_pixellt7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_0_a2_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010000000"
        )
    port map (
            in0 => \N__8763\,
            in1 => \N__9271\,
            in2 => \N__9057\,
            in3 => \N__9494\,
            lcout => OPEN,
            ltout => \un115_pixel_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un117_pixel_2_7_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8515\,
            in2 => \N__6634\,
            in3 => \N__6667\,
            lcout => \N_281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_1_0_a2_5_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000010000000"
        )
    port map (
            in0 => \N__8697\,
            in1 => \N__9217\,
            in2 => \N__9030\,
            in3 => \N__9488\,
            lcout => \N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_62_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011111101101"
        )
    port map (
            in0 => \N__9219\,
            in1 => \N__8976\,
            in2 => \N__6607\,
            in3 => \N__8698\,
            lcout => \Pixel_1_RNOZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_86_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010000000"
        )
    port map (
            in0 => \N__8696\,
            in1 => \N__9216\,
            in2 => \N__9029\,
            in3 => \N__9487\,
            lcout => \N_275_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_70_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9486\,
            in1 => \N__8969\,
            in2 => \_gnd_net_\,
            in3 => \N__8695\,
            lcout => \Pixel_1_RNOZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__m3_a0_0_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8952\,
            in2 => \_gnd_net_\,
            in3 => \N__9484\,
            lcout => \un115_pixel_13_15__m3_a0Z0Z_0\,
            ltout => \un115_pixel_13_15__m3_a0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_88_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111011101"
        )
    port map (
            in0 => \N__9212\,
            in1 => \N__8967\,
            in2 => \N__6598\,
            in3 => \N__8693\,
            lcout => \Pixel_1_RNOZ0Z_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_63_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111111"
        )
    port map (
            in0 => \N__8699\,
            in1 => \N__9218\,
            in2 => \N__9031\,
            in3 => \N__9489\,
            lcout => \Pixel_1_RNOZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_2_0_5__m13_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000100010"
        )
    port map (
            in0 => \N__9485\,
            in1 => \N__8968\,
            in2 => \N__9269\,
            in3 => \N__8694\,
            lcout => \un115_pixel_2_0_5__N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_cry_1_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13057\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un82_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6660\,
            in2 => \N__6646\,
            in3 => \N__9176\,
            lcout => \G_370\,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un82_sum_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_cry_3_c_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7324\,
            in2 => \N__9259\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_cry_4_c_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6661\,
            in2 => \N__7315\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_s_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7303\,
            in2 => \_gnd_net_\,
            in3 => \N__6652\,
            lcout => \un4_pixel_N_3\,
            ltout => \un4_pixel_N_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_74_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9024\,
            in1 => \N__9180\,
            in2 => \N__6649\,
            in3 => \N__9491\,
            lcout => \N_208_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_i_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14092\,
            lcout => \un4_pixel_if_generate_plus_mult1_un75_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__g0_0_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000000000"
        )
    port map (
            in0 => \N__9211\,
            in1 => \N__8700\,
            in2 => \N__9053\,
            in3 => \N__9490\,
            lcout => \N_192_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_75_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111010100"
        )
    port map (
            in0 => \N__10124\,
            in1 => \N__7375\,
            in2 => \N__8783\,
            in3 => \N__9027\,
            lcout => OPEN,
            ltout => \N_1260_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_49_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__6706\,
            in1 => \N__10126\,
            in2 => \N__6700\,
            in3 => \N__8576\,
            lcout => \N_307_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_78_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9263\,
            in1 => \N__9028\,
            in2 => \N__8784\,
            in3 => \N__9479\,
            lcout => OPEN,
            ltout => \Z_decfrac2_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_51_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111010001"
        )
    port map (
            in0 => \N__6691\,
            in1 => \N__8577\,
            in2 => \N__6697\,
            in3 => \N__10127\,
            lcout => \N_303_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_3_0_3__g0_0_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011010000010"
        )
    port map (
            in0 => \N__9262\,
            in1 => \N__9025\,
            in2 => \N__8782\,
            in3 => \N__9477\,
            lcout => OPEN,
            ltout => \un115_pixel_3_0_3__N_8_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_79_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10123\,
            in2 => \N__6694\,
            in3 => \N__8357\,
            lcout => un117_pixel_3_1_0_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_3_0_3__m4_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8739\,
            in1 => \N__9026\,
            in2 => \_gnd_net_\,
            in3 => \N__9478\,
            lcout => OPEN,
            ltout => \m4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_59_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10125\,
            in2 => \N__6685\,
            in3 => \N__7353\,
            lcout => \N_316_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_8_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7620\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13221\,
            ce => \N__13274\,
            sr => \_gnd_net_\
        );

    \beamY_fast_8_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13221\,
            ce => \N__13274\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7929\,
            in2 => \_gnd_net_\,
            in3 => \N__7810\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13221\,
            ce => \N__13274\,
            sr => \_gnd_net_\
        );

    \beamY_fast_4_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__7808\,
            in1 => \_gnd_net_\,
            in2 => \N__7754\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13218\,
            ce => \N__13272\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIRPUB_4_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6799\,
            in1 => \N__6825\,
            in2 => \_gnd_net_\,
            in3 => \N__7662\,
            lcout => OPEN,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIT5511_6_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__7717\,
            in1 => \N__10692\,
            in2 => \N__6718\,
            in3 => \N__7695\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_9_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7606\,
            in2 => \_gnd_net_\,
            in3 => \N__7809\,
            lcout => \beamY_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13218\,
            ce => \N__13272\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7605\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13218\,
            ce => \N__13272\,
            sr => \_gnd_net_\
        );

    \beamY_RNIFIHM2_9_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__12132\,
            in2 => \N__11926\,
            in3 => \N__10363\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC4JRL_9_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11797\,
            in1 => \N__6898\,
            in2 => \N__6709\,
            in3 => \N__6919\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNICEGA_4_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__6826\,
            in1 => \N__10992\,
            in2 => \N__6812\,
            in3 => \N__10553\,
            lcout => \beamY_fast_RNICEGAZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIF1IR4_9_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11795\,
            in1 => \N__11924\,
            in2 => \N__7108\,
            in3 => \N__12135\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4DUR1_9_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__12131\,
            in2 => \_gnd_net_\,
            in3 => \N__10362\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKOS54_9_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000001111"
        )
    port map (
            in0 => \N__10364\,
            in1 => \N__10886\,
            in2 => \N__7109\,
            in3 => \N__12134\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIL92Q3_9_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11925\,
            in1 => \N__7099\,
            in2 => \_gnd_net_\,
            in3 => \N__11796\,
            lcout => OPEN,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7L40P_9_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6882\,
            in1 => \N__6899\,
            in2 => \N__6754\,
            in3 => \N__6920\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5VCS42_0_3_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001011001"
        )
    port map (
            in0 => \N__6751\,
            in1 => \N__6953\,
            in2 => \N__9751\,
            in3 => \N__6862\,
            lcout => \font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_4_rep1_RNI9H1F1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000001"
        )
    port map (
            in0 => \N__12145\,
            in1 => \N__10454\,
            in2 => \N__10554\,
            in3 => \N__10596\,
            lcout => \beamY_4_rep1_RNI9H1FZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9I1Q6_9_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__6850\,
            in1 => \N__10913\,
            in2 => \N__7110\,
            in3 => \N__10365\,
            lcout => OPEN,
            ltout => \beamY_RNI9I1Q6Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI035HO_9_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__10198\,
            in1 => \N__7024\,
            in2 => \N__7015\,
            in3 => \N__7051\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8L6E21_9_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6997\,
            in1 => \N__6881\,
            in2 => \N__6904\,
            in3 => \N__6922\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQQREO1_3_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__6952\,
            in1 => \_gnd_net_\,
            in2 => \N__6931\,
            in3 => \N__9742\,
            lcout => \beamY_RNIQQREO1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHS041_6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__10533\,
            in1 => \N__10453\,
            in2 => \_gnd_net_\,
            in3 => \N__12144\,
            lcout => \beamY_RNIHS041Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC4JRL_0_9_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010110"
        )
    port map (
            in0 => \N__6921\,
            in1 => \N__6900\,
            in2 => \N__6883\,
            in3 => \N__11787\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__11090\,
            in2 => \_gnd_net_\,
            in3 => \N__13294\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFHKL3_7_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101000"
        )
    port map (
            in0 => \N__7131\,
            in1 => \N__10986\,
            in2 => \N__10285\,
            in3 => \N__10532\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5D1R2_6_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6844\,
            in1 => \N__6838\,
            in2 => \_gnd_net_\,
            in3 => \N__10681\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIF8TM3_9_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11898\,
            in2 => \N__6829\,
            in3 => \N__10911\,
            lcout => \beamY_RNIF8TM3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_4_rep1_RNIQOGL_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110100101"
        )
    port map (
            in0 => \N__10452\,
            in1 => \N__10680\,
            in2 => \N__10552\,
            in3 => \N__10595\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVD444_9_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__11900\,
            in1 => \N__10912\,
            in2 => \N__7132\,
            in3 => \N__7995\,
            lcout => OPEN,
            ltout => \beamY_RNIVD444Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9G078_9_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7120\,
            in2 => \N__7114\,
            in3 => \N__7978\,
            lcout => OPEN,
            ltout => \font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUP21C_9_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010001"
        )
    port map (
            in0 => \N__7111\,
            in1 => \N__11786\,
            in2 => \N__7054\,
            in3 => \N__11899\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_10_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010111000"
        )
    port map (
            in0 => \N__7402\,
            in1 => \N__7171\,
            in2 => \N__7243\,
            in3 => \N__11437\,
            lcout => OPEN,
            ltout => \N_7_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_3_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__13075\,
            in1 => \N__8206\,
            in2 => \N__7045\,
            in3 => \N__7198\,
            lcout => \N_338_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4H2_6_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10458\,
            lcout => un8_beamy_3,
            ltout => \un8_beamy_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISKOB_4_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__10693\,
            in1 => \_gnd_net_\,
            in2 => \N__7042\,
            in3 => \N__7871\,
            lcout => un8_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_26_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011101010101"
        )
    port map (
            in0 => \N__11088\,
            in1 => \N__7039\,
            in2 => \N__7033\,
            in3 => \N__7156\,
            lcout => OPEN,
            ltout => \font_un127_pixel_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_11_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101100"
        )
    port map (
            in0 => \N__7207\,
            in1 => \N__7162\,
            in2 => \N__7201\,
            in3 => \N__7234\,
            lcout => \N_336_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7872\,
            in1 => \N__7192\,
            in2 => \N__7186\,
            in3 => \N__11089\,
            lcout => \beamY_RNI9DLCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_23_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__13074\,
            in1 => \_gnd_net_\,
            in2 => \N__8205\,
            in3 => \_gnd_net_\,
            lcout => g1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_41_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8562\,
            in1 => \N__7222\,
            in2 => \_gnd_net_\,
            in3 => \N__7369\,
            lcout => OPEN,
            ltout => \N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_25_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10095\,
            in2 => \N__7165\,
            in3 => \N__8151\,
            lcout => \N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEQIGK2_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__13071\,
            in1 => \N__11434\,
            in2 => \_gnd_net_\,
            in3 => \N__8195\,
            lcout => font_un13_pixel_23,
            ltout => \font_un13_pixel_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_35_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__7633\,
            in1 => \N__7150\,
            in2 => \N__7144\,
            in3 => \N__8233\,
            lcout => font_un127_pixel_m_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_39_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7141\,
            in1 => \N__8561\,
            in2 => \_gnd_net_\,
            in3 => \N__7213\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_22_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11112\,
            in2 => \N__7135\,
            in3 => \N__7249\,
            lcout => \N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_24_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__13072\,
            in1 => \N__11435\,
            in2 => \_gnd_net_\,
            in3 => \N__8196\,
            lcout => \N_5_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_45_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001000"
        )
    port map (
            in0 => \N__9446\,
            in1 => \N__9285\,
            in2 => \N__9020\,
            in3 => \N__8788\,
            lcout => OPEN,
            ltout => \g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_28_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__10087\,
            in1 => \N__8517\,
            in2 => \N__7228\,
            in3 => \N__7339\,
            lcout => \N_326_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011101000000"
        )
    port map (
            in0 => \N__7811\,
            in1 => \N__13292\,
            in2 => \N__11131\,
            in3 => \N__10088\,
            lcout => un43lto1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_4_0_1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000000000"
        )
    port map (
            in0 => \N__8785\,
            in1 => \N__8942\,
            in2 => \N__9289\,
            in3 => \N__9443\,
            lcout => OPEN,
            ltout => \N_250_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVV787O2_2_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__8516\,
            in1 => \_gnd_net_\,
            in2 => \N__7225\,
            in3 => \N__7255\,
            lcout => \beamY_RNIVV787O2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_1_i_1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9283\,
            in1 => \N__8943\,
            in2 => \_gnd_net_\,
            in3 => \N__9444\,
            lcout => \N_266_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_87_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100000101000"
        )
    port map (
            in0 => \N__9445\,
            in1 => \N__9284\,
            in2 => \N__9019\,
            in3 => \N__8786\,
            lcout => OPEN,
            ltout => \N_242_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_61_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__8787\,
            in1 => \_gnd_net_\,
            in2 => \N__7216\,
            in3 => \N__10086\,
            lcout => \Pixel_1_RNOZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_69_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111000"
        )
    port map (
            in0 => \N__8727\,
            in1 => \N__7261\,
            in2 => \N__10134\,
            in3 => \N__7279\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_69_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_44_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__8527\,
            in1 => \_gnd_net_\,
            in2 => \N__7273\,
            in3 => \N__7270\,
            lcout => \Pixel_1_RNOZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_1_i_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__9431\,
            in1 => \N__8938\,
            in2 => \N__8775\,
            in3 => \N__9252\,
            lcout => \N_268_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_91_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100101111"
        )
    port map (
            in0 => \N__9247\,
            in1 => \N__8719\,
            in2 => \N__9017\,
            in3 => \N__9428\,
            lcout => OPEN,
            ltout => \g0_35_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_76_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000111000010"
        )
    port map (
            in0 => \N__9432\,
            in1 => \N__8526\,
            in2 => \N__7264\,
            in3 => \N__9253\,
            lcout => \N_314_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15___m1_e_0_1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__8936\,
            in1 => \_gnd_net_\,
            in2 => \N__9286\,
            in3 => \N__9429\,
            lcout => \un115_pixel_13_15___m1_e_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__m9_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010001000"
        )
    port map (
            in0 => \N__9430\,
            in1 => \N__8937\,
            in2 => \N__8774\,
            in3 => \N__9251\,
            lcout => \un115_pixel_13_15__i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__g0_9_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__9254\,
            in1 => \N__8726\,
            in2 => \N__9018\,
            in3 => \N__9433\,
            lcout => \N_219_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14085\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_cry_2_s_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8262\,
            in2 => \N__11353\,
            in3 => \N__7318\,
            lcout => if_generate_plus_mult1_un75_sum_cry_2_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8868\,
            in2 => \N__8305\,
            in3 => \N__7306\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un82_sum_axb_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9181\,
            in1 => \N__8263\,
            in2 => \N__8293\,
            in3 => \N__7297\,
            lcout => \un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_s_5_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8278\,
            in2 => \_gnd_net_\,
            in3 => \N__7294\,
            lcout => un7_pixel_1_axb1,
            ltout => \un7_pixel_1_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__un115_pixel_1_i_9_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001001001100"
        )
    port map (
            in0 => \N__8872\,
            in1 => \N__8735\,
            in2 => \N__7291\,
            in3 => \N__9426\,
            lcout => OPEN,
            ltout => \N_203_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_47_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__8571\,
            in1 => \_gnd_net_\,
            in2 => \N__7288\,
            in3 => \N__7285\,
            lcout => \Pixel_1_RNOZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_92_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010110001101"
        )
    port map (
            in0 => \N__9182\,
            in1 => \N__8734\,
            in2 => \N__8951\,
            in3 => \N__9425\,
            lcout => g0_18_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__g0_7_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000100000"
        )
    port map (
            in0 => \N__9406\,
            in1 => \N__8990\,
            in2 => \N__9264\,
            in3 => \N__8688\,
            lcout => \N_192_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_72_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101111111"
        )
    port map (
            in0 => \N__8689\,
            in1 => \N__9197\,
            in2 => \N__9040\,
            in3 => \N__9408\,
            lcout => \Pixel_1_RNOZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un115_pixel_13_15__g0_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000101000"
        )
    port map (
            in0 => \N__9409\,
            in1 => \N__8995\,
            in2 => \N__9265\,
            in3 => \N__8691\,
            lcout => \N_234_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_90_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011110100001"
        )
    port map (
            in0 => \N__8991\,
            in1 => \N__10146\,
            in2 => \N__9267\,
            in3 => \N__9407\,
            lcout => g0_40_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_65_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010110001000"
        )
    port map (
            in0 => \N__9410\,
            in1 => \N__8996\,
            in2 => \N__9266\,
            in3 => \N__8692\,
            lcout => \N_206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_84_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101101111"
        )
    port map (
            in0 => \N__8690\,
            in1 => \N__10147\,
            in2 => \N__9268\,
            in3 => \N__9411\,
            lcout => OPEN,
            ltout => \g0_6_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_57_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101001111111"
        )
    port map (
            in0 => \N__9204\,
            in1 => \N__10128\,
            in2 => \N__7360\,
            in3 => \N__8997\,
            lcout => OPEN,
            ltout => \g0_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_37_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101110"
        )
    port map (
            in0 => \N__10129\,
            in1 => \N__8568\,
            in2 => \N__7357\,
            in3 => \N__7354\,
            lcout => \N_302_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_71_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001110000"
        )
    port map (
            in0 => \N__8760\,
            in1 => \N__9260\,
            in2 => \N__9051\,
            in3 => \N__9422\,
            lcout => OPEN,
            ltout => \g1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_46_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101011011111"
        )
    port map (
            in0 => \N__9423\,
            in1 => \N__8569\,
            in2 => \N__7342\,
            in3 => \N__9010\,
            lcout => g1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_85_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__9011\,
            in1 => \N__10153\,
            in2 => \_gnd_net_\,
            in3 => \N__9424\,
            lcout => OPEN,
            ltout => \g0_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_58_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100110011"
        )
    port map (
            in0 => \N__9261\,
            in1 => \N__10133\,
            in2 => \N__7327\,
            in3 => \N__8761\,
            lcout => OPEN,
            ltout => \N_309_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_38_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__8570\,
            in1 => \_gnd_net_\,
            in2 => \N__7420\,
            in3 => \N__7417\,
            lcout => OPEN,
            ltout => \N_323_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_21_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11091\,
            in2 => \N__7411\,
            in3 => \N__7408\,
            lcout => \N_5_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8022\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13225\,
            ce => \N__13275\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10160\,
            in2 => \N__11128\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_RNIAL73_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7466\,
            in2 => \_gnd_net_\,
            in3 => \N__7390\,
            lcout => \un21_beamy_cry_1_c_RNIALZ0Z73\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_2_c_RNICO83_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7566\,
            in2 => \_gnd_net_\,
            in3 => \N__7387\,
            lcout => \un21_beamy_cry_2_c_RNICOZ0Z83\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_3_c_RNIER93_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7890\,
            in2 => \_gnd_net_\,
            in3 => \N__7384\,
            lcout => \un21_beamy_cry_3_c_RNIERZ0Z93\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_4_c_RNIGUA3_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10465\,
            in2 => \_gnd_net_\,
            in3 => \N__7381\,
            lcout => \un21_beamy_cry_4_c_RNIGUAZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_5_c_RNII1C3_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10558\,
            in2 => \_gnd_net_\,
            in3 => \N__7378\,
            lcout => \un21_beamy_cry_5_c_RNII1CZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_6_c_RNIK4D3_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11004\,
            in2 => \_gnd_net_\,
            in3 => \N__7624\,
            lcout => \un21_beamy_cry_6_c_RNIK4DZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_7_c_RNIM7E3_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10793\,
            in2 => \_gnd_net_\,
            in3 => \N__7612\,
            lcout => \un21_beamy_cry_7_c_RNIM7EZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_8_c_RNIOAF3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10880\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7609\,
            lcout => \un21_beamy_cry_8_c_RNIOAFZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5NLM2_3_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11915\,
            in1 => \N__11810\,
            in2 => \N__7429\,
            in3 => \N__12146\,
            lcout => un11_visibleylto9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__12080\,
            in1 => \N__14592\,
            in2 => \_gnd_net_\,
            in3 => \N__7482\,
            lcout => \beamY_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9660\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIALEQ_0_9_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__10879\,
            in1 => \N__7996\,
            in2 => \_gnd_net_\,
            in3 => \N__7974\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_0_3_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000100010"
        )
    port map (
            in0 => \N__10464\,
            in1 => \N__7585\,
            in2 => \N__7497\,
            in3 => \N__7879\,
            lcout => un11_visibleylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9595\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIEP79_7_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10463\,
            in1 => \N__7711\,
            in2 => \_gnd_net_\,
            in3 => \N__7694\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_6_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7917\,
            lcout => \beamY_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13219\,
            ce => \N__13273\,
            sr => \_gnd_net_\
        );

    \beamY_fast_7_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7953\,
            in2 => \_gnd_net_\,
            in3 => \N__7816\,
            lcout => \beamY_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13219\,
            ce => \N__13273\,
            sr => \_gnd_net_\
        );

    \beamY_fast_5_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7731\,
            lcout => \beamY_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13219\,
            ce => \N__13273\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIRPUB_7_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7710\,
            in1 => \N__7690\,
            in2 => \_gnd_net_\,
            in3 => \N__7661\,
            lcout => un5_visibley_c6_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFC4H3_9_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10915\,
            in1 => \N__7645\,
            in2 => \_gnd_net_\,
            in3 => \N__10366\,
            lcout => un11_visibley,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI198K_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110011"
        )
    port map (
            in0 => \N__10712\,
            in1 => \N__10811\,
            in2 => \N__10597\,
            in3 => \N__10613\,
            lcout => OPEN,
            ltout => \beamY_fast_RNI198KZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQNF11_8_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__10812\,
            in1 => \_gnd_net_\,
            in2 => \N__7636\,
            in3 => \N__7973\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_54_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__10641\,
            in1 => \N__12691\,
            in2 => \N__11182\,
            in3 => \N__14422\,
            lcout => font_un127_pixel_m_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_2_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8026\,
            lcout => \beamY_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13217\,
            ce => \N__13271\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIG57D_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__10711\,
            in1 => \N__10612\,
            in2 => \N__8011\,
            in3 => \N__7853\,
            lcout => \beamY_fast_RNIG57DZ0Z_8\,
            ltout => \beamY_fast_RNIG57DZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIBV5P_8_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7981\,
            in3 => \N__7972\,
            lcout => un5_visibley_c7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_7_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7954\,
            in2 => \_gnd_net_\,
            in3 => \N__7786\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \beamY_fast_3_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7936\,
            lcout => \beamY_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7918\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7784\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \beamY_4_rep1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \beamY_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7735\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13216\,
            ce => \N__13270\,
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__13179\,
            in1 => \N__11377\,
            in2 => \N__8128\,
            in3 => \N__8056\,
            lcout => OPEN,
            ltout => \font_un127_pixel_m_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__8090\,
            in1 => \N__12787\,
            in2 => \N__8119\,
            in3 => \N__10621\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13213\,
            ce => 'H',
            sr => \N__11337\
        );

    \Pixel_1_RNO_16_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000000"
        )
    port map (
            in0 => \N__8224\,
            in1 => \N__12690\,
            in2 => \N__14421\,
            in3 => \N__8077\,
            lcout => OPEN,
            ltout => \g0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_5_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011100000"
        )
    port map (
            in0 => \N__8563\,
            in1 => \N__10144\,
            in2 => \N__8071\,
            in3 => \N__8068\,
            lcout => g0_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13066\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JF_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8215\,
            in2 => \N__8043\,
            in3 => \N__8050\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_82_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10750\,
            in2 => \N__11200\,
            in3 => \N__8047\,
            lcout => \Pixel_1_RNOZ0Z_82\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11248\,
            in2 => \N__8044\,
            in3 => \N__11195\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJ2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11218\,
            in2 => \_gnd_net_\,
            in3 => \N__8029\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2\,
            ltout => \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_31_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__13069\,
            in1 => \_gnd_net_\,
            in2 => \N__8245\,
            in3 => \_gnd_net_\,
            lcout => g1_0_0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_83_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__13180\,
            in1 => \N__13067\,
            in2 => \_gnd_net_\,
            in3 => \N__11433\,
            lcout => OPEN,
            ltout => \font_un127_pixel_m_4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_55_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110000010"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__8242\,
            in2 => \N__8236\,
            in3 => \N__8197\,
            lcout => font_un127_pixel_m_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_56_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__8950\,
            in1 => \N__9287\,
            in2 => \_gnd_net_\,
            in3 => \N__9492\,
            lcout => OPEN,
            ltout => \un7_pixel_1_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_36_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111110111"
        )
    port map (
            in0 => \N__11599\,
            in1 => \N__8796\,
            in2 => \N__8227\,
            in3 => \N__11524\,
            lcout => font_un127_pixel_m_7_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14086\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHMV0K2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13073\,
            in2 => \_gnd_net_\,
            in3 => \N__8198\,
            lcout => font_un13_pixel_0_1_0_0_22,
            ltout => \font_un13_pixel_0_1_0_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_32_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111011"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__8167\,
            in2 => \N__8155\,
            in3 => \N__8374\,
            lcout => g1_4_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_29_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001111111"
        )
    port map (
            in0 => \N__10096\,
            in1 => \N__8152\,
            in2 => \N__11129\,
            in3 => \N__8137\,
            lcout => OPEN,
            ltout => \N_1482_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_13_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11119\,
            in2 => \N__8308\,
            in3 => \N__8416\,
            lcout => \N_1870_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13970\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8331\,
            in2 => \N__11284\,
            in3 => \N__8296\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9427\,
            in2 => \N__8323\,
            in3 => \N__8281\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8867\,
            in1 => \N__8332\,
            in2 => \N__9526\,
            in3 => \N__8272\,
            lcout => \un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9511\,
            in2 => \_gnd_net_\,
            in3 => \N__8269\,
            lcout => un7_pixel_1_axb2,
            ltout => \un7_pixel_1_axb2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_pixel_1_axb2_sbtinv_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8266\,
            in3 => \_gnd_net_\,
            lcout => un7_pixel_1_axb2_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_27_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__8574\,
            in1 => \N__8254\,
            in2 => \N__10161\,
            in3 => \N__8362\,
            lcout => OPEN,
            ltout => \N_305_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_12_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11124\,
            in2 => \N__8248\,
            in3 => \N__8395\,
            lcout => \N_1869_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_77_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011111111110"
        )
    port map (
            in0 => \N__9016\,
            in1 => \N__8389\,
            in2 => \N__8578\,
            in3 => \N__8790\,
            lcout => OPEN,
            ltout => \N_321_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_50_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10151\,
            in1 => \_gnd_net_\,
            in2 => \N__8383\,
            in3 => \N__8380\,
            lcout => \N_328_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_93_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__9367\,
            in1 => \N__9255\,
            in2 => \N__9052\,
            in3 => \N__8789\,
            lcout => OPEN,
            ltout => \g1_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_80_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__10150\,
            in1 => \_gnd_net_\,
            in2 => \N__8365\,
            in3 => \N__8358\,
            lcout => OPEN,
            ltout => \un117_pixel_6_1_0_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_52_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000111110"
        )
    port map (
            in0 => \N__8567\,
            in1 => \N__10152\,
            in2 => \N__8341\,
            in3 => \N__8338\,
            lcout => \N_324_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_pixel_1_axb3_sbtinv_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9366\,
            lcout => un7_pixel_1_axb3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13868\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_cry_2_s_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8403\,
            in2 => \N__9073\,
            in3 => \N__8311\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11517\,
            in2 => \N__11611\,
            in3 => \N__9514\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_axb_5_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__8404\,
            in2 => \N__11569\,
            in3 => \N__9502\,
            lcout => \un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_s_5_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11542\,
            in2 => \_gnd_net_\,
            in3 => \N__9499\,
            lcout => un7_pixel_1_axb3,
            ltout => \un7_pixel_1_axb3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_89_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111000000"
        )
    port map (
            in0 => \N__10145\,
            in1 => \N__8989\,
            in2 => \N__9292\,
            in3 => \N__9183\,
            lcout => un117_pixel_2_6_i3_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_N_532_i_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13763\,
            lcout => \N_532_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_73_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010010011"
        )
    port map (
            in0 => \N__9064\,
            in1 => \N__9012\,
            in2 => \N__8797\,
            in3 => \N__10148\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_48_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8572\,
            in2 => \N__8587\,
            in3 => \N__8584\,
            lcout => OPEN,
            ltout => \Pixel_1_RNOZ0Z_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_30_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8573\,
            in1 => \N__10149\,
            in2 => \N__8425\,
            in3 => \N__8422\,
            lcout => \d_N_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_pixel_0_axb3_sbtinv_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11515\,
            lcout => un7_pixel_0_axb3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9740\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11687\,
            in2 => \N__9604\,
            in3 => \N__9622\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11737\,
            in2 => \N__11692\,
            in3 => \N__9619\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTA2_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11691\,
            in2 => \N__11728\,
            in3 => \N__9616\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI809T4_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9811\,
            in1 => \N__9757\,
            in2 => \N__11716\,
            in3 => \N__9613\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11704\,
            in2 => \_gnd_net_\,
            in3 => \N__9610\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2\,
            ltout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_0_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9607\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11812\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9586\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQO93_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9812\,
            in2 => \N__9673\,
            in3 => \N__9829\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFP3_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9826\,
            in2 => \N__9817\,
            in3 => \N__9820\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGC94_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9816\,
            in2 => \N__9796\,
            in3 => \N__9787\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV5NMA_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9882\,
            in1 => \N__9784\,
            in2 => \N__9778\,
            in3 => \N__9769\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9766\,
            in2 => \_gnd_net_\,
            in3 => \N__9760\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11685\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9741\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLK5_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9877\,
            in2 => \N__9937\,
            in3 => \N__9928\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAP8_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9925\,
            in2 => \N__9883\,
            in3 => \N__9919\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIB9299_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9881\,
            in2 => \N__9916\,
            in3 => \N__9907\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIVO5IK_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10247\,
            in1 => \N__9859\,
            in2 => \N__9904\,
            in3 => \N__9895\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PA_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9892\,
            in2 => \_gnd_net_\,
            in3 => \N__9886\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9876\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12072\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5B_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9853\,
            in2 => \N__10248\,
            in3 => \N__9844\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMG_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10243\,
            in2 => \N__9841\,
            in3 => \N__9832\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_18_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10270\,
            in2 => \N__10249\,
            in3 => \N__10264\,
            lcout => \Pixel_1_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10222\,
            in2 => \N__10261\,
            in3 => \N__10239\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQK_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10210\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_6_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__10207\,
            in1 => \N__12037\,
            in2 => \N__10201\,
            in3 => \N__10183\,
            lcout => \un1_beamY_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIALEQ_1_9_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10194\,
            lcout => \beamY_RNIALEQ_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_20_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010001000"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__10182\,
            in2 => \N__12084\,
            in3 => \N__10170\,
            lcout => OPEN,
            ltout => \un43lto4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_9_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__10171\,
            in1 => \N__10162\,
            in2 => \N__9949\,
            in3 => \N__12079\,
            lcout => OPEN,
            ltout => \un43lt10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011110"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__10372\,
            in2 => \N__9946\,
            in3 => \N__9943\,
            lcout => un44,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_8_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100011000100"
        )
    port map (
            in0 => \N__13882\,
            in1 => \N__10312\,
            in2 => \N__13990\,
            in3 => \N__10318\,
            lcout => un42lt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIALEQ_9_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10924\,
            in2 => \_gnd_net_\,
            in3 => \N__10361\,
            lcout => \beamY_RNIALEQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13880\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10329\,
            in2 => \N__11368\,
            in3 => \N__10336\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_19_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12031\,
            in2 => \N__11995\,
            in3 => \N__10333\,
            lcout => \Pixel_1_RNOZ0Z_19\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10330\,
            in2 => \N__12019\,
            in3 => \N__11990\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5AS_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12007\,
            in2 => \_gnd_net_\,
            in3 => \N__10321\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_7_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111110110000"
        )
    port map (
            in0 => \N__13881\,
            in1 => \N__10311\,
            in2 => \N__10300\,
            in3 => \N__10297\,
            lcout => un1_visiblex_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIHT1O_3_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__10555\,
            in1 => \N__10451\,
            in2 => \N__10567\,
            in3 => \N__10714\,
            lcout => un5_visibley_ac0_7,
            ltout => \un5_visibley_ac0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4S2S1_7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__10985\,
            in1 => \N__10556\,
            in2 => \N__10738\,
            in3 => \N__12133\,
            lcout => font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_4_rep1_RNICDQE_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__10439\,
            in1 => \N__10527\,
            in2 => \N__10991\,
            in3 => \N__10593\,
            lcout => OPEN,
            ltout => \beamY_4_rep1_RNICDQEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIB5JQ_7_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10378\,
            in2 => \N__10717\,
            in3 => \N__10665\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIBVU7_2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10713\,
            in2 => \_gnd_net_\,
            in3 => \N__10614\,
            lcout => un5_visibley_c2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__12783\,
            in1 => \N__12762\,
            in2 => \N__10645\,
            in3 => \N__10630\,
            lcout => \Pixel_1_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIK8HH_2_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__10615\,
            in1 => \N__10528\,
            in2 => \N__10462\,
            in3 => \N__10594\,
            lcout => \beamY_fast_RNIK8HHZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKOP3_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__10526\,
            in1 => \N__10969\,
            in2 => \_gnd_net_\,
            in3 => \N__10435\,
            lcout => \beamY_RNIKOP3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13982\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKB_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11014\,
            in2 => \N__12276\,
            in3 => \N__11029\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONH_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12295\,
            in2 => \N__12334\,
            in3 => \N__11026\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI0MA3B1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11259\,
            in1 => \N__12322\,
            in2 => \N__12277\,
            in3 => \N__11023\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12313\,
            in2 => \_gnd_net_\,
            in3 => \N__11020\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0\,
            ltout => \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11017\,
            in3 => \_gnd_net_\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13870\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMJIF_8_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__10925\,
            in2 => \N__10831\,
            in3 => \N__10819\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGM_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12403\,
            in2 => \N__11232\,
            in3 => \N__10741\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPC321_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11269\,
            in2 => \N__11263\,
            in3 => \N__11242\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJFAHJ2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11199\,
            in1 => \N__11239\,
            in2 => \N__11233\,
            in3 => \N__11212\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQAB1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11209\,
            in2 => \_gnd_net_\,
            in3 => \N__11203\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_81_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__13642\,
            in1 => \N__13869\,
            in2 => \N__11167\,
            in3 => \N__13765\,
            lcout => un14_visibleylt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_94_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13070\,
            in1 => \N__14091\,
            in2 => \_gnd_net_\,
            in3 => \N__13983\,
            lcout => un14_visibleylt4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__14123\,
            in1 => \N__13120\,
            in2 => \N__14038\,
            in3 => \N__13178\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_10_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13927\,
            in1 => \N__14128\,
            in2 => \N__13390\,
            in3 => \N__13118\,
            lcout => OPEN,
            ltout => \un3_beamx_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13693\,
            in1 => \N__14037\,
            in2 => \N__11158\,
            in3 => \N__13168\,
            lcout => un3_beamx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_33_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010011"
        )
    port map (
            in0 => \N__11155\,
            in1 => \N__11143\,
            in2 => \N__11130\,
            in3 => \N__11385\,
            lcout => OPEN,
            ltout => \g3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_14_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__11443\,
            in1 => \N__11436\,
            in2 => \N__11410\,
            in3 => \N__11407\,
            lcout => OPEN,
            ltout => \font_un127_pixel_6_ns_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__11401\,
            in1 => \N__11395\,
            in2 => \N__11389\,
            in3 => \N__11386\,
            lcout => \N_520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13762\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un68_sum_i_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13971\,
            lcout => \un4_pixel_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11338\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_i_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13856\,
            lcout => \un4_pixel_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13641\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_m_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__11464\,
            in1 => \N__14406\,
            in2 => \N__12523\,
            in3 => \N__11272\,
            lcout => if_generate_plus_mult1_un47_sum_m_2,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12565\,
            in2 => \N__12544\,
            in3 => \N__11473\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum1_3,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14407\,
            in2 => \N__12574\,
            in3 => \N__11470\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum1_4,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__14408\,
            in1 => \N__13521\,
            in2 => \N__14707\,
            in3 => \N__11467\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13634\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12550\,
            in2 => \N__12559\,
            in3 => \N__11458\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum0_2,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12724\,
            in2 => \N__12718\,
            in3 => \N__11455\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum0_3,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12709\,
            in2 => \N__12619\,
            in3 => \N__11452\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum0_4,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14409\,
            in2 => \_gnd_net_\,
            in3 => \N__11449\,
            lcout => un4_pixel_if_generate_plus_mult1_un47_sum0_5,
            ltout => \un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_m_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__11628\,
            in1 => \_gnd_net_\,
            in2 => \N__11446\,
            in3 => \N__14413\,
            lcout => un7_pixel_0_axb4,
            ltout => \un7_pixel_0_axb4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un54_sum_axb_5_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110100101"
        )
    port map (
            in0 => \N__11644\,
            in1 => \N__11638\,
            in2 => \N__11632\,
            in3 => \N__14411\,
            lcout => \un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_un7_pixel_0_axb4_i_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__14410\,
            in1 => \_gnd_net_\,
            in2 => \N__11629\,
            in3 => \N__11617\,
            lcout => un7_pixel_0_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13760\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => un4_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12535\,
            in2 => \N__11556\,
            in3 => \N__11602\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => un4_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11592\,
            in2 => \N__11581\,
            in3 => \N__11560\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => un4_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un61_sum_axb_5_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11516\,
            in1 => \N__11479\,
            in2 => \N__11557\,
            in3 => \N__11536\,
            lcout => \un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => un4_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => un4_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un54_sum_s_5_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11533\,
            in2 => \_gnd_net_\,
            in3 => \N__11527\,
            lcout => un7_pixel_0_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_m_3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11494\,
            in1 => \N__11485\,
            in2 => \_gnd_net_\,
            in3 => \N__14412\,
            lcout => if_generate_plus_mult1_un47_sum_m_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11811\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11947\,
            in2 => \N__11851\,
            in3 => \N__11731\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689H1_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11665\,
            in2 => \N__11953\,
            in3 => \N__11719\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11951\,
            in2 => \N__11656\,
            in3 => \N__11707\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI69052_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11686\,
            in1 => \N__11932\,
            in2 => \N__11977\,
            in3 => \N__11698\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11965\,
            in1 => \N__11952\,
            in2 => \N__12172\,
            in3 => \N__11695\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11916\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHT921_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12091\,
            in2 => \N__14606\,
            in3 => \N__11659\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11836\,
            in2 => \N__14556\,
            in3 => \N__11647\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11821\,
            in2 => \N__14607\,
            in3 => \N__11968\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12164\,
            in2 => \_gnd_net_\,
            in3 => \N__11959\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12181\,
            in2 => \_gnd_net_\,
            in3 => \N__11956\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11935\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11917\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12147\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11842\,
            in2 => \N__14608\,
            in3 => \N__11830\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11827\,
            in2 => \N__14609\,
            in3 => \N__11815\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12184\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12175\,
            in3 => \N__12168\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQNF11_0_8_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_RNIQNF11_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_17_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12085\,
            in2 => \_gnd_net_\,
            in3 => \N__12048\,
            lcout => \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13764\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VG6_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12247\,
            in2 => \N__12256\,
            in3 => \N__12022\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6N9_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12241\,
            in2 => \N__12205\,
            in3 => \N__12010\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIE7K6S_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11994\,
            in1 => \N__12262\,
            in2 => \N__12232\,
            in3 => \N__12001\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07C_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12217\,
            in2 => \_gnd_net_\,
            in3 => \N__11998\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPA_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__12231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12200\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13637\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12199\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13636\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMS983_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12342\,
            in2 => \N__12472\,
            in3 => \N__12235\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAO4_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12607\,
            in2 => \N__12460\,
            in3 => \N__12220\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI9MMPB_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12204\,
            in1 => \N__12343\,
            in2 => \N__12442\,
            in3 => \N__12211\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12208\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI8P51_4_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__13925\,
            in1 => \N__13686\,
            in2 => \N__12844\,
            in3 => \N__13808\,
            lcout => un13_beamylt7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12763\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12606\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13879\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRF156_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12301\,
            in2 => \N__12903\,
            in3 => \N__12325\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RA99_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12919\,
            in2 => \N__12973\,
            in3 => \N__12316\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIOK72M_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12294\,
            in1 => \N__12952\,
            in2 => \N__12904\,
            in3 => \N__12307\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12937\,
            in2 => \_gnd_net_\,
            in3 => \N__12304\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13761\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12293\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13635\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3D1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13231\,
            in2 => \N__12486\,
            in3 => \N__12415\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UD62_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12502\,
            in2 => \N__12394\,
            in3 => \N__12412\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIF5PB5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12889\,
            in1 => \N__12382\,
            in2 => \N__12487\,
            in3 => \N__12409\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12514\,
            in2 => \_gnd_net_\,
            in3 => \N__12406\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13975\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNISG94_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13499\,
            in2 => \_gnd_net_\,
            in3 => \N__14699\,
            lcout => \N_32\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DR_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14449\,
            in2 => \N__12583\,
            in3 => \N__12385\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3U41_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13314\,
            in2 => \N__14650\,
            in3 => \N__12376\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIOPOL2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12501\,
            in1 => \N__14493\,
            in2 => \N__13303\,
            in3 => \N__12508\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14467\,
            in1 => \N__13315\,
            in2 => \N__14414\,
            in3 => \N__12505\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251\,
            ltout => \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12490\,
            in3 => \_gnd_net_\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13500\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNISG94_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13501\,
            in2 => \_gnd_net_\,
            in3 => \N__14694\,
            lcout => \N_20_i\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3I1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14262\,
            in2 => \N__14272\,
            in3 => \N__12445\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPH2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14179\,
            in2 => \N__14254\,
            in3 => \N__12430\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7SRM5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__14263\,
            in2 => \N__14224\,
            in3 => \N__12418\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14200\,
            in2 => \_gnd_net_\,
            in3 => \N__12610\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14695\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__14361\,
            in1 => \_gnd_net_\,
            in2 => \N__12678\,
            in3 => \N__12738\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__12737\,
            in1 => \N__12662\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13502\,
            lcout => un5_visiblex_i_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__13511\,
            in1 => \N__12656\,
            in2 => \_gnd_net_\,
            in3 => \N__14355\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_m_1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13607\,
            in2 => \N__13632\,
            in3 => \N__14359\,
            lcout => if_generate_plus_mult1_un47_sum_m_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_3_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_visiblex_i_0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011111010"
        )
    port map (
            in0 => \N__12742\,
            in1 => \N__12657\,
            in2 => \N__12677\,
            in3 => \N__14358\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14356\,
            in1 => \N__12661\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => if_generate_plus_mult1_un47_sum_0_cry_3_ma,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNITTF6_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14362\,
            in2 => \_gnd_net_\,
            in3 => \N__12679\,
            lcout => \N_158_0_i\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMB_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14619\,
            in2 => \_gnd_net_\,
            in3 => \N__12703\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OB_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14631\,
            in2 => \N__14630\,
            in3 => \N__12700\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12697\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12694\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111100"
        )
    port map (
            in0 => \N__12686\,
            in1 => \N__14363\,
            in2 => \N__13522\,
            in3 => \N__14696\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14632\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12853\,
            in2 => \_gnd_net_\,
            in3 => \N__12847\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNII5M_9_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13556\,
            in1 => \N__13454\,
            in2 => \N__13423\,
            in3 => \N__13688\,
            lcout => OPEN,
            ltout => \un18_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_4_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__12840\,
            in1 => \N__13804\,
            in2 => \N__12823\,
            in3 => \N__13923\,
            lcout => OPEN,
            ltout => \un18_beamylt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNINAS01_10_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13388\,
            in1 => \N__12820\,
            in2 => \N__12811\,
            in3 => \N__12808\,
            lcout => OPEN,
            ltout => \un15_beamy_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIMPI21_7_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001010000"
        )
    port map (
            in0 => \N__13347\,
            in1 => \N__12796\,
            in2 => \N__12790\,
            in3 => \N__13557\,
            lcout => un15_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13455\,
            lcout => un1_beamx_2,
            ltout => \un1_beamx_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI34L6_10_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12748\,
            in1 => \N__13389\,
            in2 => \N__12766\,
            in3 => \N__13558\,
            lcout => un1_beamx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI6PL_3_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13924\,
            in1 => \N__13687\,
            in2 => \N__13810\,
            in3 => \N__14032\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13759\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AA63_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12859\,
            in2 => \N__12873\,
            in3 => \N__12964\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CH4_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12888\,
            in2 => \N__12961\,
            in3 => \N__12946\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIBH1VA_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12918\,
            in1 => \N__12943\,
            in2 => \N__12874\,
            in3 => \N__12931\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12928\,
            in2 => \_gnd_net_\,
            in3 => \N__12922\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5\,
            ltout => \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12907\,
            in3 => \_gnd_net_\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12887\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13633\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13164\,
            in2 => \N__13119\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14119\,
            in2 => \_gnd_net_\,
            in3 => \N__13000\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14025\,
            in2 => \_gnd_net_\,
            in3 => \N__12997\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13293\,
            in1 => \N__13916\,
            in2 => \_gnd_net_\,
            in3 => \N__12994\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13800\,
            in2 => \_gnd_net_\,
            in3 => \N__12991\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13679\,
            in2 => \_gnd_net_\,
            in3 => \N__12988\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13554\,
            in2 => \_gnd_net_\,
            in3 => \N__12985\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13450\,
            in2 => \_gnd_net_\,
            in3 => \N__12982\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__13223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13417\,
            in2 => \_gnd_net_\,
            in3 => \N__12979\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__13224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__13384\,
            in1 => \N__13291\,
            in2 => \_gnd_net_\,
            in3 => \N__12976\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13360\,
            in1 => \N__13546\,
            in2 => \N__13351\,
            in3 => \N__13799\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9TH9_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14448\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9\,
            ltout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38L_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__14494\,
            in1 => \_gnd_net_\,
            in2 => \N__13306\,
            in3 => \_gnd_net_\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13290\,
            in2 => \_gnd_net_\,
            in3 => \N__13165\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13510\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13113\,
            in2 => \_gnd_net_\,
            in3 => \N__13166\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13167\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13114\,
            in3 => \N__13003\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14127\,
            in3 => \N__14041\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14593\,
            in2 => \N__14036\,
            in3 => \N__13930\,
            lcout => un1_visiblex_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13926\,
            in3 => \N__13813\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13809\,
            in3 => \N__13696\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14594\,
            in2 => \N__13689\,
            in3 => \N__13561\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13555\,
            in2 => \_gnd_net_\,
            in3 => \N__13459\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14595\,
            in2 => \N__13456\,
            in3 => \N__13426\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13418\,
            in2 => \_gnd_net_\,
            in3 => \N__13393\,
            lcout => un1_visiblex_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14698\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14174\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14697\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UP11_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14136\,
            in2 => \N__14158\,
            in3 => \N__14239\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBB1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14148\,
            in2 => \N__14236\,
            in3 => \N__14212\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_c_RNICFTM2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14175\,
            in1 => \N__14137\,
            in2 => \N__14209\,
            in3 => \N__14191\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14188\,
            in1 => \N__14149\,
            in2 => \_gnd_net_\,
            in3 => \N__14182\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14370\,
            lcout => un1_visiblex_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14147\,
            lcout => un1_visiblex_if_generate_plus_mult1_un40_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14700\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LB_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14281\,
            in3 => \N__14635\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MB_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14623\,
            in2 => \N__14431\,
            in3 => \N__14470\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14376\,
            in2 => \_gnd_net_\,
            in3 => \N__14455\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14452\,
            lcout => \font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14375\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_2_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14374\,
            lcout => font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
