-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 19:42:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un18_beamylto9_2_cascade_\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal un20_beamy_cry_1 : std_logic;
signal un20_beamy_cry_2 : std_logic;
signal un20_beamy_cry_3 : std_logic;
signal un20_beamy_cry_4 : std_logic;
signal un20_beamy_cry_5 : std_logic;
signal un20_beamy_cry_6 : std_logic;
signal un20_beamy_cry_7 : std_logic;
signal un20_beamy_cry_8 : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \un5_beamx_4_cascade_\ : std_logic;
signal \beamY_RNI9DLCZ0Z_5_cascade_\ : std_logic;
signal un5_beamx_3 : std_logic;
signal un5_beamx_2 : std_logic;
signal \un5_beamx_2_cascade_\ : std_logic;
signal \un8_beamylto9_1_cascade_\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal \un4_beamylt8_0_cascade_\ : std_logic;
signal un3_beamx_5 : std_logic;
signal \un3_beamx_7_cascade_\ : std_logic;
signal \un1_beamxlt10_0_cascade_\ : std_logic;
signal \HSync_c\ : std_logic;
signal un18_beamylt10_0 : std_logic;
signal un8_beamy : std_logic;
signal un4_beamy_0 : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un1_beamx_2 : std_logic;
signal un13_beamylt7 : std_logic;
signal \un15_beamy_2_cascade_\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal un5_visiblex_1_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un5_visiblex_1_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un5_visiblex_1_cry_2 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un5_visiblex_1_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un5_visiblex_1_cry_4 : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un5_visiblex_1_cry_5 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un5_visiblex_1_cry_6 : std_logic;
signal un5_visiblex_1_cry_7 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un5_visiblex_1_cry_8 : std_logic;
signal \un5_visiblex_1_n_23_cascade_\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \beamY_fast_RNIGR79Z0Z_7_cascade_\ : std_logic;
signal \beamY_RNIALEQ_0Z0Z_9\ : std_logic;
signal \un20_beamy_cry_2_c_RNIBADZ0Z4\ : std_logic;
signal \un20_beamy_cry_3_c_RNIDDEZ0Z4\ : std_logic;
signal \un20_beamy_cry_6_c_RNIJMHZ0Z4\ : std_logic;
signal \beamY_RNI9DLCZ0Z_5\ : std_logic;
signal \un20_beamy_cry_4_c_RNIFGFZ0Z4\ : std_logic;
signal un13_visiblex_2_0 : std_logic;
signal un12_visiblexlt9_0 : std_logic;
signal un13_visiblex_0 : std_logic;
signal font_un7_pixellt9_0 : std_logic;
signal \font_un14_pixellt9_0_cascade_\ : std_logic;
signal un13_visiblex_5 : std_logic;
signal \Pixel_0_sqmuxa_2\ : std_logic;
signal \un13_visiblex_5_cascade_\ : std_logic;
signal un5_visiblex_1_n_31 : std_logic;
signal un5_visiblex_1_n_30 : std_logic;
signal \N_159\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_\ : std_logic;
signal un5_visiblex_1_n_i_24 : std_logic;
signal un5_visiblex_1_n_24 : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal un5_visiblex_1_n_23 : std_logic;
signal \un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\ : std_logic;
signal \un5_visibley_c3_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\ : std_logic;
signal \beamY_fastZ0Z_7\ : std_logic;
signal \beamY_fastZ0Z_5\ : std_logic;
signal un5_visibley_c6_0_0_0 : std_logic;
signal \un5_visibley_c6_0_0_0_cascade_\ : std_logic;
signal un5_visibley_c3 : std_logic;
signal \beamY_RNIBV5PZ0Z_8\ : std_logic;
signal un13_visiblex_2 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cascade_\ : std_logic;
signal \beamY_fastZ0Z_3\ : std_logic;
signal \beamY_fastZ0Z_4\ : std_logic;
signal \un5_visibley_ac0_11_0_1_cascade_\ : std_logic;
signal \beamY_fast_RNIGR79Z0Z_7\ : std_logic;
signal \beamY_RNIALEQZ0Z_9\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cascade_\ : std_logic;
signal \font_un11_pixellto9_7_0_cascade_\ : std_logic;
signal \un8_beamx_cry_1_c_RNITP5AZ0\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \font_un26_pixel_0_cascade_\ : std_logic;
signal un5_visibley_ac0_11_0_1 : std_logic;
signal un5_visibley_c7 : std_logic;
signal \Pixel_0_sqmuxa_4\ : std_logic;
signal font_un11_pixel_0_7 : std_logic;
signal \un5_visibley_c7_cascade_\ : std_logic;
signal \Pixel_0_sqmuxa_7\ : std_logic;
signal \Pixel_0_sqmuxa_6\ : std_logic;
signal un15_beamy : std_logic;
signal \Pixel_0_sqmuxa_7_cascade_\ : std_logic;
signal un13_visiblex_4 : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un1_beamylto9_1 : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \un1_beamylto9_2_cascade_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \VSync_c\ : std_logic;
signal un5_visiblex_1_n_26 : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \beamX_RNIBKAZ0Z_1\ : std_logic;
signal un5_visiblex_1_n_25 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\ : std_logic;
signal \beamY_fastZ0Z_6\ : std_logic;
signal \un20_beamy_cry_5_c_RNIHJGZ0Z4\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \un20_beamy_cry_1_c_RNI97CZ0Z4\ : std_logic;
signal \beamY_fastZ0Z_2\ : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\ : std_logic;
signal un1_visiblex_24 : std_logic;
signal \un19lto10_1_1_cascade_\ : std_logic;
signal un5_visiblex_1_n_28 : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \Pixel_1_RNOZ0Z_13\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \Pixel_1_RNOZ0Z_6\ : std_logic;
signal un5_visiblex_1_n_27 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \G_6_i_a4_0_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \Pixel_1_RNOZ0Z_10\ : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \N_11\ : std_logic;
signal un19_0_1 : std_logic;
signal \d_N_3_mux\ : std_logic;
signal \un20_0_1_cascade_\ : std_logic;
signal \Pixel_5_N_3_mux\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    Pixel <= \Pixel_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__2634\,
            RESETB => \N__5457\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5956\,
            DIN => \N__5955\,
            DOUT => \N__5954\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5956\,
            PADOUT => \N__5955\,
            PADIN => \N__5954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5625\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5947\,
            DIN => \N__5946\,
            DOUT => \N__5945\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5947\,
            PADOUT => \N__5946\,
            PADIN => \N__5945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5938\,
            DIN => \N__5937\,
            DOUT => \N__5936\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5938\,
            PADOUT => \N__5937\,
            PADIN => \N__5936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5929\,
            DIN => \N__5928\,
            DOUT => \N__5927\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5929\,
            PADOUT => \N__5928\,
            PADIN => \N__5927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5920\,
            DIN => \N__5919\,
            DOUT => \N__5918\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5920\,
            PADOUT => \N__5919\,
            PADIN => \N__5918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5911\,
            DIN => \N__5910\,
            DOUT => \N__5909\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5911\,
            PADOUT => \N__5910\,
            PADIN => \N__5909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2781\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5902\,
            DIN => \N__5901\,
            DOUT => \N__5900\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5902\,
            PADOUT => \N__5901\,
            PADIN => \N__5900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1314\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5880\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__5877\,
            I => \N__5872\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__5876\,
            I => \N__5868\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5864\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5855\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5855\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5855\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5855\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5864\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5855\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5844\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5838\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5835\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5829\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5829\,
            I => \G_6_i_a4_0_0\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__5826\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__5820\,
            I => \N__5815\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5812\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5809\
        );

    \I__1290\ : Span4Mux_s0_h
    port map (
            O => \N__5815\,
            I => \N__5804\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5812\,
            I => \N__5804\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5809\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__5804\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5796\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5789\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5786\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5789\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5786\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5777\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5774\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5777\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5774\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__5769\,
            I => \N__5764\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5761\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5758\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5755\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5752\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5758\,
            I => \beamY_i_2\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5755\,
            I => \beamY_i_2\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__5752\,
            I => \beamY_i_2\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5742\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5735\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5732\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5735\,
            I => \N__5727\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5732\,
            I => \N__5723\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5720\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__5730\,
            I => \N__5717\
        );

    \I__1260\ : Span4Mux_s1_h
    port map (
            O => \N__5727\,
            I => \N__5714\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5710\
        );

    \I__1258\ : Span4Mux_s2_h
    port map (
            O => \N__5723\,
            I => \N__5705\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5720\,
            I => \N__5705\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5700\
        );

    \I__1255\ : Span4Mux_h
    port map (
            O => \N__5714\,
            I => \N__5697\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5694\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5691\
        );

    \I__1252\ : Span4Mux_h
    port map (
            O => \N__5705\,
            I => \N__5688\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5683\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5683\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5700\,
            I => \beamYZ0Z_1\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__5697\,
            I => \beamYZ0Z_1\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5694\,
            I => \beamYZ0Z_1\
        );

    \I__1246\ : Odrv12
    port map (
            O => \N__5691\,
            I => \beamYZ0Z_1\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__5688\,
            I => \beamYZ0Z_1\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5683\,
            I => \beamYZ0Z_1\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5667\,
            I => \Pixel_1_RNOZ0Z_10\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__5664\,
            I => \N_8_cascade_\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5658\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5658\,
            I => \N_11\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5652\,
            I => un19_0_1
        );

    \I__1236\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5646\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__1234\ : Span4Mux_s1_h
    port map (
            O => \N__5643\,
            I => \N__5640\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__5640\,
            I => \d_N_3_mux\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__5637\,
            I => \un20_0_1_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__5628\,
            I => \Pixel_5_N_3_mux\
        );

    \I__1228\ : IoInMux
    port map (
            O => \N__5625\,
            I => \N__5621\
        );

    \I__1227\ : IoInMux
    port map (
            O => \N__5624\,
            I => \N__5618\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5615\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5612\
        );

    \I__1224\ : Span12Mux_s2_v
    port map (
            O => \N__5615\,
            I => \N__5609\
        );

    \I__1223\ : Span4Mux_s3_v
    port map (
            O => \N__5612\,
            I => \N__5606\
        );

    \I__1222\ : Odrv12
    port map (
            O => \N__5609\,
            I => \Pixel_c\
        );

    \I__1221\ : Odrv4
    port map (
            O => \N__5606\,
            I => \Pixel_c\
        );

    \I__1220\ : ClkMux
    port map (
            O => \N__5601\,
            I => \N__5562\
        );

    \I__1219\ : ClkMux
    port map (
            O => \N__5600\,
            I => \N__5562\
        );

    \I__1218\ : ClkMux
    port map (
            O => \N__5599\,
            I => \N__5562\
        );

    \I__1217\ : ClkMux
    port map (
            O => \N__5598\,
            I => \N__5562\
        );

    \I__1216\ : ClkMux
    port map (
            O => \N__5597\,
            I => \N__5562\
        );

    \I__1215\ : ClkMux
    port map (
            O => \N__5596\,
            I => \N__5562\
        );

    \I__1214\ : ClkMux
    port map (
            O => \N__5595\,
            I => \N__5562\
        );

    \I__1213\ : ClkMux
    port map (
            O => \N__5594\,
            I => \N__5562\
        );

    \I__1212\ : ClkMux
    port map (
            O => \N__5593\,
            I => \N__5562\
        );

    \I__1211\ : ClkMux
    port map (
            O => \N__5592\,
            I => \N__5562\
        );

    \I__1210\ : ClkMux
    port map (
            O => \N__5591\,
            I => \N__5562\
        );

    \I__1209\ : ClkMux
    port map (
            O => \N__5590\,
            I => \N__5562\
        );

    \I__1208\ : ClkMux
    port map (
            O => \N__5589\,
            I => \N__5562\
        );

    \I__1207\ : GlobalMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1206\ : gio2CtrlBuf
    port map (
            O => \N__5559\,
            I => \PixelClock_g\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__5547\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5534\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5534\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5531\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5528\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5531\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__5528\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5517\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5517\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5517\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__1191\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5508\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__5508\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__1188\ : InMux
    port map (
            O => \N__5505\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__1187\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5499\,
            I => \Pixel_1_RNOZ0Z_6\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5493\,
            I => \N__5489\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5486\
        );

    \I__1182\ : Span4Mux_s2_h
    port map (
            O => \N__5489\,
            I => \N__5480\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5486\,
            I => \N__5480\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5477\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__5480\,
            I => \N__5474\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5477\,
            I => un5_visiblex_1_n_27
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__5474\,
            I => un5_visiblex_1_n_27
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5463\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__5460\,
            I => \N__5453\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__5459\,
            I => \N__5450\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__5458\,
            I => \N__5444\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__5457\,
            I => \N__5439\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5436\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5433\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5430\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__5449\,
            I => \N__5427\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__5448\,
            I => \N__5424\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__5447\,
            I => \N__5421\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5418\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5415\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \N__5412\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5408\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5436\,
            I => \N__5405\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5400\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5400\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5397\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5392\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5392\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5418\,
            I => \N__5389\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5386\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5381\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5381\
        );

    \I__1149\ : Span12Mux_s3_v
    port map (
            O => \N__5408\,
            I => \N__5378\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__5405\,
            I => \N__5373\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__5400\,
            I => \N__5373\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5368\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5368\
        );

    \I__1144\ : Sp12to4
    port map (
            O => \N__5389\,
            I => \N__5361\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5361\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5361\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__5378\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__5373\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__5368\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1138\ : Odrv12
    port map (
            O => \N__5361\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5340\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5340\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5337\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5330\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5330\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5330\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5327\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5323\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5340\,
            I => \N__5320\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5317\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5330\,
            I => \N__5312\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5312\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5309\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5323\,
            I => \N__5303\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__5320\,
            I => \N__5300\
        );

    \I__1122\ : Span4Mux_s3_h
    port map (
            O => \N__5317\,
            I => \N__5293\
        );

    \I__1121\ : Span4Mux_h
    port map (
            O => \N__5312\,
            I => \N__5293\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5309\,
            I => \N__5293\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5286\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5286\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5286\
        );

    \I__1116\ : Odrv12
    port map (
            O => \N__5303\,
            I => \beamYZ0Z_2\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__5300\,
            I => \beamYZ0Z_2\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__5293\,
            I => \beamYZ0Z_2\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5286\,
            I => \beamYZ0Z_2\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5277\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5268\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5265\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5259\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5256\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5247\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5244\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5238\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5235\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5227\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5224\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5221\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5217\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5214\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5211\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5208\
        );

    \I__1090\ : Span4Mux_s3_h
    port map (
            O => \N__5217\,
            I => \N__5205\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__5214\,
            I => \N__5200\
        );

    \I__1088\ : Span4Mux_s3_h
    port map (
            O => \N__5211\,
            I => \N__5200\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5208\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__5205\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__5200\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5187\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5179\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5176\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5173\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5179\,
            I => \N__5170\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5176\,
            I => \N__5167\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5164\
        );

    \I__1075\ : Span4Mux_s3_h
    port map (
            O => \N__5170\,
            I => \N__5161\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__5167\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__5164\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__5161\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__5154\,
            I => \N__5151\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5148\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5141\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \N__5137\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5133\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5126\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5126\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5126\
        );

    \I__1062\ : Span12Mux_s6_v
    port map (
            O => \N__5133\,
            I => \N__5123\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5126\,
            I => \N__5120\
        );

    \I__1060\ : Odrv12
    port map (
            O => \N__5123\,
            I => un1_visiblex_24
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__5120\,
            I => un1_visiblex_24
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__5115\,
            I => \un19lto10_1_1_cascade_\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__5112\,
            I => \N__5108\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5102\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5102\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5099\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5099\,
            I => \N__5093\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5096\,
            I => \N__5087\
        );

    \I__1050\ : Span4Mux_s1_h
    port map (
            O => \N__5093\,
            I => \N__5087\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5084\
        );

    \I__1048\ : Span4Mux_h
    port map (
            O => \N__5087\,
            I => \N__5081\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5078\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__5081\,
            I => un5_visiblex_1_n_28
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5078\,
            I => un5_visiblex_1_n_28
        );

    \I__1044\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5070\,
            I => \Pixel_1_RNOZ0Z_13\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5067\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1041\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__5058\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5049\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5049\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5046\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__1034\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5040\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5037\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5031\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5028\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__5022\,
            I => \N__5017\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5012\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5003\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5003\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5003\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5003\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5012\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5003\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4992\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4989\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4983\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4980\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__4977\,
            I => \N__4973\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4964\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4964\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4964\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4961\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4964\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4961\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4950\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4947\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4941\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5\
        );

    \I__999\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__4932\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\
        );

    \I__996\ : InMux
    port map (
            O => \N__4929\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__4926\,
            I => \N__4922\
        );

    \I__994\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4914\
        );

    \I__993\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4914\
        );

    \I__992\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4914\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4910\
        );

    \I__990\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4907\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__4910\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4907\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__986\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__4893\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81\
        );

    \I__983\ : InMux
    port map (
            O => \N__4890\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__982\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__4881\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__978\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__4869\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\
        );

    \I__975\ : InMux
    port map (
            O => \N__4866\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__974\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__4857\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\
        );

    \I__971\ : InMux
    port map (
            O => \N__4854\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__970\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4848\,
            I => \N__4842\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__4847\,
            I => \N__4839\
        );

    \I__967\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4834\
        );

    \I__966\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4834\
        );

    \I__965\ : Span4Mux_s1_v
    port map (
            O => \N__4842\,
            I => \N__4831\
        );

    \I__964\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4828\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4834\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__4831\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4828\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__959\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4815\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\
        );

    \I__957\ : InMux
    port map (
            O => \N__4812\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\
        );

    \I__956\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4806\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\
        );

    \I__954\ : InMux
    port map (
            O => \N__4803\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__952\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4794\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\
        );

    \I__950\ : InMux
    port map (
            O => \N__4791\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__949\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4785\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__946\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4776\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i
        );

    \I__944\ : InMux
    port map (
            O => \N__4773\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__942\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4764\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52\
        );

    \I__940\ : InMux
    port map (
            O => \N__4761\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__939\ : InMux
    port map (
            O => \N__4758\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__938\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4752\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__936\ : InMux
    port map (
            O => \N__4749\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__4746\,
            I => \N__4742\
        );

    \I__934\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4737\
        );

    \I__933\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4737\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4737\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2\
        );

    \I__931\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4729\
        );

    \I__930\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4726\
        );

    \I__929\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4723\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4729\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4726\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4723\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63\
        );

    \I__925\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4713\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5\
        );

    \I__923\ : InMux
    port map (
            O => \N__4710\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\
        );

    \I__922\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4704\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\
        );

    \I__920\ : InMux
    port map (
            O => \N__4701\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__919\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4694\
        );

    \I__918\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4691\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4694\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4691\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4686\,
            I => \N__4683\
        );

    \I__914\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4680\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1\
        );

    \I__912\ : InMux
    port map (
            O => \N__4677\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__911\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4671\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__909\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4665\,
            I => \N__4660\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \N__4657\
        );

    \I__906\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4654\
        );

    \I__905\ : Span4Mux_s1_v
    port map (
            O => \N__4660\,
            I => \N__4651\
        );

    \I__904\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4648\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4654\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__4651\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4648\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4641\,
            I => \N__4636\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4640\,
            I => \N__4633\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__4639\,
            I => \N__4629\
        );

    \I__897\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4620\
        );

    \I__896\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4620\
        );

    \I__895\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4620\
        );

    \I__894\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4620\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4620\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\
        );

    \I__892\ : InMux
    port map (
            O => \N__4617\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4614\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\
        );

    \I__890\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4606\
        );

    \I__889\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4603\
        );

    \I__888\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4600\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4606\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4603\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4600\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__884\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4590\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__881\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4580\
        );

    \I__880\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4580\,
            I => \beamY_fastZ0Z_6\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4577\,
            I => \beamY_fastZ0Z_6\
        );

    \I__877\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__876\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4566\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4563\,
            I => \un20_beamy_cry_5_c_RNIHJGZ0Z4\
        );

    \I__873\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4551\
        );

    \I__872\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4551\
        );

    \I__871\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4548\
        );

    \I__870\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4545\
        );

    \I__869\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4542\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4539\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4548\,
            I => \N__4534\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4534\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4542\,
            I => \N__4527\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__4539\,
            I => \N__4527\
        );

    \I__863\ : Span4Mux_h
    port map (
            O => \N__4534\,
            I => \N__4524\
        );

    \I__862\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4519\
        );

    \I__861\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4519\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__4527\,
            I => \beamYZ0Z_6\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__4524\,
            I => \beamYZ0Z_6\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4519\,
            I => \beamYZ0Z_6\
        );

    \I__857\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4509\,
            I => \N__4505\
        );

    \I__855\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4502\
        );

    \I__854\ : Span4Mux_h
    port map (
            O => \N__4505\,
            I => \N__4499\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4502\,
            I => \N__4496\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__4499\,
            I => \un20_beamy_cry_1_c_RNI97CZ0Z4\
        );

    \I__851\ : Odrv12
    port map (
            O => \N__4496\,
            I => \un20_beamy_cry_1_c_RNI97CZ0Z4\
        );

    \I__850\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4484\
        );

    \I__849\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4484\
        );

    \I__848\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4481\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4484\,
            I => \beamY_fastZ0Z_2\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4481\,
            I => \beamY_fastZ0Z_2\
        );

    \I__845\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4472\
        );

    \I__844\ : CEMux
    port map (
            O => \N__4475\,
            I => \N__4464\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4472\,
            I => \N__4461\
        );

    \I__842\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4458\
        );

    \I__841\ : CEMux
    port map (
            O => \N__4470\,
            I => \N__4454\
        );

    \I__840\ : CEMux
    port map (
            O => \N__4469\,
            I => \N__4451\
        );

    \I__839\ : CEMux
    port map (
            O => \N__4468\,
            I => \N__4448\
        );

    \I__838\ : CEMux
    port map (
            O => \N__4467\,
            I => \N__4443\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4464\,
            I => \N__4440\
        );

    \I__836\ : Span4Mux_h
    port map (
            O => \N__4461\,
            I => \N__4435\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4435\
        );

    \I__834\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4432\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4427\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4427\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4448\,
            I => \N__4424\
        );

    \I__830\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4421\
        );

    \I__829\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4418\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4415\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4440\,
            I => \N__4412\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__4435\,
            I => \N__4403\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4432\,
            I => \N__4403\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__4427\,
            I => \N__4403\
        );

    \I__823\ : Span4Mux_s2_v
    port map (
            O => \N__4424\,
            I => \N__4403\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4421\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4418\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__4415\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__4412\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__4403\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__817\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4386\
        );

    \I__816\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4386\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4386\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__4383\,
            I => \N__4380\
        );

    \I__813\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4377\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1\
        );

    \I__811\ : InMux
    port map (
            O => \N__4374\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__810\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4368\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__808\ : InMux
    port map (
            O => \N__4365\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4362\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__805\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4349\
        );

    \I__804\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4346\
        );

    \I__803\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4341\
        );

    \I__802\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4341\
        );

    \I__801\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4334\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4327\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4327\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4327\
        );

    \I__797\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4320\
        );

    \I__796\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4320\
        );

    \I__795\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4320\
        );

    \I__794\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4317\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4334\,
            I => \beamXZ0Z_0\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__4327\,
            I => \beamXZ0Z_0\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4320\,
            I => \beamXZ0Z_0\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4317\,
            I => \beamXZ0Z_0\
        );

    \I__789\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4304\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__4307\,
            I => \N__4301\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4294\
        );

    \I__786\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4291\
        );

    \I__785\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4284\
        );

    \I__784\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4284\
        );

    \I__783\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4284\
        );

    \I__782\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4281\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__4294\,
            I => \beamXZ0Z_1\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4291\,
            I => \beamXZ0Z_1\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4284\,
            I => \beamXZ0Z_1\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4281\,
            I => \beamXZ0Z_1\
        );

    \I__777\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__775\ : Odrv4
    port map (
            O => \N__4266\,
            I => \beamX_RNIBKAZ0Z_1\
        );

    \I__774\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4258\
        );

    \I__773\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4252\
        );

    \I__772\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4252\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4249\
        );

    \I__770\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4246\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4252\,
            I => un5_visiblex_1_n_25
        );

    \I__768\ : Odrv4
    port map (
            O => \N__4249\,
            I => un5_visiblex_1_n_25
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4246\,
            I => un5_visiblex_1_n_25
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__765\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4233\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i
        );

    \I__763\ : InMux
    port map (
            O => \N__4230\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__761\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4221\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0\
        );

    \I__759\ : InMux
    port map (
            O => \N__4218\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\
        );

    \I__758\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__757\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4209\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4209\,
            I => \Pixel_0_sqmuxa_6\
        );

    \I__755\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__754\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4200\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__752\ : Span4Mux_h
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__4194\,
            I => un15_beamy
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4191\,
            I => \Pixel_0_sqmuxa_7_cascade_\
        );

    \I__749\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4185\,
            I => un13_visiblex_4
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__4182\,
            I => \N__4177\
        );

    \I__746\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4173\
        );

    \I__745\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4170\
        );

    \I__744\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4165\
        );

    \I__743\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4162\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4173\,
            I => \N__4157\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4170\,
            I => \N__4157\
        );

    \I__740\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4154\
        );

    \I__739\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4151\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4148\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4162\,
            I => \beamYZ0Z_4\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__4157\,
            I => \beamYZ0Z_4\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4154\,
            I => \beamYZ0Z_4\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4151\,
            I => \beamYZ0Z_4\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__4148\,
            I => \beamYZ0Z_4\
        );

    \I__732\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4130\
        );

    \I__731\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4127\
        );

    \I__730\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4120\
        );

    \I__729\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4115\
        );

    \I__728\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4115\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4130\,
            I => \N__4110\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4127\,
            I => \N__4110\
        );

    \I__725\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4103\
        );

    \I__724\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4103\
        );

    \I__723\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4103\
        );

    \I__722\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4099\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4120\,
            I => \N__4094\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4094\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__4110\,
            I => \N__4089\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4103\,
            I => \N__4089\
        );

    \I__717\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4086\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4099\,
            I => \beamYZ0Z_8\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__4094\,
            I => \beamYZ0Z_8\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__4089\,
            I => \beamYZ0Z_8\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4086\,
            I => \beamYZ0Z_8\
        );

    \I__712\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4073\
        );

    \I__711\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4069\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4062\
        );

    \I__709\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4059\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4069\,
            I => \N__4056\
        );

    \I__707\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4053\
        );

    \I__706\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4050\
        );

    \I__705\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4045\
        );

    \I__704\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4045\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__4062\,
            I => \N__4042\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4059\,
            I => \N__4037\
        );

    \I__701\ : Span4Mux_s1_v
    port map (
            O => \N__4056\,
            I => \N__4037\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4053\,
            I => \beamYZ0Z_7\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4050\,
            I => \beamYZ0Z_7\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4045\,
            I => \beamYZ0Z_7\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__4042\,
            I => \beamYZ0Z_7\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__4037\,
            I => \beamYZ0Z_7\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__694\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4017\
        );

    \I__693\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4010\
        );

    \I__692\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4010\
        );

    \I__691\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4007\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4017\,
            I => \N__4001\
        );

    \I__689\ : InMux
    port map (
            O => \N__4016\,
            I => \N__3998\
        );

    \I__688\ : InMux
    port map (
            O => \N__4015\,
            I => \N__3995\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4010\,
            I => \N__3990\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4007\,
            I => \N__3990\
        );

    \I__685\ : InMux
    port map (
            O => \N__4006\,
            I => \N__3987\
        );

    \I__684\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3982\
        );

    \I__683\ : InMux
    port map (
            O => \N__4004\,
            I => \N__3982\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__4001\,
            I => \beamYZ0Z_3\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3998\,
            I => \beamYZ0Z_3\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3995\,
            I => \beamYZ0Z_3\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__3990\,
            I => \beamYZ0Z_3\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3987\,
            I => \beamYZ0Z_3\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3982\,
            I => \beamYZ0Z_3\
        );

    \I__676\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3966\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3966\,
            I => un1_beamylto9_1
        );

    \I__674\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3958\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \N__3954\
        );

    \I__672\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3949\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3958\,
            I => \N__3944\
        );

    \I__670\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3941\
        );

    \I__669\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3938\
        );

    \I__668\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3933\
        );

    \I__667\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3933\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3949\,
            I => \N__3930\
        );

    \I__665\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3927\
        );

    \I__664\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3924\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__3944\,
            I => \beamYZ0Z_5\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3941\,
            I => \beamYZ0Z_5\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3938\,
            I => \beamYZ0Z_5\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3933\,
            I => \beamYZ0Z_5\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__3930\,
            I => \beamYZ0Z_5\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3927\,
            I => \beamYZ0Z_5\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3924\,
            I => \beamYZ0Z_5\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3909\,
            I => \un1_beamylto9_2_cascade_\
        );

    \I__655\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3899\
        );

    \I__654\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3896\
        );

    \I__653\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3892\
        );

    \I__652\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3889\
        );

    \I__651\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3883\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3899\,
            I => \N__3878\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3896\,
            I => \N__3878\
        );

    \I__648\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3875\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3892\,
            I => \N__3872\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3889\,
            I => \N__3869\
        );

    \I__645\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3864\
        );

    \I__644\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3864\
        );

    \I__643\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3861\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3883\,
            I => \N__3854\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__3878\,
            I => \N__3854\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3875\,
            I => \N__3854\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__3872\,
            I => \beamYZ0Z_9\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__3869\,
            I => \beamYZ0Z_9\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3864\,
            I => \beamYZ0Z_9\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3861\,
            I => \beamYZ0Z_9\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3854\,
            I => \beamYZ0Z_9\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3836\
        );

    \I__632\ : IoInMux
    port map (
            O => \N__3839\,
            I => \N__3833\
        );

    \I__631\ : Span12Mux_s11_v
    port map (
            O => \N__3836\,
            I => \N__3830\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3827\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__3830\,
            I => \VSync_c\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3827\,
            I => \VSync_c\
        );

    \I__627\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3818\
        );

    \I__626\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3815\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3818\,
            I => \N__3808\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3815\,
            I => \N__3808\
        );

    \I__623\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3805\
        );

    \I__622\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3802\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__3808\,
            I => \N__3799\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3805\,
            I => un5_visiblex_1_n_26
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3802\,
            I => un5_visiblex_1_n_26
        );

    \I__618\ : Odrv4
    port map (
            O => \N__3799\,
            I => un5_visiblex_1_n_26
        );

    \I__617\ : InMux
    port map (
            O => \N__3792\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__616\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3785\
        );

    \I__615\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3782\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3785\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3782\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__611\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3771\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0\
        );

    \I__609\ : InMux
    port map (
            O => \N__3768\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__608\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3758\
        );

    \I__607\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3758\
        );

    \I__606\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3755\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3758\,
            I => \beamY_fastZ0Z_3\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3755\,
            I => \beamY_fastZ0Z_3\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3750\,
            I => \N__3746\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__3749\,
            I => \N__3743\
        );

    \I__601\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3737\
        );

    \I__600\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3737\
        );

    \I__599\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3734\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3737\,
            I => \beamY_fastZ0Z_4\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3734\,
            I => \beamY_fastZ0Z_4\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__3729\,
            I => \un5_visibley_ac0_11_0_1_cascade_\
        );

    \I__595\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3723\,
            I => \beamY_fast_RNIGR79Z0Z_7\
        );

    \I__593\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3717\,
            I => \beamY_RNIALEQZ0Z_9\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__3714\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cascade_\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__3711\,
            I => \font_un11_pixellto9_7_0_cascade_\
        );

    \I__589\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3705\,
            I => \N__3701\
        );

    \I__587\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3698\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3698\,
            I => \un8_beamx_cry_1_c_RNITP5AZ0\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3695\,
            I => \un8_beamx_cry_1_c_RNITP5AZ0\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__3690\,
            I => \N__3686\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3689\,
            I => \N__3682\
        );

    \I__581\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3678\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__3685\,
            I => \N__3674\
        );

    \I__579\ : InMux
    port map (
            O => \N__3682\,
            I => \N__3671\
        );

    \I__578\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3668\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3678\,
            I => \N__3665\
        );

    \I__576\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3660\
        );

    \I__575\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3660\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3671\,
            I => \N__3657\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3668\,
            I => \beamYZ0Z_0\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__3665\,
            I => \beamYZ0Z_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3660\,
            I => \beamYZ0Z_0\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__3657\,
            I => \beamYZ0Z_0\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__3648\,
            I => \font_un26_pixel_0_cascade_\
        );

    \I__568\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3641\
        );

    \I__567\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3638\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3641\,
            I => un5_visibley_ac0_11_0_1
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3638\,
            I => un5_visibley_ac0_11_0_1
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__563\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3627\,
            I => un5_visibley_c7
        );

    \I__561\ : InMux
    port map (
            O => \N__3624\,
            I => \N__3621\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__3618\,
            I => \Pixel_0_sqmuxa_4\
        );

    \I__558\ : InMux
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3612\,
            I => font_un11_pixel_0_7
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__3609\,
            I => \un5_visibley_c7_cascade_\
        );

    \I__555\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3603\,
            I => \Pixel_0_sqmuxa_7\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__3600\,
            I => \un5_visibley_c3_cascade_\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3597\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__550\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3588\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3585\,
            I => \N__3581\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__3584\,
            I => \N__3578\
        );

    \I__546\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3575\
        );

    \I__545\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3572\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3575\,
            I => \beamY_fastZ0Z_7\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3572\,
            I => \beamY_fastZ0Z_7\
        );

    \I__542\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3562\
        );

    \I__541\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3557\
        );

    \I__540\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3557\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3562\,
            I => \beamY_fastZ0Z_5\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3557\,
            I => \beamY_fastZ0Z_5\
        );

    \I__537\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3546\
        );

    \I__536\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3546\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3546\,
            I => un5_visibley_c6_0_0_0
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3543\,
            I => \un5_visibley_c6_0_0_0_cascade_\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__532\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3528\
        );

    \I__531\ : InMux
    port map (
            O => \N__3536\,
            I => \N__3528\
        );

    \I__530\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3528\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3528\,
            I => un5_visibley_c3
        );

    \I__528\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3522\,
            I => \beamY_RNIBV5PZ0Z_8\
        );

    \I__526\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3516\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3516\,
            I => un13_visiblex_2
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3513\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3504\
        );

    \I__522\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3504\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3504\,
            I => \N__3498\
        );

    \I__520\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3495\
        );

    \I__519\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3490\
        );

    \I__518\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3490\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__3498\,
            I => un5_visiblex_1_n_23
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3495\,
            I => un5_visiblex_1_n_23
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3490\,
            I => un5_visiblex_1_n_23
        );

    \I__514\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3480\,
            I => \un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0\
        );

    \I__512\ : InMux
    port map (
            O => \N__3477\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\
        );

    \I__511\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3471\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3471\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\
        );

    \I__509\ : InMux
    port map (
            O => \N__3468\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\
        );

    \I__508\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3462\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\
        );

    \I__506\ : InMux
    port map (
            O => \N__3459\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\
        );

    \I__505\ : InMux
    port map (
            O => \N__3456\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\
        );

    \I__504\ : InMux
    port map (
            O => \N__3453\,
            I => \N__3450\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3450\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__502\ : InMux
    port map (
            O => \N__3447\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__3444\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3441\,
            I => \N__3438\
        );

    \I__499\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3435\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3435\,
            I => un5_visiblex_1_n_i_24
        );

    \I__497\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3429\,
            I => \N__3424\
        );

    \I__495\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3421\
        );

    \I__494\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3418\
        );

    \I__493\ : Odrv4
    port map (
            O => \N__3424\,
            I => un5_visiblex_1_n_24
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3421\,
            I => un5_visiblex_1_n_24
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3418\,
            I => un5_visiblex_1_n_24
        );

    \I__490\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3408\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__487\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3399\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0\
        );

    \I__485\ : InMux
    port map (
            O => \N__3396\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__483\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3387\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3387\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0\
        );

    \I__481\ : InMux
    port map (
            O => \N__3384\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__479\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3375\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\
        );

    \I__477\ : InMux
    port map (
            O => \N__3372\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__476\ : InMux
    port map (
            O => \N__3369\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__475\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3363\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3363\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__3360\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\
        );

    \I__472\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3353\
        );

    \I__471\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3350\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3353\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3350\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3345\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3339\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3339\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__465\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3333\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3333\,
            I => un13_visiblex_5
        );

    \I__463\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3327\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3327\,
            I => \Pixel_0_sqmuxa_2\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__3324\,
            I => \un13_visiblex_5_cascade_\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__459\ : InMux
    port map (
            O => \N__3318\,
            I => \N__3309\
        );

    \I__458\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3309\
        );

    \I__457\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3309\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3309\,
            I => un5_visiblex_1_n_31
        );

    \I__455\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3297\
        );

    \I__454\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3297\
        );

    \I__453\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3297\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3297\,
            I => un5_visiblex_1_n_30
        );

    \I__451\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N_159\
        );

    \I__449\ : InMux
    port map (
            O => \N__3288\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__448\ : InMux
    port map (
            O => \N__3285\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__447\ : InMux
    port map (
            O => \N__3282\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__446\ : InMux
    port map (
            O => \N__3279\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__3276\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3267\
        );

    \I__443\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3267\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3267\,
            I => \un20_beamy_cry_4_c_RNIFGFZ0Z4\
        );

    \I__441\ : InMux
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3261\,
            I => un13_visiblex_2_0
        );

    \I__439\ : InMux
    port map (
            O => \N__3258\,
            I => \N__3255\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3255\,
            I => un12_visiblexlt9_0
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__436\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3246\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3246\,
            I => un13_visiblex_0
        );

    \I__434\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3240\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3240\,
            I => font_un7_pixellt9_0
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__3237\,
            I => \font_un14_pixellt9_0_cascade_\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__3234\,
            I => \beamY_fast_RNIGR79Z0Z_7_cascade_\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__429\ : InMux
    port map (
            O => \N__3228\,
            I => \N__3225\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3225\,
            I => \beamY_RNIALEQ_0Z0Z_9\
        );

    \I__427\ : InMux
    port map (
            O => \N__3222\,
            I => \N__3216\
        );

    \I__426\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3216\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3216\,
            I => \un20_beamy_cry_2_c_RNIBADZ0Z4\
        );

    \I__424\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3207\
        );

    \I__423\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3207\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3207\,
            I => \un20_beamy_cry_3_c_RNIDDEZ0Z4\
        );

    \I__421\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3200\
        );

    \I__420\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3197\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3200\,
            I => \un20_beamy_cry_6_c_RNIJMHZ0Z4\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3197\,
            I => \un20_beamy_cry_6_c_RNIJMHZ0Z4\
        );

    \I__417\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3182\
        );

    \I__416\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3179\
        );

    \I__415\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3166\
        );

    \I__414\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3166\
        );

    \I__413\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3166\
        );

    \I__412\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3166\
        );

    \I__411\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3166\
        );

    \I__410\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3166\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3182\,
            I => \beamY_RNI9DLCZ0Z_5\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3179\,
            I => \beamY_RNI9DLCZ0Z_5\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3166\,
            I => \beamY_RNI9DLCZ0Z_5\
        );

    \I__406\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3151\
        );

    \I__405\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3144\
        );

    \I__404\ : InMux
    port map (
            O => \N__3157\,
            I => \N__3144\
        );

    \I__403\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3144\
        );

    \I__402\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3141\
        );

    \I__401\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3138\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3151\,
            I => \beamXZ0Z_7\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3144\,
            I => \beamXZ0Z_7\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3141\,
            I => \beamXZ0Z_7\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3138\,
            I => \beamXZ0Z_7\
        );

    \I__396\ : InMux
    port map (
            O => \N__3129\,
            I => un5_visiblex_1_cry_6
        );

    \I__395\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3120\
        );

    \I__394\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3117\
        );

    \I__393\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3114\
        );

    \I__392\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3111\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3120\,
            I => \beamXZ0Z_8\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3117\,
            I => \beamXZ0Z_8\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3114\,
            I => \beamXZ0Z_8\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3111\,
            I => \beamXZ0Z_8\
        );

    \I__387\ : InMux
    port map (
            O => \N__3102\,
            I => \bfn_6_8_0_\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3099\,
            I => \N__3095\
        );

    \I__385\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3091\
        );

    \I__384\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3088\
        );

    \I__383\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3084\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3091\,
            I => \N__3081\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3088\,
            I => \N__3078\
        );

    \I__380\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3075\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3084\,
            I => \beamXZ0Z_9\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__3081\,
            I => \beamXZ0Z_9\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__3078\,
            I => \beamXZ0Z_9\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3075\,
            I => \beamXZ0Z_9\
        );

    \I__375\ : InMux
    port map (
            O => \N__3066\,
            I => un5_visiblex_1_cry_8
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__3063\,
            I => \un5_visiblex_1_n_23_cascade_\
        );

    \I__373\ : InMux
    port map (
            O => \N__3060\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\
        );

    \I__372\ : InMux
    port map (
            O => \N__3057\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\
        );

    \I__371\ : InMux
    port map (
            O => \N__3054\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__3051\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__369\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__3042\,
            I => un8_beamy
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__365\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3033\,
            I => un4_beamy_0
        );

    \I__363\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3023\
        );

    \I__362\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3023\
        );

    \I__361\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3019\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3023\,
            I => \N__3016\
        );

    \I__359\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3013\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3019\,
            I => \N__3010\
        );

    \I__357\ : Span4Mux_h
    port map (
            O => \N__3016\,
            I => \N__3007\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3013\,
            I => \beamXZ0Z_10\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__3010\,
            I => \beamXZ0Z_10\
        );

    \I__354\ : Odrv4
    port map (
            O => \N__3007\,
            I => \beamXZ0Z_10\
        );

    \I__353\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2991\
        );

    \I__352\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2991\
        );

    \I__351\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2991\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2991\,
            I => un1_beamx_2
        );

    \I__349\ : InMux
    port map (
            O => \N__2988\,
            I => \N__2985\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2985\,
            I => un13_beamylt7
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2982\,
            I => \un15_beamy_2_cascade_\
        );

    \I__346\ : InMux
    port map (
            O => \N__2979\,
            I => un5_visiblex_1_cry_0
        );

    \I__345\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2969\
        );

    \I__344\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2969\
        );

    \I__343\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2965\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2969\,
            I => \N__2962\
        );

    \I__341\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2959\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2965\,
            I => \beamXZ0Z_2\
        );

    \I__339\ : Odrv4
    port map (
            O => \N__2962\,
            I => \beamXZ0Z_2\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2959\,
            I => \beamXZ0Z_2\
        );

    \I__337\ : InMux
    port map (
            O => \N__2952\,
            I => un5_visiblex_1_cry_1
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__2949\,
            I => \N__2943\
        );

    \I__335\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2939\
        );

    \I__334\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2934\
        );

    \I__333\ : InMux
    port map (
            O => \N__2946\,
            I => \N__2934\
        );

    \I__332\ : InMux
    port map (
            O => \N__2943\,
            I => \N__2931\
        );

    \I__331\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2928\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2939\,
            I => \beamXZ0Z_3\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2934\,
            I => \beamXZ0Z_3\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2931\,
            I => \beamXZ0Z_3\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2928\,
            I => \beamXZ0Z_3\
        );

    \I__326\ : InMux
    port map (
            O => \N__2919\,
            I => un5_visiblex_1_cry_2
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2916\,
            I => \N__2912\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2915\,
            I => \N__2908\
        );

    \I__323\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2902\
        );

    \I__322\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2899\
        );

    \I__321\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2892\
        );

    \I__320\ : InMux
    port map (
            O => \N__2907\,
            I => \N__2892\
        );

    \I__319\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2892\
        );

    \I__318\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2889\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2902\,
            I => \beamXZ0Z_4\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2899\,
            I => \beamXZ0Z_4\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2892\,
            I => \beamXZ0Z_4\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2889\,
            I => \beamXZ0Z_4\
        );

    \I__313\ : InMux
    port map (
            O => \N__2880\,
            I => un5_visiblex_1_cry_3
        );

    \I__312\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2869\
        );

    \I__311\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2864\
        );

    \I__310\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2864\
        );

    \I__309\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2861\
        );

    \I__308\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2858\
        );

    \I__307\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2855\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2869\,
            I => \beamXZ0Z_5\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2864\,
            I => \beamXZ0Z_5\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2861\,
            I => \beamXZ0Z_5\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2858\,
            I => \beamXZ0Z_5\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2855\,
            I => \beamXZ0Z_5\
        );

    \I__301\ : InMux
    port map (
            O => \N__2844\,
            I => un5_visiblex_1_cry_4
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2841\,
            I => \N__2835\
        );

    \I__299\ : InMux
    port map (
            O => \N__2840\,
            I => \N__2830\
        );

    \I__298\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2825\
        );

    \I__297\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2825\
        );

    \I__296\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2822\
        );

    \I__295\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2819\
        );

    \I__294\ : InMux
    port map (
            O => \N__2833\,
            I => \N__2816\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2830\,
            I => \beamXZ0Z_6\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2825\,
            I => \beamXZ0Z_6\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2822\,
            I => \beamXZ0Z_6\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2819\,
            I => \beamXZ0Z_6\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2816\,
            I => \beamXZ0Z_6\
        );

    \I__288\ : InMux
    port map (
            O => \N__2805\,
            I => un5_visiblex_1_cry_5
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2802\,
            I => \un4_beamylt6_cascade_\
        );

    \I__286\ : CascadeMux
    port map (
            O => \N__2799\,
            I => \un4_beamylt8_0_cascade_\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__2796\,
            I => \N__2793\
        );

    \I__284\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2790\,
            I => un3_beamx_5
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__2787\,
            I => \un3_beamx_7_cascade_\
        );

    \I__281\ : CascadeMux
    port map (
            O => \N__2784\,
            I => \un1_beamxlt10_0_cascade_\
        );

    \I__280\ : IoInMux
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__278\ : Span4Mux_s2_v
    port map (
            O => \N__2775\,
            I => \N__2771\
        );

    \I__277\ : IoInMux
    port map (
            O => \N__2774\,
            I => \N__2768\
        );

    \I__276\ : Span4Mux_h
    port map (
            O => \N__2771\,
            I => \N__2765\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2768\,
            I => \N__2762\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__2765\,
            I => \N__2759\
        );

    \I__273\ : IoSpan4Mux
    port map (
            O => \N__2762\,
            I => \N__2756\
        );

    \I__272\ : Span4Mux_v
    port map (
            O => \N__2759\,
            I => \N__2753\
        );

    \I__271\ : Span4Mux_s3_v
    port map (
            O => \N__2756\,
            I => \N__2750\
        );

    \I__270\ : Odrv4
    port map (
            O => \N__2753\,
            I => \HSync_c\
        );

    \I__269\ : Odrv4
    port map (
            O => \N__2750\,
            I => \HSync_c\
        );

    \I__268\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2742\,
            I => un18_beamylt10_0
        );

    \I__266\ : InMux
    port map (
            O => \N__2739\,
            I => un20_beamy_cry_7
        );

    \I__265\ : InMux
    port map (
            O => \N__2736\,
            I => \bfn_6_3_0_\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__2733\,
            I => \un5_beamx_4_cascade_\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2730\,
            I => \beamY_RNI9DLCZ0Z_5_cascade_\
        );

    \I__262\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2724\,
            I => un5_beamx_3
        );

    \I__260\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2718\,
            I => un5_beamx_2
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__2715\,
            I => \un5_beamx_2_cascade_\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2712\,
            I => \un8_beamylto9_1_cascade_\
        );

    \I__256\ : InMux
    port map (
            O => \N__2709\,
            I => un8_beamx_cry_9
        );

    \I__255\ : InMux
    port map (
            O => \N__2706\,
            I => un20_beamy_cry_1
        );

    \I__254\ : InMux
    port map (
            O => \N__2703\,
            I => un20_beamy_cry_2
        );

    \I__253\ : InMux
    port map (
            O => \N__2700\,
            I => un20_beamy_cry_3
        );

    \I__252\ : InMux
    port map (
            O => \N__2697\,
            I => un20_beamy_cry_4
        );

    \I__251\ : InMux
    port map (
            O => \N__2694\,
            I => un20_beamy_cry_5
        );

    \I__250\ : InMux
    port map (
            O => \N__2691\,
            I => un20_beamy_cry_6
        );

    \I__249\ : InMux
    port map (
            O => \N__2688\,
            I => un8_beamx_cry_1
        );

    \I__248\ : InMux
    port map (
            O => \N__2685\,
            I => un8_beamx_cry_2
        );

    \I__247\ : InMux
    port map (
            O => \N__2682\,
            I => un8_beamx_cry_3
        );

    \I__246\ : InMux
    port map (
            O => \N__2679\,
            I => un8_beamx_cry_4
        );

    \I__245\ : InMux
    port map (
            O => \N__2676\,
            I => un8_beamx_cry_5
        );

    \I__244\ : InMux
    port map (
            O => \N__2673\,
            I => un8_beamx_cry_6
        );

    \I__243\ : InMux
    port map (
            O => \N__2670\,
            I => un8_beamx_cry_7
        );

    \I__242\ : InMux
    port map (
            O => \N__2667\,
            I => \bfn_5_8_0_\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__2664\,
            I => \un18_beamylto9_2_cascade_\
        );

    \I__240\ : InMux
    port map (
            O => \N__2661\,
            I => \N__2655\
        );

    \I__239\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2655\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2655\,
            I => un18_beamylt4
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2652\,
            I => \N__2649\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2649\,
            I => \N__2646\
        );

    \I__235\ : IoSpan4Mux
    port map (
            O => \N__2646\,
            I => \N__2643\
        );

    \I__234\ : IoSpan4Mux
    port map (
            O => \N__2643\,
            I => \N__2640\
        );

    \I__233\ : IoSpan4Mux
    port map (
            O => \N__2640\,
            I => \N__2637\
        );

    \I__232\ : Odrv4
    port map (
            O => \N__2637\,
            I => \Clock50MHz.PixelClock\
        );

    \I__231\ : IoInMux
    port map (
            O => \N__2634\,
            I => \N__2631\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2631\,
            I => \N__2628\
        );

    \I__229\ : IoSpan4Mux
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__228\ : Odrv4
    port map (
            O => \N__2625\,
            I => \Clock12MHz_c\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_1_cry_7,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un20_beamy_cry_8,
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_3_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2652\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__2975\,
            in1 => \N__4298\,
            in2 => \N__2949\,
            in3 => \N__4338\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4447\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4300\,
            in2 => \_gnd_net_\,
            in3 => \N__4340\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNII5M_9_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3124\,
            in1 => \N__3155\,
            in2 => \N__3099\,
            in3 => \N__2834\,
            lcout => OPEN,
            ltout => \un18_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__2660\,
            in1 => \N__2873\,
            in2 => \N__2664\,
            in3 => \N__2906\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI8P51_4_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__2907\,
            in1 => \N__2661\,
            in2 => \N__2841\,
            in3 => \N__2874\,
            lcout => un13_beamylt7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_10_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4299\,
            in1 => \N__2976\,
            in2 => \N__2915\,
            in3 => \N__3028\,
            lcout => un3_beamx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4352\,
            in2 => \N__4307\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_RNITP5A_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__2688\,
            lcout => \un8_beamx_cry_1_c_RNITP5AZ0\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2948\,
            in2 => \_gnd_net_\,
            in3 => \N__2685\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4476\,
            in1 => \N__2911\,
            in2 => \_gnd_net_\,
            in3 => \N__2682\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2877\,
            in2 => \_gnd_net_\,
            in3 => \N__2679\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2840\,
            in2 => \_gnd_net_\,
            in3 => \N__2676\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3159\,
            in2 => \_gnd_net_\,
            in3 => \N__2673\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3126\,
            in2 => \_gnd_net_\,
            in3 => \N__2670\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__5590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3094\,
            in2 => \_gnd_net_\,
            in3 => \N__2667\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__5589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4471\,
            in1 => \N__3022\,
            in2 => \_gnd_net_\,
            in3 => \N__2709\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3704\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_1_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5726\,
            in2 => \N__3689\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => un20_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_1_c_RNI97C4_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5345\,
            in2 => \_gnd_net_\,
            in3 => \N__2706\,
            lcout => \un20_beamy_cry_1_c_RNI97CZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_1,
            carryout => un20_beamy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_2_c_RNIBAD4_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4016\,
            in2 => \_gnd_net_\,
            in3 => \N__2703\,
            lcout => \un20_beamy_cry_2_c_RNIBADZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_2,
            carryout => un20_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_3_c_RNIDDE4_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4176\,
            in2 => \_gnd_net_\,
            in3 => \N__2700\,
            lcout => \un20_beamy_cry_3_c_RNIDDEZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_3,
            carryout => un20_beamy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_4_c_RNIFGF4_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3957\,
            in2 => \_gnd_net_\,
            in3 => \N__2697\,
            lcout => \un20_beamy_cry_4_c_RNIFGFZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_4,
            carryout => un20_beamy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_5_c_RNIHJG4_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4556\,
            in2 => \_gnd_net_\,
            in3 => \N__2694\,
            lcout => \un20_beamy_cry_5_c_RNIHJGZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_5,
            carryout => un20_beamy_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_6_c_RNIJMH4_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4068\,
            in2 => \_gnd_net_\,
            in3 => \N__2691\,
            lcout => \un20_beamy_cry_6_c_RNIJMHZ0Z4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_6,
            carryout => un20_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_8_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4123\,
            in2 => \_gnd_net_\,
            in3 => \N__2739\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un20_beamy_cry_7,
            carryout => un20_beamy_cry_8,
            clk => \N__5597\,
            ce => \N__4467\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3902\,
            in1 => \N__3191\,
            in2 => \_gnd_net_\,
            in3 => \N__2736\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5595\,
            ce => \N__4468\,
            sr => \_gnd_net_\
        );

    \beamY_RNID825_6_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__2721\,
            in1 => \N__4560\,
            in2 => \_gnd_net_\,
            in3 => \N__4134\,
            lcout => OPEN,
            ltout => \un5_beamx_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_5_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5352\,
            in1 => \N__2727\,
            in2 => \N__2733\,
            in3 => \N__3953\,
            lcout => \beamY_RNI9DLCZ0Z_5\,
            ltout => \beamY_RNI9DLCZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3677\,
            in2 => \N__2730\,
            in3 => \N__4457\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9425_0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5713\,
            in1 => \N__3888\,
            in2 => \N__3685\,
            in3 => \N__4066\,
            lcout => un5_beamx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0H2_4_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4169\,
            in2 => \_gnd_net_\,
            in3 => \N__4015\,
            lcout => un5_beamx_2,
            ltout => \un5_beamx_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5NA6_5_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__5351\,
            in1 => \N__3887\,
            in2 => \N__2715\,
            in3 => \N__3952\,
            lcout => OPEN,
            ltout => \un8_beamylto9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_6_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4065\,
            in1 => \N__4559\,
            in2 => \N__2712\,
            in3 => \N__4133\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5346\,
            lcout => OPEN,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_4_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4180\,
            in1 => \N__3961\,
            in2 => \N__2802\,
            in3 => \N__4557\,
            lcout => OPEN,
            ltout => \un4_beamylt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_7_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__4077\,
            in1 => \N__3903\,
            in2 => \N__2799\,
            in3 => \N__4135\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001001110000"
        )
    port map (
            in0 => \N__4446\,
            in1 => \N__3192\,
            in2 => \N__5730\,
            in3 => \N__3681\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_3_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2838\,
            in1 => \N__2946\,
            in2 => \N__2796\,
            in3 => \N__4358\,
            lcout => OPEN,
            ltout => \un3_beamx_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2999\,
            in1 => \N__3157\,
            in2 => \N__2787\,
            in3 => \N__2875\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_RNO_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2947\,
            in1 => \N__2876\,
            in2 => \N__2916\,
            in3 => \N__2839\,
            lcout => OPEN,
            ltout => \un1_beamxlt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__3158\,
            in1 => \N__3030\,
            in2 => \N__2784\,
            in3 => \N__3000\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3098\,
            in2 => \_gnd_net_\,
            in3 => \N__3125\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIT9ER_10_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2745\,
            in1 => \N__3048\,
            in2 => \N__3039\,
            in3 => \N__3029\,
            lcout => OPEN,
            ltout => \un15_beamy_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNISO4T_7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001010000"
        )
    port map (
            in0 => \N__2998\,
            in1 => \N__2988\,
            in2 => \N__2982\,
            in3 => \N__3156\,
            lcout => un15_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_0_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4337\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => un5_visiblex_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_0_c_RNI1IJC_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4297\,
            in2 => \_gnd_net_\,
            in3 => \N__2979\,
            lcout => un5_visiblex_1_n_31,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_0,
            carryout => un5_visiblex_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_1_c_RNI3LKC_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2968\,
            in2 => \_gnd_net_\,
            in3 => \N__2952\,
            lcout => un5_visiblex_1_n_30,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_1,
            carryout => un5_visiblex_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_2_c_RNI5OLC_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2942\,
            in2 => \N__5458\,
            in3 => \N__2919\,
            lcout => un1_visiblex_24,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_2,
            carryout => un5_visiblex_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_3_c_RNI7RMC_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2905\,
            in2 => \_gnd_net_\,
            in3 => \N__2880\,
            lcout => un5_visiblex_1_n_28,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_3,
            carryout => un5_visiblex_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_4_c_RNI9UNC_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2872\,
            in2 => \_gnd_net_\,
            in3 => \N__2844\,
            lcout => un5_visiblex_1_n_27,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_4,
            carryout => un5_visiblex_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_5_c_RNIB1PC_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2833\,
            in2 => \N__5459\,
            in3 => \N__2805\,
            lcout => un5_visiblex_1_n_26,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_5,
            carryout => un5_visiblex_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_6_c_RNID4QC_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3154\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => un5_visiblex_1_n_25,
            ltout => OPEN,
            carryin => un5_visiblex_1_cry_6,
            carryout => un5_visiblex_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_7_c_RNIF7RC_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3123\,
            in2 => \N__5460\,
            in3 => \N__3102\,
            lcout => un5_visiblex_1_n_24,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => un5_visiblex_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_8_c_RNIHASC_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3087\,
            in2 => \_gnd_net_\,
            in3 => \N__3066\,
            lcout => un5_visiblex_1_n_23,
            ltout => \un5_visiblex_1_n_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_8_c_RNIHASC_1_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3063\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3594\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5411\,
            in2 => \N__3231\,
            in3 => \N__3060\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3720\,
            in2 => \N__5442\,
            in3 => \N__3057\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3051\,
            in3 => \N__4663\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIGR79_7_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4102\,
            in1 => \_gnd_net_\,
            in2 => \N__3585\,
            in3 => \N__3567\,
            lcout => \beamY_fast_RNIGR79Z0Z_7\,
            ltout => \beamY_fast_RNIGR79Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIALEQ_0_9_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3886\,
            in2 => \N__3234\,
            in3 => \N__3644\,
            lcout => \beamY_RNIALEQ_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_3_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3221\,
            in2 => \_gnd_net_\,
            in3 => \N__3185\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_fast_7_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3190\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3204\,
            lcout => \beamY_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_fast_4_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3189\,
            lcout => \beamY_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3272\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_fast_3_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3222\,
            in2 => \_gnd_net_\,
            in3 => \N__3188\,
            lcout => \beamY_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3212\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3203\,
            in2 => \_gnd_net_\,
            in3 => \N__3187\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \beamY_fast_5_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3273\,
            lcout => \beamY_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5598\,
            ce => \N__4469\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_16_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4022\,
            in2 => \_gnd_net_\,
            in3 => \N__5348\,
            lcout => un12_visiblexlt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__3264\,
            in1 => \N__3904\,
            in2 => \N__3633\,
            in3 => \N__3336\,
            lcout => un13_visiblex_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8CP3_1_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011001100"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__4021\,
            in2 => \_gnd_net_\,
            in3 => \N__5347\,
            lcout => font_un7_pixellt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_RNO_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__5704\,
            in1 => \N__4181\,
            in2 => \_gnd_net_\,
            in3 => \N__5349\,
            lcout => un1_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_11_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4262\,
            in1 => \N__3814\,
            in2 => \N__3252\,
            in3 => \N__3509\,
            lcout => un13_visiblex_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_15_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__5140\,
            in1 => \N__3258\,
            in2 => \N__3321\,
            in3 => \N__3306\,
            lcout => un13_visiblex_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIU8361_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__3304\,
            in1 => \N__5136\,
            in2 => \N__4359\,
            in3 => \N__3316\,
            lcout => OPEN,
            ltout => \font_un14_pixellt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIUQF32_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3243\,
            in1 => \N__3813\,
            in2 => \N__3237\,
            in3 => \N__4261\,
            lcout => \Pixel_0_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_4_c_RNIAG3A1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5485\,
            in1 => \N__5231\,
            in2 => \N__5092\,
            in3 => \N__3432\,
            lcout => un13_visiblex_5,
            ltout => \un13_visiblex_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNINUI05_0_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3294\,
            in1 => \N__3330\,
            in2 => \N__3324\,
            in3 => \N__3510\,
            lcout => \Pixel_0_sqmuxa_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIU8361_0_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3317\,
            in1 => \N__4356\,
            in2 => \N__5144\,
            in3 => \N__3305\,
            lcout => \N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4257\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKV_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3366\,
            in2 => \N__3441\,
            in3 => \N__3288\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUD1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3356\,
            in2 => \N__3405\,
            in3 => \N__3285\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISJ3S2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3788\,
            in1 => \N__3342\,
            in2 => \N__3393\,
            in3 => \N__3282\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3357\,
            in1 => \N__3503\,
            in2 => \N__3381\,
            in3 => \N__3279\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3276\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_7_c_RNIF7RC_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3428\,
            lcout => un5_visiblex_1_n_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3427\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3R_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3411\,
            in2 => \_gnd_net_\,
            in3 => \N__3396\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4R_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3483\,
            in2 => \N__5443\,
            in3 => \N__3384\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3502\,
            in2 => \_gnd_net_\,
            in3 => \N__3372\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3369\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3360\,
            in3 => \_gnd_net_\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3345\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_8_c_RNIHASC_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3501\,
            lcout => \un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4609\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250Q_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3525\,
            in2 => \N__5447\,
            in3 => \N__3477\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3474\,
            in2 => \N__5449\,
            in3 => \N__3468\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3465\,
            in2 => \N__5448\,
            in3 => \N__3459\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4664\,
            in3 => \N__3456\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3453\,
            in2 => \_gnd_net_\,
            in3 => \N__3447\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIH1_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__4698\,
            in1 => \_gnd_net_\,
            in2 => \N__3444\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIIGUB_2_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4491\,
            in1 => \_gnd_net_\,
            in2 => \N__3750\,
            in3 => \N__3765\,
            lcout => un5_visibley_c3,
            ltout => \un5_visibley_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIJ9FI_5_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__3566\,
            in1 => \N__4076\,
            in2 => \N__3600\,
            in3 => \N__4532\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_0_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3749\,
            in3 => \N__3764\,
            lcout => OPEN,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010010101"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__4490\,
            in2 => \N__3597\,
            in3 => \N__3551\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIU8LB1_8_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110010"
        )
    port map (
            in0 => \N__3552\,
            in1 => \N__4611\,
            in2 => \N__3540\,
            in3 => \N__4126\,
            lcout => un13_visiblex_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9LFE_6_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__3947\,
            in1 => \N__4533\,
            in2 => \_gnd_net_\,
            in3 => \N__3536\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIRPUB_6_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4583\,
            in2 => \N__3584\,
            in3 => \N__3565\,
            lcout => un5_visibley_c6_0_0_0,
            ltout => \un5_visibley_c6_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBV5P_8_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011010"
        )
    port map (
            in0 => \N__4125\,
            in1 => \_gnd_net_\,
            in2 => \N__3543\,
            in3 => \N__3535\,
            lcout => \beamY_RNIBV5PZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_4_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__4004\,
            in1 => \N__5306\,
            in2 => \N__4182\,
            in3 => \N__3948\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum\,
            ltout => \un1_beamY_if_generate_plus_mult1_un54_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDV6V1_8_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__3519\,
            in1 => \_gnd_net_\,
            in2 => \N__3513\,
            in3 => \N__4846\,
            lcout => \Pixel_0_sqmuxa_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIR3UF_6_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3763\,
            in1 => \N__3742\,
            in2 => \N__4587\,
            in3 => \N__4489\,
            lcout => un5_visibley_ac0_11_0_1,
            ltout => \un5_visibley_ac0_11_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIALEQ_9_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3895\,
            in2 => \N__3729\,
            in3 => \N__3726\,
            lcout => \beamY_RNIALEQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__5307\,
            in1 => \N__4005\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum\,
            ltout => \un1_beamY_if_generate_plus_mult1_un68_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0R15_1_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5731\,
            in2 => \N__3714\,
            in3 => \N__5308\,
            lcout => OPEN,
            ltout => \font_un11_pixellto9_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ0DS_1_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5220\,
            in1 => \N__5183\,
            in2 => \N__3711\,
            in3 => \N__4845\,
            lcout => font_un11_pixel_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_5_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__3708\,
            in1 => \N__4272\,
            in2 => \N__3690\,
            in3 => \N__5818\,
            lcout => OPEN,
            ltout => \font_un26_pixel_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_1_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4206\,
            in1 => \N__4215\,
            in2 => \N__3648\,
            in3 => \N__3606\,
            lcout => \d_N_3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUNJ_7_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__3645\,
            in2 => \N__3962\,
            in3 => \N__4136\,
            lcout => un5_visibley_c7,
            ltout => \un5_visibley_c7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1K0I6_9_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__3624\,
            in1 => \N__3615\,
            in2 => \N__3609\,
            in3 => \N__3905\,
            lcout => \Pixel_0_sqmuxa_7\,
            ltout => \Pixel_0_sqmuxa_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001100"
        )
    port map (
            in0 => \N__4214\,
            in1 => \N__4205\,
            in2 => \N__4191\,
            in3 => \N__4188\,
            lcout => \Pixel_5_N_3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_4_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5326\,
            in1 => \N__4168\,
            in2 => \_gnd_net_\,
            in3 => \N__4006\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_RNO_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4137\,
            in1 => \N__4072\,
            in2 => \N__4026\,
            in3 => \N__4558\,
            lcout => OPEN,
            ltout => \un1_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__3969\,
            in1 => \N__3963\,
            in2 => \N__3909\,
            in3 => \N__3906\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_5_c_RNIB1PC_0_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3822\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3821\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05J52_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4391\,
            in2 => \N__4239\,
            in3 => \N__3792\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEO2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3789\,
            in2 => \N__3777\,
            in3 => \N__3768\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3NMD6_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4733\,
            in1 => \N__4392\,
            in2 => \N__4383\,
            in3 => \N__4374\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4371\,
            in2 => \_gnd_net_\,
            in3 => \N__4365\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4362\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIBKA_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4357\,
            in1 => \N__4308\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamX_RNIBKAZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_6_c_RNID4QC_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4263\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4847\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4593\,
            in2 => \N__4639\,
            in3 => \N__4230\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFV81_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4632\,
            in2 => \N__4227\,
            in3 => \N__4218\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4707\,
            in2 => \N__4640\,
            in3 => \N__4701\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI37VA3_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4913\,
            in1 => \N__4697\,
            in2 => \N__4686\,
            in3 => \N__4677\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4674\,
            in1 => \N__4668\,
            in2 => \N__4641\,
            in3 => \N__4617\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4614\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4610\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_6_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5600\,
            ce => \N__4475\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4571\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5600\,
            ce => \N__4475\,
            sr => \_gnd_net_\
        );

    \beamY_2_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4508\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5600\,
            ce => \N__4475\,
            sr => \_gnd_net_\
        );

    \beamY_fast_2_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4512\,
            lcout => \beamY_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5599\,
            ce => \N__4470\,
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5492\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOS04_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4788\,
            in2 => \N__4782\,
            in3 => \N__4773\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNP5_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4734\,
            in2 => \N__4770\,
            in3 => \N__4761\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_12_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5539\,
            in1 => \N__4716\,
            in2 => \N__4746\,
            in3 => \N__4758\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0R6_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4755\,
            in2 => \_gnd_net_\,
            in3 => \N__4749\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBV5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__4745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4732\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4921\,
            in2 => \N__4821\,
            in3 => \N__4710\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4938\,
            in2 => \N__4926\,
            in3 => \N__4929\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJ22_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4925\,
            in2 => \N__4902\,
            in3 => \N__4890\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI5U736_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5021\,
            in1 => \N__4887\,
            in2 => \N__4878\,
            in3 => \N__4866\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4863\,
            in2 => \_gnd_net_\,
            in3 => \N__4854\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4851\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5230\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONF4_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5016\,
            in2 => \N__5154\,
            in3 => \N__4812\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEV4_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4809\,
            in2 => \N__5022\,
            in3 => \N__4803\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBF5_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5020\,
            in2 => \N__4800\,
            in3 => \N__4791\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIA9BQC_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4971\,
            in1 => \N__5043\,
            in2 => \N__4998\,
            in3 => \N__5037\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5034\,
            in2 => \_gnd_net_\,
            in3 => \N__5028\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6\,
            ltout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_0_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5025\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5015\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5819\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQ6_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4972\,
            in2 => \N__5193\,
            in3 => \N__4989\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85B_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4986\,
            in2 => \N__4977\,
            in3 => \N__4980\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LB_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4976\,
            in2 => \N__4956\,
            in3 => \N__4947\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNI4ON1P_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5875\,
            in1 => \N__4944\,
            in2 => \N__5253\,
            in3 => \N__5244\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSC_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \N__5235\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5232\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_7_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101110011"
        )
    port map (
            in0 => \N__5145\,
            in1 => \N__5073\,
            in2 => \N__5112\,
            in3 => \N__5054\,
            lcout => OPEN,
            ltout => \un19lto10_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_2_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000101010000"
        )
    port map (
            in0 => \N__5055\,
            in1 => \N__5111\,
            in2 => \N__5115\,
            in3 => \N__5502\,
            lcout => un19_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5107\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_13_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5522\,
            in2 => \N__5469\,
            in3 => \N__5067\,
            lcout => \Pixel_1_RNOZ0Z_13\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVA_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5064\,
            in2 => \N__5544\,
            in3 => \N__5046\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5523\,
            in2 => \N__5556\,
            in3 => \N__5540\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_6_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5514\,
            in2 => \_gnd_net_\,
            in3 => \N__5505\,
            lcout => \Pixel_1_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_1_cry_4_c_RNI9UNC_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5496\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__5456\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \N__5350\,
            lcout => \beamY_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_14_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5768\,
            in2 => \_gnd_net_\,
            in3 => \N__5738\,
            lcout => \G_6_i_a4_0_0\,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9D_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5799\,
            in2 => \N__5876\,
            in3 => \N__5277\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00K_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5871\,
            in2 => \N__5274\,
            in3 => \N__5265\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_10_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5262\,
            in2 => \N__5877\,
            in3 => \N__5256\,
            lcout => \Pixel_1_RNOZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5883\,
            in2 => \N__5850\,
            in3 => \N__5867\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAP_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5841\,
            in2 => \_gnd_net_\,
            in3 => \N__5835\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_9_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5832\,
            in1 => \N__5793\,
            in2 => \N__5826\,
            in3 => \N__5781\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5823\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_8_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__5780\,
            in2 => \N__5769\,
            in3 => \N__5745\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_3_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__5739\,
            in1 => \N__5670\,
            in2 => \N__5664\,
            in3 => \N__5661\,
            lcout => OPEN,
            ltout => \un20_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__5655\,
            in1 => \N__5649\,
            in2 => \N__5637\,
            in3 => \N__5634\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5601\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
