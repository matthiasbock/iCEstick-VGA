-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 19 2015 15:42:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal un5_beamx_3 : std_logic;
signal \un5_beamx_4_cascade_\ : std_logic;
signal \beamY_RNIMA24P1Z0Z_5\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_\ : std_logic;
signal \un3_beamx_5_cascade_\ : std_logic;
signal \un3_beamx_7_cascade_\ : std_logic;
signal \beamX_RNI5457Z0Z_5_cascade_\ : std_logic;
signal \un13_beamylto2_0_cascade_\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \N_7_1_cascade_\ : std_logic;
signal g2_1_0 : std_logic;
signal \N_14_cascade_\ : std_logic;
signal \beamY_fast_RNIG57DZ0Z_4_cascade_\ : std_logic;
signal \un5_visibley_c5_cascade_\ : std_logic;
signal \un21_beamy_cry_2_c_RNICOZ0Z83\ : std_logic;
signal \un21_beamy_cry_3_c_RNIERZ0Z93\ : std_logic;
signal \un21_beamy_cry_1_c_RNIALZ0Z73\ : std_logic;
signal \un5_visibley_ac0_11_d_cascade_\ : std_logic;
signal \beamY_fastZ0Z_8\ : std_logic;
signal \beamY_fastZ0Z_4\ : std_logic;
signal \beamY_fast_RNI24GAZ0Z_2_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cascade_\ : std_logic;
signal \beamY_RNI2GUN3Z0Z_9\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_\ : std_logic;
signal \beamY_RNI2GUN3_0Z0Z_9\ : std_logic;
signal d_i4_mux : std_logic;
signal \beamY_RNICDD7FZ0Z_5_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3 : std_logic;
signal \beamY_RNIUBM4FZ0Z_7_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un54_sum_c5 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i : std_logic;
signal \beamY_RNIID28F1_0Z0Z_3_cascade_\ : std_logic;
signal un18_beamylt5_0 : std_logic;
signal \un18_beamylto9_2_cascade_\ : std_logic;
signal \beamY_RNIID28F1Z0Z_3\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_\ : std_logic;
signal g0_0_2_0 : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \beamY_fast_RNIM4P7_0Z0Z_2_cascade_\ : std_logic;
signal \beamY_fast_RNIO71DZ0Z_3\ : std_logic;
signal \beamY_fastZ0Z_2\ : std_logic;
signal \beamY_fast_RNIM4P7Z0Z_2_cascade_\ : std_logic;
signal \beamY_fastZ0Z_3\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \beamY_fast_RNIG57D_0Z0Z_4\ : std_logic;
signal \beamY_fast_RNI45FMZ0Z_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_\ : std_logic;
signal \beamY_RNIK0NV_0Z0Z_9\ : std_logic;
signal un5_visibley_ac0_11_d : std_logic;
signal \un5_visibley_c7_cascade_\ : std_logic;
signal \un21_beamy_cry_8_c_RNIOAFZ0Z3\ : std_logic;
signal \un21_beamy_cry_6_c_RNIK4DZ0Z3\ : std_logic;
signal \un21_beamy_cry_7_c_RNIM7EZ0Z3\ : std_logic;
signal un5_visibley_c5 : std_logic;
signal \beamY_fastZ0Z_9\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6 : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i : std_logic;
signal \beamY_RNI779U3Z0Z_5\ : std_logic;
signal \beamY_RNIUBM4FZ0Z_7\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un61_sum_c4 : std_logic;
signal \beamY_RNI9N7M7Z0Z_5\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal \beamY_RNI5F8A81Z0Z_3_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0 : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_\ : std_logic;
signal \beamY_RNIKUC181_0Z0Z_5\ : std_logic;
signal \beamY_RNIKPNA02Z0Z_5\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3 : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_\ : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un68_sum_c4 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_\ : std_logic;
signal un22_visibleylt9_0_0_0 : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_i : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_\ : std_logic;
signal \un5_visiblex_cry_7_c_RNIVZ0Z952\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \beamY_RNI9KEQ_0Z0Z_8\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\ : std_logic;
signal \beamY_fastZ0Z_7\ : std_logic;
signal un5_visibley_c6_0_0_0 : std_logic;
signal \un11_visibleylto9_1_cascade_\ : std_logic;
signal \un11_visibleylto9_4_cascade_\ : std_logic;
signal \un21_beamy_cry_5_c_RNII1CZ0Z3\ : std_logic;
signal \beamY_fastZ0Z_6\ : std_logic;
signal un5_visibley_c6_0_0 : std_logic;
signal \un21_beamy_cry_4_c_RNIGUAZ0Z3\ : std_logic;
signal \beamY_fastZ0Z_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\ : std_logic;
signal \beamY_RNIECTA3Z0Z_8_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1 : std_logic;
signal un1_beamylto9_2 : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0 : std_logic;
signal \beamY_RNIECTA3Z0Z_8\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un47_sum_c5 : std_logic;
signal \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2 : std_logic;
signal un1_beamylto9_1 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\ : std_logic;
signal \Pixel_1_esr_RNOZ0Z_60\ : std_logic;
signal \g1_0_cascade_\ : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0 : std_logic;
signal \beamY_RNIAJLT9AZ0Z_3\ : std_logic;
signal \r_i1_mux_cascade_\ : std_logic;
signal font_un78_pixellto3 : std_logic;
signal \Pixel_3_sqmuxa_1_1_cascade_\ : std_logic;
signal \G_25_i_a8_0_0\ : std_logic;
signal \Pixel_7_sqmuxa_1_cascade_\ : std_logic;
signal g0_0_0_1 : std_logic;
signal g1 : std_logic;
signal \g0_0_4_0_cascade_\ : std_logic;
signal \N_11\ : std_logic;
signal g0_0_2 : std_logic;
signal \Pixel_3_sqmuxa_1_1\ : std_logic;
signal \N_7_0\ : std_logic;
signal \G_25_i_a8_1_1\ : std_logic;
signal \G_25_i_o8_0_2\ : std_logic;
signal \Pixel_7_sqmuxa_1\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5\ : std_logic;
signal \g0_10_0_cascade_\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \Pixel_9_sn_N_7_mux_1_tz\ : std_logic;
signal \un16_visibleylt9_0_cascade_\ : std_logic;
signal un16_visibley_4 : std_logic;
signal un28_visibleylt9_0 : std_logic;
signal \Pixel_7_sqmuxa_3_0_1\ : std_logic;
signal un22_visibley_3 : std_logic;
signal \un22_visibleylt9_0_cascade_\ : std_logic;
signal un22_visibley_2 : std_logic;
signal un22_visibley : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\ : std_logic;
signal \beamY_fast_RNI1QVSZ0Z_9\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum\ : std_logic;
signal font_un42_pixel_if_generate_plus_mult1_un47_sum_c4 : std_logic;
signal un5_visibley_c2 : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal un5_beamx : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un4_beamylt6 : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \un4_beamylt8_0_cascade_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal un8_beamylto9_1 : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal \Pixel_1_sqmuxa_i_cascade_\ : std_logic;
signal un1_beamx : std_logic;
signal \HSync_c\ : std_logic;
signal un4_beamy_0 : std_logic;
signal un18_beamylt10_0 : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un8_beamy : std_logic;
signal un15_beamy_2 : std_logic;
signal un1_beamx_2 : std_logic;
signal un13_beamylt10_0 : std_logic;
signal \un15_beamy_2_cascade_\ : std_logic;
signal un11_visibley : std_logic;
signal un27lt10 : std_logic;
signal un1_visiblex_27 : std_logic;
signal \Pixel_9_sqmuxa_0_cascade_\ : std_logic;
signal \Pixel_9_sqmuxa\ : std_logic;
signal g0_i_o4_3 : std_logic;
signal \Pixel_9_u_ns_sn\ : std_logic;
signal \N_163_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \Pixel_1_sqmuxa_i_0\ : std_logic;
signal g1_0_0 : std_logic;
signal g0_0_4 : std_logic;
signal \G_25_i_a8_2_0\ : std_logic;
signal \g0_0_5_cascade_\ : std_logic;
signal \G_25_i_3_0\ : std_logic;
signal \N_20\ : std_logic;
signal \G_25_i_2_0_cascade_\ : std_logic;
signal \G_25_i_0\ : std_logic;
signal \Pixel_9_u_ns_rn_0\ : std_logic;
signal g2_1 : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_\ : std_logic;
signal g1_0_1_1 : std_logic;
signal \font_un19_pixel_0_0_0_23_cascade_\ : std_logic;
signal g2_0 : std_logic;
signal g1_0_2 : std_logic;
signal \font_un237_pixel_6_ns_1_0_0_cascade_\ : std_logic;
signal g1_2_0 : std_logic;
signal font_un237_pixel_0_0 : std_logic;
signal \g2_cascade_\ : std_logic;
signal font_un83_pixel_0_0 : std_logic;
signal font_un19_pixel_23 : std_logic;
signal \font_un19_pixel_23_cascade_\ : std_logic;
signal font_un160_pixel_6_1 : std_logic;
signal \g0_1_0_cascade_\ : std_logic;
signal g3_0_0 : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6 : std_logic;
signal g0_i_o4_2 : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \un28lto4_1_cascade_\ : std_logic;
signal \Pixel_1_esr_RNOZ0Z_62\ : std_logic;
signal \un28lt10_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0\ : std_logic;
signal un28_0_1 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5\ : std_logic;
signal \beamY_RNIJ0DBZ0Z_9\ : std_logic;
signal \VSync_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \g1_1_cascade_\ : std_logic;
signal \Pixel_1_esr_RNOZ0Z_39\ : std_logic;
signal \N_1304_0_cascade_\ : std_logic;
signal g1_0_1 : std_logic;
signal \N_17_cascade_\ : std_logic;
signal \G_25_i_a8_1\ : std_logic;
signal \g1_3_cascade_\ : std_logic;
signal \N_1302_0_0_0_cascade_\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \N_159_0_0_cascade_\ : std_logic;
signal \N_156_0\ : std_logic;
signal font_un314_pixel_0 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\ : std_logic;
signal g1_3_0_0 : std_logic;
signal un28lto1 : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal font_un42_pixel_23 : std_logic;
signal \N_1303_0_0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96\ : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9\ : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i : std_logic;
signal un1_visiblex_24 : std_logic;
signal font_un19_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    HSyncDebug <= \HSyncDebug_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__4687\,
            RESETB => \N__9094\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11180\,
            DIN => \N__11179\,
            DOUT => \N__11178\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11180\,
            PADOUT => \N__11179\,
            PADIN => \N__11178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9223\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11171\,
            DIN => \N__11170\,
            DOUT => \N__11169\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11171\,
            PADOUT => \N__11170\,
            PADIN => \N__11169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9855\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11162\,
            DIN => \N__11161\,
            DOUT => \N__11160\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11162\,
            PADOUT => \N__11161\,
            PADIN => \N__11160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8676\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11153\,
            DIN => \N__11152\,
            DOUT => \N__11151\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11153\,
            PADOUT => \N__11152\,
            PADIN => \N__11151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8683\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11144\,
            DIN => \N__11143\,
            DOUT => \N__11142\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11144\,
            PADOUT => \N__11143\,
            PADIN => \N__11142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11135\,
            DIN => \N__11134\,
            DOUT => \N__11133\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11135\,
            PADOUT => \N__11134\,
            PADIN => \N__11133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9859\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11126\,
            DIN => \N__11125\,
            DOUT => \N__11124\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11126\,
            PADOUT => \N__11125\,
            PADIN => \N__11124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2546\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11100\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11097\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11092\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11089\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11086\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11081\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11081\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11078\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11075\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__11092\,
            I => \N__11067\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11089\,
            I => \N__11067\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__11086\,
            I => \N__11067\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__11081\,
            I => \N__11062\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11062\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11075\,
            I => \N__11059\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11056\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__11067\,
            I => \N__11053\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__11062\,
            I => \N__11048\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__11059\,
            I => \N__11048\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11056\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__11053\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__11048\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2524\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11038\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11038\,
            I => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11035\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__2521\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11028\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11025\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11028\,
            I => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__11025\,
            I => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__11020\,
            I => \N__11017\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11014\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__11014\,
            I => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11008\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11008\,
            I => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0\
        );

    \I__2512\ : InMux
    port map (
            O => \N__11005\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__2511\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10999\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10999\,
            I => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__10996\,
            I => \N__10992\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__10995\,
            I => \N__10989\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10984\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10984\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10984\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__2504\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10978\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__2502\ : InMux
    port map (
            O => \N__10975\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__2501\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10969\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10969\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__2499\ : InMux
    port map (
            O => \N__10966\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__10963\,
            I => \N__10959\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10955\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10950\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10950\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10955\,
            I => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10950\,
            I => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10938\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10935\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10929\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10926\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__10941\,
            I => \N__10921\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10938\,
            I => \N__10916\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10916\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__10934\,
            I => \N__10913\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__10933\,
            I => \N__10910\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__10932\,
            I => \N__10907\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10929\,
            I => \N__10904\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10901\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10896\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10896\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10893\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__10916\,
            I => \N__10890\
        );

    \I__2476\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10887\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10882\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10882\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__10904\,
            I => \N__10879\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10901\,
            I => \N__10872\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10872\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10872\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__10890\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10887\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10882\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__10879\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__10872\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__10861\,
            I => \N__10858\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10855\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10855\,
            I => \N__10852\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__10852\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__10849\,
            I => \N__10840\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10837\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10833\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10830\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10824\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10824\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10821\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10817\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10837\,
            I => \N__10814\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10811\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10805\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10805\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10802\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10824\,
            I => \N__10799\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10821\,
            I => \N__10796\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10793\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10790\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__10814\,
            I => \N__10785\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10785\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10782\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__10805\,
            I => \N__10779\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10802\,
            I => \N__10772\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__10799\,
            I => \N__10772\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__10796\,
            I => \N__10772\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10793\,
            I => \N__10765\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__10790\,
            I => \N__10765\
        );

    \I__2434\ : Span4Mux_h
    port map (
            O => \N__10785\,
            I => \N__10765\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10782\,
            I => un1_visiblex_24
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__10779\,
            I => un1_visiblex_24
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__10772\,
            I => un1_visiblex_24
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__10765\,
            I => un1_visiblex_24
        );

    \I__2429\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10753\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10753\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__2427\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10747\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10747\,
            I => g1_0_1
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__10744\,
            I => \N_17_cascade_\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10738\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10738\,
            I => \G_25_i_a8_1\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__10735\,
            I => \g1_3_cascade_\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__10732\,
            I => \N_1302_0_0_0_cascade_\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__10729\,
            I => \N__10719\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10716\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10713\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10710\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10705\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10705\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10700\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10700\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10697\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10716\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10713\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10710\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10705\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10700\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10697\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10678\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10670\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10670\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10667\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10678\,
            I => \N__10664\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10677\,
            I => \N__10659\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10659\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10656\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10670\,
            I => \N__10651\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10651\
        );

    \I__2395\ : Span4Mux_s3_h
    port map (
            O => \N__10664\,
            I => \N__10645\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10659\,
            I => \N__10640\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10640\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10651\,
            I => \N__10637\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__10650\,
            I => \N__10631\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10628\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10625\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__10645\,
            I => \N__10622\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10617\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__10637\,
            I => \N__10617\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10610\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10610\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10610\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10607\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10628\,
            I => \beamXZ0Z_0\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10625\,
            I => \beamXZ0Z_0\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__10622\,
            I => \beamXZ0Z_0\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__10617\,
            I => \beamXZ0Z_0\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10610\,
            I => \beamXZ0Z_0\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10607\,
            I => \beamXZ0Z_0\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__10594\,
            I => \N_159_0_0_cascade_\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10588\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10588\,
            I => \N_156_0\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10582\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10582\,
            I => font_un314_pixel_0
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__10579\,
            I => \N__10568\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__10578\,
            I => \N__10565\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10558\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10558\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10551\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10551\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10551\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10540\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10537\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10534\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10527\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10527\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10527\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10524\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10521\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10516\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10516\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10513\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10506\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10506\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10506\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10501\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10501\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10498\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10493\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10493\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10489\
        );

    \I__2343\ : Span4Mux_s3_h
    port map (
            O => \N__10524\,
            I => \N__10482\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__10521\,
            I => \N__10482\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10516\,
            I => \N__10482\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10479\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10506\,
            I => \N__10474\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10501\,
            I => \N__10474\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__10498\,
            I => \N__10469\
        );

    \I__2336\ : Span4Mux_v
    port map (
            O => \N__10493\,
            I => \N__10469\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10466\
        );

    \I__2334\ : Span4Mux_h
    port map (
            O => \N__10489\,
            I => \N__10461\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__10482\,
            I => \N__10461\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10479\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2331\ : Odrv12
    port map (
            O => \N__10474\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__10469\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10466\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__10461\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \N__10439\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__10449\,
            I => \N__10435\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10432\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__10447\,
            I => \N__10426\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__10446\,
            I => \N__10423\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10419\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10412\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10412\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10412\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10407\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10407\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10400\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10400\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10400\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10395\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10395\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10388\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10388\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10388\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__10419\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10412\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10407\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10400\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10395\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10388\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10372\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10372\,
            I => g1_3_0_0
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__10369\,
            I => \N__10364\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10360\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10347\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10342\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10339\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10360\,
            I => \N__10336\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10333\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10330\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10327\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10324\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__10355\,
            I => \N__10321\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10316\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10311\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10311\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10306\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10306\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10302\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \N__10299\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__10345\,
            I => \N__10296\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__10342\,
            I => \N__10293\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10339\,
            I => \N__10280\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__10336\,
            I => \N__10280\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10333\,
            I => \N__10280\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10330\,
            I => \N__10280\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__10327\,
            I => \N__10280\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10324\,
            I => \N__10280\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10277\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10272\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10272\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10265\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10311\,
            I => \N__10265\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10306\,
            I => \N__10265\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10262\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__10302\,
            I => \N__10258\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10255\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10252\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__10293\,
            I => \N__10247\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__10280\,
            I => \N__10247\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10238\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10238\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__10265\,
            I => \N__10238\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10262\,
            I => \N__10238\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10261\,
            I => \N__10235\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__10258\,
            I => \N__10232\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10255\,
            I => un28lto1
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__10252\,
            I => un28lto1
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__10247\,
            I => un28lto1
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__10238\,
            I => un28lto1
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__10235\,
            I => un28lto1
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__10232\,
            I => un28lto1
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__10219\,
            I => \N__10206\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10203\
        );

    \I__2248\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10200\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10193\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10193\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10193\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10187\
        );

    \I__2243\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10184\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10181\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10176\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10176\
        );

    \I__2239\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10172\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10167\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__10200\,
            I => \N__10167\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10164\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10161\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10158\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__10190\,
            I => \N__10155\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10152\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10145\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__10181\,
            I => \N__10145\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10176\,
            I => \N__10145\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__10175\,
            I => \N__10142\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10139\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__10167\,
            I => \N__10134\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__10164\,
            I => \N__10134\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10161\,
            I => \N__10130\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10158\,
            I => \N__10127\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10124\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__10152\,
            I => \N__10119\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__10145\,
            I => \N__10119\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10116\
        );

    \I__2218\ : Span4Mux_h
    port map (
            O => \N__10139\,
            I => \N__10111\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__10134\,
            I => \N__10111\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10108\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__10130\,
            I => \N__10103\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__10127\,
            I => \N__10103\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10100\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__10119\,
            I => \N__10097\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__10116\,
            I => \N__10092\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__10111\,
            I => \N__10092\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10087\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__10103\,
            I => \N__10087\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__10100\,
            I => \beamYZ0Z_0\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__10097\,
            I => \beamYZ0Z_0\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__10092\,
            I => \beamYZ0Z_0\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__10087\,
            I => \beamYZ0Z_0\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10065\
        );

    \I__2202\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10065\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10060\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10057\
        );

    \I__2199\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10054\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10047\
        );

    \I__2197\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10047\
        );

    \I__2196\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10047\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10043\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__10065\,
            I => \N__10040\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10035\
        );

    \I__2192\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10035\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__10027\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10027\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10054\,
            I => \N__10022\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__10047\,
            I => \N__10022\
        );

    \I__2187\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10019\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10012\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__10040\,
            I => \N__10012\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10012\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10009\
        );

    \I__2182\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10004\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10004\
        );

    \I__2180\ : Span4Mux_h
    port map (
            O => \N__10027\,
            I => \N__10001\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__10022\,
            I => \N__9998\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__10019\,
            I => \N__9995\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__10012\,
            I => \N__9992\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__10009\,
            I => font_un42_pixel_23
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__10004\,
            I => font_un42_pixel_23
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__10001\,
            I => font_un42_pixel_23
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__9998\,
            I => font_un42_pixel_23
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__9995\,
            I => font_un42_pixel_23
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__9992\,
            I => font_un42_pixel_23
        );

    \I__2170\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9976\,
            I => \N_1303_0_0\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__9973\,
            I => \un28lto4_1_cascade_\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9967\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9967\,
            I => \Pixel_1_esr_RNOZ0Z_62\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__9964\,
            I => \un28lt10_cascade_\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9952\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9952\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9952\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9952\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9946\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9946\,
            I => un28_0_1
        );

    \I__2158\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9937\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9937\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9937\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9928\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9928\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9928\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__9925\,
            I => \N__9918\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__9924\,
            I => \N__9915\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9912\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9905\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9905\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9905\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9902\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9912\,
            I => \beamY_i_2\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9905\,
            I => \beamY_i_2\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9902\,
            I => \beamY_i_2\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9892\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9892\,
            I => \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5\
        );

    \I__2140\ : SRMux
    port map (
            O => \N__9889\,
            I => \N__9885\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9882\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9885\,
            I => \N__9879\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9882\,
            I => \N__9876\
        );

    \I__2136\ : Span4Mux_h
    port map (
            O => \N__9879\,
            I => \N__9872\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9876\,
            I => \N__9869\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9866\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__9872\,
            I => \beamY_RNIJ0DBZ0Z_9\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__9869\,
            I => \beamY_RNIJ0DBZ0Z_9\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9866\,
            I => \beamY_RNIJ0DBZ0Z_9\
        );

    \I__2130\ : IoInMux
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9856\,
            I => \N__9852\
        );

    \I__2128\ : IoInMux
    port map (
            O => \N__9855\,
            I => \N__9849\
        );

    \I__2127\ : Span4Mux_s0_v
    port map (
            O => \N__9852\,
            I => \N__9846\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9843\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__9846\,
            I => \N__9840\
        );

    \I__2124\ : IoSpan4Mux
    port map (
            O => \N__9843\,
            I => \N__9837\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__2122\ : Span4Mux_s3_v
    port map (
            O => \N__9837\,
            I => \N__9831\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__9834\,
            I => \VSync_c\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__9831\,
            I => \VSync_c\
        );

    \I__2119\ : ClkMux
    port map (
            O => \N__9826\,
            I => \N__9781\
        );

    \I__2118\ : ClkMux
    port map (
            O => \N__9825\,
            I => \N__9781\
        );

    \I__2117\ : ClkMux
    port map (
            O => \N__9824\,
            I => \N__9781\
        );

    \I__2116\ : ClkMux
    port map (
            O => \N__9823\,
            I => \N__9781\
        );

    \I__2115\ : ClkMux
    port map (
            O => \N__9822\,
            I => \N__9781\
        );

    \I__2114\ : ClkMux
    port map (
            O => \N__9821\,
            I => \N__9781\
        );

    \I__2113\ : ClkMux
    port map (
            O => \N__9820\,
            I => \N__9781\
        );

    \I__2112\ : ClkMux
    port map (
            O => \N__9819\,
            I => \N__9781\
        );

    \I__2111\ : ClkMux
    port map (
            O => \N__9818\,
            I => \N__9781\
        );

    \I__2110\ : ClkMux
    port map (
            O => \N__9817\,
            I => \N__9781\
        );

    \I__2109\ : ClkMux
    port map (
            O => \N__9816\,
            I => \N__9781\
        );

    \I__2108\ : ClkMux
    port map (
            O => \N__9815\,
            I => \N__9781\
        );

    \I__2107\ : ClkMux
    port map (
            O => \N__9814\,
            I => \N__9781\
        );

    \I__2106\ : ClkMux
    port map (
            O => \N__9813\,
            I => \N__9781\
        );

    \I__2105\ : ClkMux
    port map (
            O => \N__9812\,
            I => \N__9781\
        );

    \I__2104\ : GlobalMux
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__2103\ : gio2CtrlBuf
    port map (
            O => \N__9778\,
            I => \PixelClock_g\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__9775\,
            I => \g1_1_cascade_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9769\,
            I => \Pixel_1_esr_RNOZ0Z_39\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \N_1304_0_cascade_\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__9763\,
            I => \N__9755\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9749\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9744\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9744\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9741\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9738\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9733\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9733\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9730\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9727\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9749\,
            I => \N__9720\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9744\,
            I => \N__9720\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9741\,
            I => \N__9715\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9738\,
            I => \N__9712\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9733\,
            I => \N__9709\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9730\,
            I => \N__9704\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9727\,
            I => \N__9704\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9701\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9698\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__9720\,
            I => \N__9695\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9690\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9690\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__9715\,
            I => \N__9685\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__9712\,
            I => \N__9685\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__9709\,
            I => \N__9680\
        );

    \I__2073\ : Span4Mux_h
    port map (
            O => \N__9704\,
            I => \N__9680\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9701\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9698\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__9695\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9690\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__9685\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__9680\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__2066\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9664\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9664\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__2064\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9658\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9658\,
            I => \N__9652\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9649\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9642\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9642\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__9652\,
            I => \N__9633\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9649\,
            I => \N__9633\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9630\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9627\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9624\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9619\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9619\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9616\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9613\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__9633\,
            I => \N__9610\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9630\,
            I => \N__9605\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9605\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__9624\,
            I => \N__9602\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9619\,
            I => \N__9599\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9616\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9613\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__9610\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__9605\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9602\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__9599\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9586\,
            I => \N__9581\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9576\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9569\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9569\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9569\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__9579\,
            I => \N__9566\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9576\,
            I => \N__9556\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9556\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9553\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9550\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__9564\,
            I => \N__9547\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__9563\,
            I => \N__9541\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9534\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9534\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__9556\,
            I => \N__9531\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9553\,
            I => \N__9528\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9550\,
            I => \N__9525\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9522\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9513\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9513\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9513\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9513\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9508\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9508\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9534\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__9531\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__9528\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__9525\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9522\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9513\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9508\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6
        );

    \I__2008\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9490\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9487\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__9487\,
            I => g0_i_o4_2
        );

    \I__2005\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9481\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9481\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9478\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9469\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9466\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9460\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9460\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9457\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9454\,
            I => \N__9451\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9448\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9448\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__9445\,
            I => \N__9440\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__9444\,
            I => \N__9436\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9432\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9423\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9423\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9423\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9423\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9432\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9423\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9415\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__9415\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9409\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9409\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9406\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__9403\,
            I => \g0_1_0_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9397\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9397\,
            I => g3_0_0
        );

    \I__1975\ : InMux
    port map (
            O => \N__9394\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__1974\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9387\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9384\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9387\,
            I => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9384\,
            I => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9373\,
            I => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9370\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__1966\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9364\,
            I => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__9361\,
            I => \N__9357\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__9360\,
            I => \N__9354\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9349\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9349\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9349\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__1959\ : InMux
    port map (
            O => \N__9346\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__1958\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__9340\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__1956\ : InMux
    port map (
            O => \N__9337\,
            I => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__9334\,
            I => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__9331\,
            I => \N__9327\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__9330\,
            I => \N__9324\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9319\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9319\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9319\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__1949\ : InMux
    port map (
            O => \N__9316\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__9313\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9307\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9307\,
            I => g1_0_1_1
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__9304\,
            I => \font_un19_pixel_0_0_0_23_cascade_\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__9298\,
            I => g2_0
        );

    \I__1942\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9292\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__9292\,
            I => g1_0_2
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__9289\,
            I => \font_un237_pixel_6_ns_1_0_0_cascade_\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9283\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9283\,
            I => g1_2_0
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__9280\,
            I => \N__9277\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9274\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__9274\,
            I => font_un237_pixel_0_0
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__9271\,
            I => \g2_cascade_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9265\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9265\,
            I => font_un83_pixel_0_0
        );

    \I__1931\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9259\,
            I => font_un19_pixel_23
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__9256\,
            I => \font_un19_pixel_23_cascade_\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9250\,
            I => \N__9247\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__9247\,
            I => font_un160_pixel_6_1
        );

    \I__1925\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__9235\,
            I => g0_i_o4_3
        );

    \I__1921\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9229\,
            I => \Pixel_9_u_ns_sn\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N_163_cascade_\
        );

    \I__1918\ : IoInMux
    port map (
            O => \N__9223\,
            I => \N__9219\
        );

    \I__1917\ : IoInMux
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9219\,
            I => \N__9213\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9216\,
            I => \N__9210\
        );

    \I__1914\ : Span4Mux_s3_v
    port map (
            O => \N__9213\,
            I => \N__9207\
        );

    \I__1913\ : Span4Mux_s3_v
    port map (
            O => \N__9210\,
            I => \N__9204\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__9207\,
            I => \N__9201\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__9201\,
            I => \Pixel_c\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__9198\,
            I => \Pixel_c\
        );

    \I__1908\ : CEMux
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9190\,
            I => \Pixel_1_sqmuxa_i_0\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__9184\,
            I => g1_0_0
        );

    \I__1904\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__9178\,
            I => g0_0_4
        );

    \I__1902\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9172\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9172\,
            I => \G_25_i_a8_2_0\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__9169\,
            I => \g0_0_5_cascade_\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__9163\,
            I => \G_25_i_3_0\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9157\,
            I => \N_20\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \G_25_i_2_0_cascade_\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9148\,
            I => \G_25_i_0\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9142\,
            I => \Pixel_9_u_ns_rn_0\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9133\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__9133\,
            I => g2_1
        );

    \I__1887\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9127\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9127\,
            I => font_un19_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__1885\ : InMux
    port map (
            O => \N__9124\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__1884\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__9118\,
            I => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9115\,
            I => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__9111\,
            I => \N__9103\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \N__9099\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9096\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9091\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9086\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9086\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9083\
        );

    \I__1873\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9080\
        );

    \I__1872\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9077\
        );

    \I__1871\ : IoInMux
    port map (
            O => \N__9094\,
            I => \N__9072\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9063\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9063\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9063\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9063\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9060\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9057\
        );

    \I__1864\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9054\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__9072\,
            I => \N__9049\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__9063\,
            I => \N__9046\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__9060\,
            I => \N__9039\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9039\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9039\
        );

    \I__1858\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9036\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__9052\,
            I => \N__9032\
        );

    \I__1856\ : Span12Mux_s11_v
    port map (
            O => \N__9049\,
            I => \N__9029\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__9046\,
            I => \N__9022\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__9039\,
            I => \N__9022\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9022\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9019\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9016\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__9029\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__9022\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9019\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__9016\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8997\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8997\
        );

    \I__1844\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8997\
        );

    \I__1843\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8987\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8984\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8981\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8976\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8976\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8973\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8970\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8966\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8963\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8954\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8984\,
            I => \N__8954\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8954\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8976\,
            I => \N__8954\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8973\,
            I => \N__8949\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8949\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8946\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8942\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8963\,
            I => \N__8933\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8954\,
            I => \N__8933\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__8949\,
            I => \N__8933\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8933\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8930\
        );

    \I__1821\ : Odrv12
    port map (
            O => \N__8942\,
            I => \beamYZ0Z_2\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__8933\,
            I => \beamYZ0Z_2\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8930\,
            I => \beamYZ0Z_2\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8915\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8915\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8911\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8908\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8905\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8902\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8911\,
            I => \N__8898\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8895\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__8905\,
            I => \N__8890\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8890\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8883\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__8898\,
            I => \N__8880\
        );

    \I__1806\ : Span4Mux_h
    port map (
            O => \N__8895\,
            I => \N__8875\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__8890\,
            I => \N__8875\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8872\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8865\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8865\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8865\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8883\,
            I => \beamYZ0Z_5\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__8880\,
            I => \beamYZ0Z_5\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__8875\,
            I => \beamYZ0Z_5\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8872\,
            I => \beamYZ0Z_5\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8865\,
            I => \beamYZ0Z_5\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8851\,
            I => un8_beamylto9_1
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__8848\,
            I => \N__8843\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8839\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8835\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8832\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8829\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8839\,
            I => \N__8823\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8820\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8813\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8832\,
            I => \N__8813\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8829\,
            I => \N__8813\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__8828\,
            I => \N__8809\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__8827\,
            I => \N__8804\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__8826\,
            I => \N__8801\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8823\,
            I => \N__8794\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8820\,
            I => \N__8794\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8813\,
            I => \N__8794\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8791\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8788\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8785\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8778\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8778\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8778\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__8794\,
            I => \beamYZ0Z_6\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8791\,
            I => \beamYZ0Z_6\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8788\,
            I => \beamYZ0Z_6\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8785\,
            I => \beamYZ0Z_6\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8778\,
            I => \beamYZ0Z_6\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8760\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8755\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8755\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8752\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8747\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8742\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8755\,
            I => \N__8742\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8752\,
            I => \N__8738\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__8751\,
            I => \N__8734\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8731\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8728\
        );

    \I__1755\ : Span4Mux_h
    port map (
            O => \N__8742\,
            I => \N__8725\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8722\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8738\,
            I => \N__8719\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8714\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8714\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8731\,
            I => \beamYZ0Z_7\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__8728\,
            I => \beamYZ0Z_7\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__8725\,
            I => \beamYZ0Z_7\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8722\,
            I => \beamYZ0Z_7\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__8719\,
            I => \beamYZ0Z_7\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8714\,
            I => \beamYZ0Z_7\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__8701\,
            I => \Pixel_1_sqmuxa_i_cascade_\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__8698\,
            I => \N__8694\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8689\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8689\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__8686\,
            I => un1_beamx
        );

    \I__1738\ : IoInMux
    port map (
            O => \N__8683\,
            I => \N__8680\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8677\
        );

    \I__1736\ : Span4Mux_s2_v
    port map (
            O => \N__8677\,
            I => \N__8673\
        );

    \I__1735\ : IoInMux
    port map (
            O => \N__8676\,
            I => \N__8670\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__8673\,
            I => \N__8667\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8664\
        );

    \I__1732\ : Sp12to4
    port map (
            O => \N__8667\,
            I => \N__8661\
        );

    \I__1731\ : Span4Mux_s3_v
    port map (
            O => \N__8664\,
            I => \N__8658\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__8661\,
            I => \HSync_c\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__8658\,
            I => \HSync_c\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8650\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8650\,
            I => un4_beamy_0
        );

    \I__1726\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__8641\,
            I => un18_beamylt10_0
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__8638\,
            I => \N__8633\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8637\,
            I => \N__8630\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8627\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8624\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8620\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8617\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8624\,
            I => \N__8614\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8611\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8620\,
            I => \N__8608\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__8617\,
            I => \N__8603\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8614\,
            I => \N__8603\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8611\,
            I => \beamXZ0Z_10\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8608\,
            I => \beamXZ0Z_10\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__8603\,
            I => \beamXZ0Z_10\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8593\,
            I => un8_beamy
        );

    \I__1707\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8587\,
            I => un15_beamy_2
        );

    \I__1705\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8578\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8573\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8573\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8570\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8565\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8565\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8570\,
            I => un1_beamx_2
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__8565\,
            I => un1_beamx_2
        );

    \I__1697\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8554\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8554\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__8551\,
            I => un13_beamylt10_0
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__8548\,
            I => \un15_beamy_2_cascade_\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8541\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8538\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8535\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8532\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__8535\,
            I => un11_visibley
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__8532\,
            I => un11_visibley
        );

    \I__1686\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8524\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8524\,
            I => un27lt10
        );

    \I__1684\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8518\,
            I => un1_visiblex_27
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8515\,
            I => \Pixel_9_sqmuxa_0_cascade_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8509\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8509\,
            I => \Pixel_9_sqmuxa\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__8506\,
            I => \N__8501\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8496\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8487\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8487\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8487\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8487\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8496\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8487\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8479\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__8476\,
            I => \N__8471\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8466\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__8474\,
            I => \N__8462\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8458\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8455\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8469\,
            I => \N__8451\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8466\,
            I => \N__8448\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8445\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8440\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8440\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8437\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8434\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8429\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8429\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__8448\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8445\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__8440\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__8437\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8434\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8429\,
            I => \beamY_fast_RNI1QVSZ0Z_9\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8403\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8399\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8394\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8394\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8385\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8385\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8385\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8385\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8378\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8378\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8378\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__8403\,
            I => \N__8374\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8371\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8399\,
            I => \N__8366\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8394\,
            I => \N__8366\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8361\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8361\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8358\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__8374\,
            I => \N__8353\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8353\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__8366\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__8361\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8358\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__8353\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8334\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8334\
        );

    \I__1623\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8328\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8325\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8321\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8318\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8334\,
            I => \N__8315\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8308\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8308\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8308\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8328\,
            I => \N__8303\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8303\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8300\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8321\,
            I => \N__8297\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8318\,
            I => \N__8288\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__8315\,
            I => \N__8288\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8288\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__8303\,
            I => \N__8288\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8300\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__8297\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__8288\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__8272\,
            I => font_un42_pixel_if_generate_plus_mult1_un47_sum_c4
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__8269\,
            I => \N__8266\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8263\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1597\ : Span4Mux_h
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__8257\,
            I => un5_visibley_c2
        );

    \I__1595\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1593\ : CEMux
    port map (
            O => \N__8250\,
            I => \N__8242\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8238\
        );

    \I__1591\ : CEMux
    port map (
            O => \N__8248\,
            I => \N__8235\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__8245\,
            I => \N__8230\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8230\
        );

    \I__1588\ : CEMux
    port map (
            O => \N__8241\,
            I => \N__8225\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8238\,
            I => \N__8219\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8235\,
            I => \N__8219\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__8230\,
            I => \N__8216\
        );

    \I__1584\ : CEMux
    port map (
            O => \N__8229\,
            I => \N__8213\
        );

    \I__1583\ : CEMux
    port map (
            O => \N__8228\,
            I => \N__8210\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8225\,
            I => \N__8207\
        );

    \I__1581\ : CEMux
    port map (
            O => \N__8224\,
            I => \N__8204\
        );

    \I__1580\ : Span4Mux_v
    port map (
            O => \N__8219\,
            I => \N__8196\
        );

    \I__1579\ : Span4Mux_s3_h
    port map (
            O => \N__8216\,
            I => \N__8196\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8196\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8192\
        );

    \I__1576\ : Span4Mux_s3_v
    port map (
            O => \N__8207\,
            I => \N__8187\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8204\,
            I => \N__8187\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8184\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__8196\,
            I => \N__8181\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8178\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__8192\,
            I => \N__8175\
        );

    \I__1570\ : Span4Mux_h
    port map (
            O => \N__8187\,
            I => \N__8172\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8167\
        );

    \I__1568\ : Span4Mux_s3_h
    port map (
            O => \N__8181\,
            I => \N__8167\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8178\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__8175\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__8172\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__8167\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8149\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8146\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8139\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8139\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8139\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8134\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8134\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8128\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__8146\,
            I => \N__8123\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__8139\,
            I => \N__8123\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8134\,
            I => \N__8120\
        );

    \I__1552\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8113\
        );

    \I__1551\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8113\
        );

    \I__1550\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8113\
        );

    \I__1549\ : Odrv12
    port map (
            O => \N__8128\,
            I => un5_beamx
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__8123\,
            I => un5_beamx
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__8120\,
            I => un5_beamx
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__8113\,
            I => un5_beamx
        );

    \I__1545\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8099\
        );

    \I__1544\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8096\
        );

    \I__1543\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8093\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__8099\,
            I => \N__8087\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8087\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8084\
        );

    \I__1539\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8081\
        );

    \I__1538\ : Span4Mux_h
    port map (
            O => \N__8087\,
            I => \N__8078\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__8084\,
            I => \N__8075\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8072\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__8078\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__8075\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__8072\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8056\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8049\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8049\
        );

    \I__1528\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8049\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__8056\,
            I => \N__8041\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__8049\,
            I => \N__8041\
        );

    \I__1525\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8038\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8035\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8030\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__8041\,
            I => \N__8023\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8023\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8023\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8020\
        );

    \I__1518\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8014\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__8030\,
            I => \N__8007\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__8023\,
            I => \N__8007\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__8020\,
            I => \N__8007\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__8019\,
            I => \N__8004\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8018\,
            I => \N__8001\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8017\,
            I => \N__7998\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7993\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__8007\,
            I => \N__7993\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7990\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8001\,
            I => \beamYZ0Z_3\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7998\,
            I => \beamYZ0Z_3\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__7993\,
            I => \beamYZ0Z_3\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7990\,
            I => \beamYZ0Z_3\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7978\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__1502\ : Span4Mux_h
    port map (
            O => \N__7975\,
            I => \N__7972\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7972\,
            I => un4_beamylt6
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7969\,
            I => \un4_beamylt6_cascade_\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7966\,
            I => \N__7962\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7955\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7952\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7948\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7943\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7943\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7940\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7933\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7933\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7951\,
            I => \N__7927\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7948\,
            I => \N__7922\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7922\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7919\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7916\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7913\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__7933\,
            I => \N__7910\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7932\,
            I => \N__7907\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7931\,
            I => \N__7902\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7902\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7893\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__7922\,
            I => \N__7893\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__7919\,
            I => \N__7893\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7893\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7913\,
            I => \beamYZ0Z_4\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7910\,
            I => \beamYZ0Z_4\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7907\,
            I => \beamYZ0Z_4\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7902\,
            I => \beamYZ0Z_4\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__7893\,
            I => \beamYZ0Z_4\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7877\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7874\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7871\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7865\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7862\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7871\,
            I => \N__7859\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7856\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__7869\,
            I => \N__7850\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7846\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__7865\,
            I => \N__7837\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__7862\,
            I => \N__7837\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7859\,
            I => \N__7837\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7856\,
            I => \N__7837\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7832\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7854\,
            I => \N__7832\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7829\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7824\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7824\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7846\,
            I => \beamYZ0Z_8\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7837\,
            I => \beamYZ0Z_8\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7832\,
            I => \beamYZ0Z_8\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7829\,
            I => \beamYZ0Z_8\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7824\,
            I => \beamYZ0Z_8\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__7813\,
            I => \un4_beamylt8_0_cascade_\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7806\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7802\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7806\,
            I => \N__7797\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7794\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7791\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7788\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7782\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__7797\,
            I => \N__7775\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7775\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__7791\,
            I => \N__7775\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7788\,
            I => \N__7772\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7769\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7766\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7763\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7782\,
            I => \beamYZ0Z_9\
        );

    \I__1432\ : Odrv4
    port map (
            O => \N__7775\,
            I => \beamYZ0Z_9\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__7772\,
            I => \beamYZ0Z_9\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7769\,
            I => \beamYZ0Z_9\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7766\,
            I => \beamYZ0Z_9\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7763\,
            I => \beamYZ0Z_9\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7747\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7747\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__7744\,
            I => \N__7741\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7738\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7738\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7735\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7729\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7729\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7726\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7723\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7717\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7717\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7714\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__7711\,
            I => \N__7708\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7705\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7705\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7702\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7693\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7693\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7690\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7684\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7681\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__7678\,
            I => \N__7674\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7677\,
            I => \N__7669\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7659\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7659\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7659\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7654\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7668\,
            I => \N__7654\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__7667\,
            I => \N__7650\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7647\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7659\,
            I => \N__7644\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7654\,
            I => \N__7641\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7636\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7636\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7626\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__7644\,
            I => \N__7626\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__7641\,
            I => \N__7626\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7636\,
            I => \N__7626\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7623\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7626\,
            I => \N__7619\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7616\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7622\,
            I => \N__7613\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__7619\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__7616\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7613\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7600\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__7591\,
            I => un28_visibleylt9_0
        );

    \I__1373\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7585\,
            I => \Pixel_7_sqmuxa_3_0_1\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7582\,
            I => \N__7579\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7576\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__7573\,
            I => \N__7568\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7572\,
            I => \N__7565\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7562\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__7568\,
            I => un22_visibley_3
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7565\,
            I => un22_visibley_3
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7562\,
            I => un22_visibley_3
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__7555\,
            I => \un22_visibleylt9_0_cascade_\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7545\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7545\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7542\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7537\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7537\
        );

    \I__1356\ : Span4Mux_v
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__7534\,
            I => un22_visibley_2
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__7531\,
            I => \N__7528\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7525\,
            I => un22_visibley
        );

    \I__1351\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7511\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7511\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7499\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7499\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7499\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7495\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7492\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7489\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7484\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7484\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7477\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7477\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7477\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7499\,
            I => \N__7474\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7498\,
            I => \N__7471\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7495\,
            I => \N__7466\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7492\,
            I => \N__7466\
        );

    \I__1334\ : Span4Mux_v
    port map (
            O => \N__7489\,
            I => \N__7463\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7484\,
            I => \N__7452\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7477\,
            I => \N__7452\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7474\,
            I => \N__7452\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7452\
        );

    \I__1329\ : Span4Mux_h
    port map (
            O => \N__7466\,
            I => \N__7452\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7463\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7452\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__7447\,
            I => \N__7444\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7441\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7438\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7432\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7429\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__7426\,
            I => \N__7422\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7412\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7412\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7412\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7409\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7406\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7412\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7409\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7406\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7393\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7393\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7390\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7384\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7384\,
            I => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__7381\,
            I => \N__7377\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__7380\,
            I => \N__7374\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7369\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7369\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7369\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__1299\ : InMux
    port map (
            O => \N__7366\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__1298\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7360\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7360\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__1296\ : InMux
    port map (
            O => \N__7357\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__7354\,
            I => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1293\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7344\
        );

    \I__1292\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7341\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7344\,
            I => \N__7338\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__7341\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__7338\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7330\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7330\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7323\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__7326\,
            I => \N__7319\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7315\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7312\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7307\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7307\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__7315\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7312\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7307\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7297\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__1275\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7291\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7288\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__7285\,
            I => \Pixel_9_sn_N_7_mux_1_tz\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__7282\,
            I => \un16_visibleylt9_0_cascade_\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7272\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7275\,
            I => \N__7269\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__7272\,
            I => un16_visibley_4
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7269\,
            I => un16_visibley_4
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__7264\,
            I => \N__7261\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7258\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__7255\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__7243\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7240\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__1256\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7234\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__7234\,
            I => \N__7231\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__7231\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__1253\ : InMux
    port map (
            O => \N__7228\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__1252\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7222\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__7219\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__1249\ : InMux
    port map (
            O => \N__7216\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__1248\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7206\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7206\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7203\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7200\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__7203\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__7200\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__7195\,
            I => \g0_10_0_cascade_\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7189\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__1239\ : InMux
    port map (
            O => \N__7186\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__1238\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7179\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7176\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__7179\,
            I => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7176\,
            I => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7165\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__7165\,
            I => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7162\,
            I => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__1230\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7156\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__7153\,
            I => \N_7_0\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__7141\,
            I => \G_25_i_a8_1_1\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1222\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7128\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7125\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__7128\,
            I => \G_25_i_o8_0_2\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7125\,
            I => \G_25_i_o8_0_2\
        );

    \I__1217\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1216\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7114\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__7114\,
            I => \Pixel_7_sqmuxa_1\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__7111\,
            I => \N__7108\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7105\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7102\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__7102\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\
        );

    \I__1210\ : InMux
    port map (
            O => \N__7099\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__7096\,
            I => \r_i1_mux_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7090\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__7090\,
            I => font_un78_pixellto3
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__7087\,
            I => \Pixel_3_sqmuxa_1_1_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7081\,
            I => \N__7078\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__7078\,
            I => \G_25_i_a8_0_0\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__7075\,
            I => \Pixel_7_sqmuxa_1_cascade_\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__7066\,
            I => \N__7063\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__7060\,
            I => g0_0_0_1
        );

    \I__1196\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__7054\,
            I => g1
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__7051\,
            I => \g0_0_4_0_cascade_\
        );

    \I__1193\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7045\,
            I => \N_11\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__7039\,
            I => g0_0_2
        );

    \I__1189\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7030\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7030\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7030\,
            I => \Pixel_3_sqmuxa_1_1\
        );

    \I__1186\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7016\
        );

    \I__1185\ : InMux
    port map (
            O => \N__7026\,
            I => \N__7016\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7025\,
            I => \N__7016\
        );

    \I__1183\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7011\
        );

    \I__1182\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7011\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__7016\,
            I => \N__7008\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__7011\,
            I => \beamY_RNIECTA3Z0Z_8\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__7008\,
            I => \beamY_RNIECTA3Z0Z_8\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6996\
        );

    \I__1177\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6985\
        );

    \I__1176\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6985\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6985\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6985\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6982\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6977\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6977\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6985\,
            I => font_un42_pixel_if_generate_plus_mult1_un47_sum_c5
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6982\,
            I => font_un42_pixel_if_generate_plus_mult1_un47_sum_c5
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6977\,
            I => font_un42_pixel_if_generate_plus_mult1_un47_sum_c5
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6970\,
            I => \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6964\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2
        );

    \I__1164\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6958\,
            I => un1_beamylto9_1
        );

    \I__1162\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6949\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6949\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6940\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6940\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6940\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6934\,
            I => \Pixel_1_esr_RNOZ0Z_60\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \g1_0_cascade_\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6919\,
            I => un1_beamxlt10_0
        );

    \I__1149\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__6912\,
            I => \N__6904\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6899\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6896\
        );

    \I__1144\ : Span4Mux_h
    port map (
            O => \N__6907\,
            I => \N__6893\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6888\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6888\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6885\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6899\,
            I => \beamXZ0Z_7\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6896\,
            I => \beamXZ0Z_7\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__6893\,
            I => \beamXZ0Z_7\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6888\,
            I => \beamXZ0Z_7\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6885\,
            I => \beamXZ0Z_7\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__6874\,
            I => \N__6869\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6862\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6862\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6862\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6862\,
            I => font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6846\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6846\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6846\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6843\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6846\,
            I => \beamY_RNIAJLT9AZ0Z_3\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6843\,
            I => \beamY_RNIAJLT9AZ0Z_3\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6835\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__1121\ : Span4Mux_h
    port map (
            O => \N__6832\,
            I => \N__6828\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6825\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6828\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6825\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6815\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6812\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6809\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6815\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6812\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6809\,
            I => \beamY_fastZ0Z_6\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6799\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6799\,
            I => \N__6795\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6792\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__6795\,
            I => un5_visibley_c6_0_0
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6792\,
            I => un5_visibley_c6_0_0
        );

    \I__1106\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6784\,
            I => \N__6781\
        );

    \I__1104\ : Span4Mux_h
    port map (
            O => \N__6781\,
            I => \N__6777\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6774\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__6777\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6774\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6763\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6763\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6759\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6754\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__6759\,
            I => \N__6751\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6748\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6745\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6754\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__6751\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6748\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6745\,
            I => \beamY_fastZ0Z_5\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6724\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6721\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6718\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6730\,
            I => \N__6715\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6712\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6709\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6706\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6724\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6721\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6718\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__6715\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6712\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6709\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6706\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6686\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6690\,
            I => \N__6681\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6677\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6674\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6671\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6668\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6681\,
            I => \N__6665\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6662\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6677\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__6674\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6671\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6668\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__6665\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6662\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \beamY_RNIECTA3Z0Z_8_cascade_\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6642\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6639\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6642\,
            I => \N__6632\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6639\,
            I => \N__6632\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6627\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6627\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__6632\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6627\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6616\,
            I => \N__6613\
        );

    \I__1048\ : Odrv12
    port map (
            O => \N__6613\,
            I => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6604\,
            I => un1_beamylto9_2
        );

    \I__1044\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6598\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0
        );

    \I__1042\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6592\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6583\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6580\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6574\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6565\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6562\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \N__6555\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6551\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6548\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6545\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6551\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6548\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6545\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6535\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6532\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6526\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6523\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6520\,
            I => \N__6515\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6505\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6505\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6505\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6505\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6505\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6502\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6496\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6496\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6485\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6482\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6479\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6485\,
            I => \beamY_fastZ0Z_7\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6482\,
            I => \beamY_fastZ0Z_7\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6479\,
            I => \beamY_fastZ0Z_7\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6469\,
            I => un5_visibley_c6_0_0_0
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__6466\,
            I => \un11_visibleylto9_1_cascade_\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \un11_visibleylto9_4_cascade_\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__996\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6454\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6454\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1\
        );

    \I__994\ : InMux
    port map (
            O => \N__6451\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__992\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6442\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1\
        );

    \I__990\ : InMux
    port map (
            O => \N__6439\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__989\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6433\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\
        );

    \I__987\ : InMux
    port map (
            O => \N__6430\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__986\ : InMux
    port map (
            O => \N__6427\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__6424\,
            I => \N__6420\
        );

    \I__984\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6411\
        );

    \I__983\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6411\
        );

    \I__982\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6411\
        );

    \I__981\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6408\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6411\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6408\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__6403\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\
        );

    \I__977\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__6397\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__974\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6388\,
            I => \beamY_RNI9KEQ_0Z0Z_8\
        );

    \I__972\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6382\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0\
        );

    \I__970\ : InMux
    port map (
            O => \N__6379\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\
        );

    \I__969\ : InMux
    port map (
            O => \N__6376\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\
        );

    \I__968\ : InMux
    port map (
            O => \N__6373\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\
        );

    \I__967\ : InMux
    port map (
            O => \N__6370\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__966\ : InMux
    port map (
            O => \N__6367\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__965\ : InMux
    port map (
            O => \N__6364\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__963\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6355\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__960\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6346\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6340\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\
        );

    \I__956\ : InMux
    port map (
            O => \N__6337\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\
        );

    \I__955\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6331\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6331\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__953\ : InMux
    port map (
            O => \N__6328\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__952\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6321\
        );

    \I__951\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6318\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6321\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6318\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__947\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6307\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\
        );

    \I__945\ : InMux
    port map (
            O => \N__6304\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__944\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__943\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6295\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6295\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__940\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6286\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\
        );

    \I__938\ : InMux
    port map (
            O => \N__6283\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__937\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6277\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__935\ : InMux
    port map (
            O => \N__6274\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__934\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6267\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__6270\,
            I => \N__6264\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6267\,
            I => \N__6258\
        );

    \I__931\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6255\
        );

    \I__930\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6249\
        );

    \I__929\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6244\
        );

    \I__928\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6244\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__6258\,
            I => \N__6241\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6238\
        );

    \I__925\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6235\
        );

    \I__924\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6230\
        );

    \I__923\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6230\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__6249\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__921\ : LocalMux
    port map (
            O => \N__6244\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__920\ : Odrv4
    port map (
            O => \N__6241\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__919\ : Odrv12
    port map (
            O => \N__6238\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6235\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6230\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__915\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__6211\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i
        );

    \I__913\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__6205\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__911\ : InMux
    port map (
            O => \N__6202\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6199\,
            I => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_\
        );

    \I__909\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6188\
        );

    \I__908\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6181\
        );

    \I__907\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6181\
        );

    \I__906\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6176\
        );

    \I__905\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6176\
        );

    \I__904\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6173\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6170\
        );

    \I__902\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6167\
        );

    \I__901\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6164\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6181\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6176\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__6173\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__6170\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6167\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6164\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__893\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6144\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__6147\,
            I => \N__6141\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6138\
        );

    \I__890\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6135\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__6138\,
            I => un5_visiblex_i_24
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6135\,
            I => un5_visiblex_i_24
        );

    \I__887\ : InMux
    port map (
            O => \N__6130\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__886\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6123\
        );

    \I__885\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6120\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__6123\,
            I => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__6120\,
            I => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__881\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__6109\,
            I => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0\
        );

    \I__879\ : InMux
    port map (
            O => \N__6106\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__878\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__6100\,
            I => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__6097\,
            I => \N__6093\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__6096\,
            I => \N__6090\
        );

    \I__874\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6085\
        );

    \I__873\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6085\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6085\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__871\ : InMux
    port map (
            O => \N__6082\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__870\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__6076\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__868\ : InMux
    port map (
            O => \N__6073\,
            I => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__6070\,
            I => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_\
        );

    \I__866\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__6064\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\
        );

    \I__864\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__863\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6055\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__6055\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3\
        );

    \I__861\ : InMux
    port map (
            O => \N__6052\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__6049\,
            I => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6043\,
            I => un22_visibleylt9_0_0_0
        );

    \I__857\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6037\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6037\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_i
        );

    \I__855\ : InMux
    port map (
            O => \N__6034\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__854\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6027\
        );

    \I__853\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6024\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__6027\,
            I => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__6024\,
            I => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__849\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__6013\,
            I => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0\
        );

    \I__847\ : InMux
    port map (
            O => \N__6010\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__846\ : InMux
    port map (
            O => \N__6007\,
            I => \N__6004\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__6004\,
            I => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__6001\,
            I => \N__5997\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__6000\,
            I => \N__5994\
        );

    \I__842\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5989\
        );

    \I__841\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5989\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5989\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__839\ : InMux
    port map (
            O => \N__5986\,
            I => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__838\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5977\
        );

    \I__837\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5977\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5977\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__835\ : InMux
    port map (
            O => \N__5974\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__834\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5967\
        );

    \I__833\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5964\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5967\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5964\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__830\ : InMux
    port map (
            O => \N__5959\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5956\,
            I => \N__5953\
        );

    \I__828\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5950\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5\
        );

    \I__826\ : InMux
    port map (
            O => \N__5947\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__825\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5940\
        );

    \I__824\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5937\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5940\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5937\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__820\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5926\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9\
        );

    \I__818\ : InMux
    port map (
            O => \N__5923\,
            I => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__817\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__816\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5911\
        );

    \I__815\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5906\
        );

    \I__814\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5906\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5914\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c5
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5911\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c5
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5906\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c5
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__5899\,
            I => \beamY_RNI5F8A81Z0Z_3_cascade_\
        );

    \I__809\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5887\
        );

    \I__808\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5887\
        );

    \I__807\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5884\
        );

    \I__806\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5879\
        );

    \I__805\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5879\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5887\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5884\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5879\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i
        );

    \I__801\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5869\,
            I => font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__5866\,
            I => \font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_\
        );

    \I__798\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5860\,
            I => \beamY_RNIKUC181_0Z0Z_5\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__795\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__794\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5848\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5848\,
            I => \beamY_RNIKPNA02Z0Z_5\
        );

    \I__792\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__791\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5839\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5839\,
            I => font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3
        );

    \I__789\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5832\
        );

    \I__788\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5829\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5832\,
            I => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5829\,
            I => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__5824\,
            I => \font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_\
        );

    \I__784\ : InMux
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__782\ : Span4Mux_h
    port map (
            O => \N__5815\,
            I => \N__5811\
        );

    \I__781\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5808\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__5811\,
            I => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5808\,
            I => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10\
        );

    \I__778\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5800\,
            I => font_un42_pixel_if_generate_plus_mult1_un68_sum_c4
        );

    \I__776\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5794\,
            I => font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5791\,
            I => \N__5787\
        );

    \I__773\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5782\
        );

    \I__772\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5782\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5782\,
            I => font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__769\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__5767\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i
        );

    \I__765\ : InMux
    port map (
            O => \N__5764\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__764\ : InMux
    port map (
            O => \N__5761\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__763\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5751\
        );

    \I__762\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5751\
        );

    \I__761\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5748\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5751\,
            I => \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5748\,
            I => \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__756\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5730\
        );

    \I__754\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5727\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__5730\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5727\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5722\,
            I => \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__5719\,
            I => \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_\
        );

    \I__749\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__5710\,
            I => font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i
        );

    \I__746\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__745\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5701\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5701\,
            I => \beamY_RNI779U3Z0Z_5\
        );

    \I__743\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5694\
        );

    \I__742\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5691\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5683\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5683\
        );

    \I__739\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5680\
        );

    \I__738\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5675\
        );

    \I__737\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5675\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__5683\,
            I => \beamY_RNIUBM4FZ0Z_7\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5680\,
            I => \beamY_RNIUBM4FZ0Z_7\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5675\,
            I => \beamY_RNIUBM4FZ0Z_7\
        );

    \I__733\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5662\
        );

    \I__732\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5662\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__730\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5653\
        );

    \I__729\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5650\
        );

    \I__728\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5647\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__5656\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5653\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5650\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5647\,
            I => font_un42_pixel_if_generate_plus_mult1_un61_sum_c4
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__5638\,
            I => \N__5634\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__5637\,
            I => \N__5629\
        );

    \I__721\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5624\
        );

    \I__720\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5624\
        );

    \I__719\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5619\
        );

    \I__718\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5619\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5624\,
            I => \beamY_RNI9N7M7Z0Z_5\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5619\,
            I => \beamY_RNI9N7M7Z0Z_5\
        );

    \I__715\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5611\,
            I => \beamY_fast_RNIG57D_0Z0Z_4\
        );

    \I__713\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5605\,
            I => \beamY_fast_RNI45FMZ0Z_7\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__5602\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_\
        );

    \I__710\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5596\,
            I => \beamY_RNIK0NV_0Z0Z_9\
        );

    \I__708\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5590\,
            I => un5_visibley_ac0_11_d
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__5587\,
            I => \un5_visibley_c7_cascade_\
        );

    \I__705\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__5578\,
            I => \N__5574\
        );

    \I__702\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5571\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__5574\,
            I => \un21_beamy_cry_8_c_RNIOAFZ0Z3\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5571\,
            I => \un21_beamy_cry_8_c_RNIOAFZ0Z3\
        );

    \I__699\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5563\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5559\
        );

    \I__697\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5556\
        );

    \I__696\ : Span4Mux_h
    port map (
            O => \N__5559\,
            I => \N__5551\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5551\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__5551\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__693\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5545\,
            I => \N__5541\
        );

    \I__691\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5538\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__5541\,
            I => \N__5533\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5533\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__5533\,
            I => \un21_beamy_cry_7_c_RNIM7EZ0Z3\
        );

    \I__687\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__5524\,
            I => un5_visibley_c5
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__683\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__681\ : Span4Mux_v
    port map (
            O => \N__5512\,
            I => \N__5509\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__5509\,
            I => \beamY_fastZ0Z_9\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__5506\,
            I => \beamY_fast_RNIM4P7_0Z0Z_2_cascade_\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__677\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__675\ : Span4Mux_h
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__5491\,
            I => \beamY_fast_RNIO71DZ0Z_3\
        );

    \I__673\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5479\
        );

    \I__672\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5474\
        );

    \I__671\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5474\
        );

    \I__670\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5471\
        );

    \I__669\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5464\
        );

    \I__668\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5464\
        );

    \I__667\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5464\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5479\,
            I => \beamY_fastZ0Z_2\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5474\,
            I => \beamY_fastZ0Z_2\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5471\,
            I => \beamY_fastZ0Z_2\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5464\,
            I => \beamY_fastZ0Z_2\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \beamY_fast_RNIM4P7Z0Z_2_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5446\
        );

    \I__660\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5440\
        );

    \I__659\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5435\
        );

    \I__658\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5435\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5432\
        );

    \I__656\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5425\
        );

    \I__655\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5425\
        );

    \I__654\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5425\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5440\,
            I => \beamY_fastZ0Z_3\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5435\,
            I => \beamY_fastZ0Z_3\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__5432\,
            I => \beamY_fastZ0Z_3\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5425\,
            I => \beamY_fastZ0Z_3\
        );

    \I__649\ : InMux
    port map (
            O => \N__5416\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\
        );

    \I__648\ : InMux
    port map (
            O => \N__5413\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\
        );

    \I__647\ : InMux
    port map (
            O => \N__5410\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__645\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5401\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__643\ : InMux
    port map (
            O => \N__5398\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__641\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5389\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5389\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\
        );

    \I__639\ : InMux
    port map (
            O => \N__5386\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__637\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5377\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\
        );

    \I__635\ : InMux
    port map (
            O => \N__5374\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__634\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5368\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\
        );

    \I__632\ : InMux
    port map (
            O => \N__5365\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\
        );

    \I__630\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5350\
        );

    \I__629\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5350\
        );

    \I__628\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5350\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5350\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\
        );

    \I__626\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5344\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__623\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5335\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\
        );

    \I__621\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5329\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5329\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf
        );

    \I__619\ : InMux
    port map (
            O => \N__5326\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__618\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5320\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\
        );

    \I__616\ : InMux
    port map (
            O => \N__5317\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__615\ : InMux
    port map (
            O => \N__5314\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__614\ : InMux
    port map (
            O => \N__5311\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__5308\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__5305\,
            I => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_\
        );

    \I__611\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5299\,
            I => g0_0_2_0
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__5296\,
            I => \N__5293\
        );

    \I__608\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5290\,
            I => font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf
        );

    \I__606\ : InMux
    port map (
            O => \N__5287\,
            I => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__605\ : InMux
    port map (
            O => \N__5284\,
            I => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__604\ : InMux
    port map (
            O => \N__5281\,
            I => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__603\ : InMux
    port map (
            O => \N__5278\,
            I => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5269\
        );

    \I__601\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5266\
        );

    \I__600\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5261\
        );

    \I__599\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5261\
        );

    \I__598\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5258\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5266\,
            I => \beamXZ0Z_2\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5261\,
            I => \beamXZ0Z_2\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5258\,
            I => \beamXZ0Z_2\
        );

    \I__594\ : InMux
    port map (
            O => \N__5251\,
            I => un5_visiblex_cry_1
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__5248\,
            I => \N__5241\
        );

    \I__592\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5238\
        );

    \I__591\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5231\
        );

    \I__590\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5231\
        );

    \I__589\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5231\
        );

    \I__588\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5228\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5238\,
            I => \beamXZ0Z_3\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5231\,
            I => \beamXZ0Z_3\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__5228\,
            I => \beamXZ0Z_3\
        );

    \I__584\ : InMux
    port map (
            O => \N__5221\,
            I => un5_visiblex_cry_2
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5218\,
            I => \N__5211\
        );

    \I__582\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5208\
        );

    \I__581\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5205\
        );

    \I__580\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5200\
        );

    \I__579\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5200\
        );

    \I__578\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5197\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__5208\,
            I => \beamXZ0Z_4\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5205\,
            I => \beamXZ0Z_4\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5200\,
            I => \beamXZ0Z_4\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__5197\,
            I => \beamXZ0Z_4\
        );

    \I__573\ : InMux
    port map (
            O => \N__5188\,
            I => un5_visiblex_cry_3
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__5185\,
            I => \N__5179\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__5184\,
            I => \N__5174\
        );

    \I__570\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5171\
        );

    \I__569\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5168\
        );

    \I__568\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5165\
        );

    \I__567\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5160\
        );

    \I__566\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5160\
        );

    \I__565\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5157\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__5171\,
            I => \beamXZ0Z_5\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5168\,
            I => \beamXZ0Z_5\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5165\,
            I => \beamXZ0Z_5\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5160\,
            I => \beamXZ0Z_5\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5157\,
            I => \beamXZ0Z_5\
        );

    \I__559\ : InMux
    port map (
            O => \N__5146\,
            I => un5_visiblex_cry_4
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__5143\,
            I => \N__5135\
        );

    \I__557\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5132\
        );

    \I__556\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5127\
        );

    \I__555\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5127\
        );

    \I__554\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5122\
        );

    \I__553\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5122\
        );

    \I__552\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5119\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__5132\,
            I => \beamXZ0Z_6\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__5127\,
            I => \beamXZ0Z_6\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__5122\,
            I => \beamXZ0Z_6\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5119\,
            I => \beamXZ0Z_6\
        );

    \I__547\ : InMux
    port map (
            O => \N__5110\,
            I => un5_visiblex_cry_5
        );

    \I__546\ : InMux
    port map (
            O => \N__5107\,
            I => un5_visiblex_cry_6
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__544\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5095\
        );

    \I__543\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5092\
        );

    \I__542\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5089\
        );

    \I__541\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5086\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5095\,
            I => \beamXZ0Z_8\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__5092\,
            I => \beamXZ0Z_8\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__5089\,
            I => \beamXZ0Z_8\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__5086\,
            I => \beamXZ0Z_8\
        );

    \I__536\ : InMux
    port map (
            O => \N__5077\,
            I => \bfn_5_10_0_\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__5074\,
            I => \N__5070\
        );

    \I__534\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5066\
        );

    \I__533\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5063\
        );

    \I__532\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5059\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5066\,
            I => \N__5054\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__5063\,
            I => \N__5054\
        );

    \I__529\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5051\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__5059\,
            I => \beamXZ0Z_9\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__5054\,
            I => \beamXZ0Z_9\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__5051\,
            I => \beamXZ0Z_9\
        );

    \I__525\ : InMux
    port map (
            O => \N__5044\,
            I => un5_visiblex_cry_8
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__5041\,
            I => \beamY_RNIID28F1_0Z0Z_3_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__522\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5032\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__5032\,
            I => un18_beamylt5_0
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__5029\,
            I => \un18_beamylto9_2_cascade_\
        );

    \I__519\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__5023\,
            I => \beamY_RNIID28F1Z0Z_3\
        );

    \I__517\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5015\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__5019\,
            I => \N__5012\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__5018\,
            I => \N__5007\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5015\,
            I => \N__5004\
        );

    \I__513\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5001\
        );

    \I__512\ : InMux
    port map (
            O => \N__5011\,
            I => \N__4996\
        );

    \I__511\ : InMux
    port map (
            O => \N__5010\,
            I => \N__4996\
        );

    \I__510\ : InMux
    port map (
            O => \N__5007\,
            I => \N__4993\
        );

    \I__509\ : Odrv4
    port map (
            O => \N__5004\,
            I => \beamXZ0Z_1\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__5001\,
            I => \beamXZ0Z_1\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4996\,
            I => \beamXZ0Z_1\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4993\,
            I => \beamXZ0Z_1\
        );

    \I__505\ : InMux
    port map (
            O => \N__4984\,
            I => un5_visiblex_cry_0
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__4981\,
            I => \beamY_RNICDD7FZ0Z_5_cascade_\
        );

    \I__503\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4974\
        );

    \I__502\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4971\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4966\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4971\,
            I => \N__4966\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4966\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4963\,
            I => \beamY_RNIUBM4FZ0Z_7_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4956\
        );

    \I__496\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4953\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4956\,
            I => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4953\,
            I => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__492\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4942\,
            I => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__4939\,
            I => \N__4933\
        );

    \I__489\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4921\
        );

    \I__488\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4921\
        );

    \I__487\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4921\
        );

    \I__486\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4921\
        );

    \I__485\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4921\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4921\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_c5
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__4918\,
            I => \N__4914\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__4917\,
            I => \N__4910\
        );

    \I__481\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4900\
        );

    \I__480\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4900\
        );

    \I__479\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4900\
        );

    \I__478\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4900\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4900\,
            I => font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__475\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4891\,
            I => \beamY_fastZ0Z_8\
        );

    \I__473\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4883\
        );

    \I__472\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4878\
        );

    \I__471\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4878\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4883\,
            I => \beamY_fastZ0Z_4\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4878\,
            I => \beamY_fastZ0Z_4\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \beamY_fast_RNI24GAZ0Z_2_cascade_\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__4870\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cascade_\
        );

    \I__466\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4864\,
            I => \beamY_RNI2GUN3Z0Z_9\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__4861\,
            I => \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_\
        );

    \I__463\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4855\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4855\,
            I => \beamY_RNI2GUN3_0Z0Z_9\
        );

    \I__461\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4849\,
            I => d_i4_mux
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__4846\,
            I => \beamY_fast_RNIG57DZ0Z_4_cascade_\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \un5_visibley_c5_cascade_\
        );

    \I__457\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4836\
        );

    \I__456\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4833\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4836\,
            I => \N__4830\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4833\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__4830\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__452\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4819\
        );

    \I__451\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4819\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4819\,
            I => \un21_beamy_cry_3_c_RNIERZ0Z93\
        );

    \I__449\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4813\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4813\,
            I => \N__4809\
        );

    \I__447\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__4809\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4806\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4801\,
            I => \un5_visibley_ac0_11_d_cascade_\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__4798\,
            I => \N_7_1_cascade_\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__441\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4789\,
            I => g2_1_0
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \N_14_cascade_\
        );

    \I__438\ : InMux
    port map (
            O => \N__4783\,
            I => un8_beamx_cry_1
        );

    \I__437\ : InMux
    port map (
            O => \N__4780\,
            I => un8_beamx_cry_2
        );

    \I__436\ : InMux
    port map (
            O => \N__4777\,
            I => un8_beamx_cry_3
        );

    \I__435\ : InMux
    port map (
            O => \N__4774\,
            I => un8_beamx_cry_4
        );

    \I__434\ : InMux
    port map (
            O => \N__4771\,
            I => un8_beamx_cry_5
        );

    \I__433\ : InMux
    port map (
            O => \N__4768\,
            I => un8_beamx_cry_6
        );

    \I__432\ : InMux
    port map (
            O => \N__4765\,
            I => un8_beamx_cry_7
        );

    \I__431\ : InMux
    port map (
            O => \N__4762\,
            I => \bfn_4_10_0_\
        );

    \I__430\ : InMux
    port map (
            O => \N__4759\,
            I => un8_beamx_cry_9
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4756\,
            I => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__4753\,
            I => \un3_beamx_5_cascade_\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4750\,
            I => \un3_beamx_7_cascade_\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4747\,
            I => \beamX_RNI5457Z0Z_5_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4744\,
            I => \un13_beamylto2_0_cascade_\
        );

    \I__424\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4738\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4738\,
            I => un5_beamx_3
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4735\,
            I => \un5_beamx_4_cascade_\
        );

    \I__421\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4729\,
            I => \beamY_RNIMA24P1Z0Z_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__4726\,
            I => un21_beamy_cry_2
        );

    \I__418\ : InMux
    port map (
            O => \N__4723\,
            I => un21_beamy_cry_3
        );

    \I__417\ : InMux
    port map (
            O => \N__4720\,
            I => un21_beamy_cry_4
        );

    \I__416\ : InMux
    port map (
            O => \N__4717\,
            I => un21_beamy_cry_5
        );

    \I__415\ : InMux
    port map (
            O => \N__4714\,
            I => un21_beamy_cry_6
        );

    \I__414\ : InMux
    port map (
            O => \N__4711\,
            I => un21_beamy_cry_7
        );

    \I__413\ : InMux
    port map (
            O => \N__4708\,
            I => \bfn_4_4_0_\
        );

    \I__412\ : IoInMux
    port map (
            O => \N__4705\,
            I => \N__4702\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__410\ : IoSpan4Mux
    port map (
            O => \N__4699\,
            I => \N__4696\
        );

    \I__409\ : IoSpan4Mux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__4690\,
            I => \Clock50MHz.PixelClock\
        );

    \I__406\ : IoInMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__404\ : IoSpan4Mux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__403\ : Odrv4
    port map (
            O => \N__4678\,
            I => \Clock12MHz_c\
        );

    \I__402\ : InMux
    port map (
            O => \N__4675\,
            I => un21_beamy_cry_1
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4705\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10367\,
            in2 => \N__10190\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_RNIAL73_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8990\,
            in2 => \_gnd_net_\,
            in3 => \N__4675\,
            lcout => \un21_beamy_cry_1_c_RNIALZ0Z73\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_2_c_RNICO83_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8046\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => \un21_beamy_cry_2_c_RNICOZ0Z83\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_3_c_RNIER93_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7938\,
            in2 => \_gnd_net_\,
            in3 => \N__4723\,
            lcout => \un21_beamy_cry_3_c_RNIERZ0Z93\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_4_c_RNIGUA3_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8901\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \un21_beamy_cry_4_c_RNIGUAZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_5_c_RNII1C3_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8838\,
            in2 => \_gnd_net_\,
            in3 => \N__4717\,
            lcout => \un21_beamy_cry_5_c_RNII1CZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_6_c_RNIK4D3_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8763\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \un21_beamy_cry_6_c_RNIK4DZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_7_c_RNIM7E3_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7881\,
            in2 => \_gnd_net_\,
            in3 => \N__4711\,
            lcout => \un21_beamy_cry_7_c_RNIM7EZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_8_c_RNIOAF3_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7810\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => \un21_beamy_cry_8_c_RNIOAFZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__8157\,
            in1 => \N__8249\,
            in2 => \_gnd_net_\,
            in3 => \N__10133\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_5_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110011"
        )
    port map (
            in0 => \N__8945\,
            in1 => \N__8889\,
            in2 => \N__8019\,
            in3 => \N__7932\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_3_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__8248\,
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8017\,
            in2 => \_gnd_net_\,
            in3 => \N__8992\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_9_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8133\,
            in2 => \_gnd_net_\,
            in3 => \N__5577\,
            lcout => \beamY_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__8248\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9817\,
            ce => \N__8248\,
            sr => \_gnd_net_\
        );

    \beamY_RNIC725_9_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8018\,
            in1 => \N__7805\,
            in2 => \N__10369\,
            in3 => \N__8750\,
            lcout => un5_beamx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5025_5_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8993\,
            in1 => \N__8847\,
            in2 => \N__10175\,
            in3 => \N__8920\,
            lcout => OPEN,
            ltout => \un5_beamx_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_8_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4741\,
            in1 => \N__7951\,
            in2 => \N__4735\,
            in3 => \N__7882\,
            lcout => un5_beamx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMA24P1_5_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__5690\,
            in1 => \N__5660\,
            in2 => \N__4948\,
            in3 => \N__7509\,
            lcout => \beamY_RNIMA24P1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMM6891_5_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001011010"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__6646\,
            in2 => \N__5740\,
            in3 => \N__7510\,
            lcout => OPEN,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPFUEA4_3_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101000001"
        )
    port map (
            in0 => \N__4732\,
            in1 => \N__5919\,
            in2 => \N__4756\,
            in3 => \N__8033\,
            lcout => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI6PL_3_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5245\,
            in1 => \N__5215\,
            in2 => \N__5185\,
            in3 => \N__5140\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5073\,
            in2 => \_gnd_net_\,
            in3 => \N__5102\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_10_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5216\,
            in1 => \N__5273\,
            in2 => \N__8637\,
            in3 => \N__5011\,
            lcout => OPEN,
            ltout => \un3_beamx_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_3_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__5246\,
            in2 => \N__4753\,
            in3 => \N__10635\,
            lcout => OPEN,
            ltout => \un3_beamx_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8581\,
            in1 => \N__6910\,
            in2 => \N__4750\,
            in3 => \N__5182\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => \beamX_RNI5457Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4747\,
            in3 => \N__10636\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIDMA_1_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5272\,
            in2 => \_gnd_net_\,
            in3 => \N__5010\,
            lcout => OPEN,
            ltout => \un13_beamylto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIJQQ_3_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__5214\,
            in1 => \N__5244\,
            in2 => \N__4744\,
            in3 => \N__10634\,
            lcout => un18_beamylt5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10648\,
            in2 => \N__5019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5274\,
            in2 => \_gnd_net_\,
            in3 => \N__4783\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5247\,
            in2 => \_gnd_net_\,
            in3 => \N__4780\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8195\,
            in1 => \N__5217\,
            in2 => \_gnd_net_\,
            in3 => \N__4777\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5183\,
            in2 => \_gnd_net_\,
            in3 => \N__4774\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5142\,
            in2 => \_gnd_net_\,
            in3 => \N__4771\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6911\,
            in2 => \_gnd_net_\,
            in3 => \N__4768\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5103\,
            in2 => \_gnd_net_\,
            in3 => \N__4765\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__9812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5069\,
            in2 => \_gnd_net_\,
            in3 => \N__4762\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__9813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8623\,
            in1 => \N__8203\,
            in2 => \_gnd_net_\,
            in3 => \N__4759\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_66_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001110"
        )
    port map (
            in0 => \N__10810\,
            in1 => \N__9725\,
            in2 => \N__4795\,
            in3 => \N__9638\,
            lcout => OPEN,
            ltout => \N_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_51_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4798\,
            in3 => \N__5302\,
            lcout => g0_0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_70_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10492\,
            in2 => \_gnd_net_\,
            in3 => \N__11074\,
            lcout => g2_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_53_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__10820\,
            in1 => \N__10572\,
            in2 => \_gnd_net_\,
            in3 => \N__11096\,
            lcout => OPEN,
            ltout => \N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_30_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__9648\,
            in1 => \_gnd_net_\,
            in2 => \N__4786\,
            in3 => \N__9759\,
            lcout => \G_25_i_a8_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9647\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4812\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__8241\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6780\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__8241\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6831\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => \N__8241\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIG57D_4_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__6768\,
            in1 => \N__4888\,
            in2 => \N__8828\,
            in3 => \N__5488\,
            lcout => OPEN,
            ltout => \beamY_fast_RNIG57DZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIQQEM_5_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__8812\,
            in1 => \N__6769\,
            in2 => \N__4846\,
            in3 => \N__5451\,
            lcout => un5_visibley_c5,
            ltout => \un5_visibley_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIK3TH2_7_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100010010"
        )
    port map (
            in0 => \N__8741\,
            in1 => \N__6733\,
            in2 => \N__4843\,
            in3 => \N__6684\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_4_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8156\,
            lcout => \beamY_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__8224\,
            sr => \_gnd_net_\
        );

    \beamY_fast_3_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4839\,
            lcout => \beamY_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__8224\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8154\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => \N__8224\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIBVU7_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5445\,
            in2 => \_gnd_net_\,
            in3 => \N__5484\,
            lcout => un5_visibley_c2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__8228\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIT5UF_8_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4886\,
            in1 => \N__5443\,
            in2 => \N__4897\,
            in3 => \N__5482\,
            lcout => un5_visibley_ac0_11_d,
            ltout => \un5_visibley_ac0_11_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI45FM_7_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__6488\,
            in1 => \N__7785\,
            in2 => \N__4801\,
            in3 => \N__7849\,
            lcout => \beamY_fast_RNI45FMZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_8_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5544\,
            lcout => \beamY_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => \N__8228\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIG57D_0_4_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__4887\,
            in1 => \N__5444\,
            in2 => \N__7869\,
            in3 => \N__5483\,
            lcout => \beamY_fast_RNIG57D_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI24GA_2_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__7939\,
            in1 => \N__5452\,
            in2 => \N__8751\,
            in3 => \N__5485\,
            lcout => OPEN,
            ltout => \beamY_fast_RNI24GAZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGTNJ_7_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8737\,
            in2 => \N__4873\,
            in3 => \N__6802\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum\,
            ltout => \un1_beamY_if_generate_plus_mult1_un40_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2GUN3_9_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001000010110"
        )
    port map (
            in0 => \N__8461\,
            in1 => \N__5757\,
            in2 => \N__4870\,
            in3 => \N__8406\,
            lcout => \beamY_RNI2GUN3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIO3Q1A_7_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4977\,
            in1 => \N__4858\,
            in2 => \_gnd_net_\,
            in3 => \N__4867\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNITVFT2_3_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000100"
        )
    port map (
            in0 => \N__8333\,
            in1 => \N__8454\,
            in2 => \N__5503\,
            in3 => \N__6685\,
            lcout => OPEN,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI47PR6_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__4852\,
            in1 => \N__6691\,
            in2 => \N__4861\,
            in3 => \N__6734\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un54_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2GUN3_0_9_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110111101001"
        )
    port map (
            in0 => \N__8332\,
            in1 => \N__5758\,
            in2 => \N__8474\,
            in3 => \N__8407\,
            lcout => \beamY_RNI2GUN3_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIAI342_9_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100010000101"
        )
    port map (
            in0 => \N__8408\,
            in1 => \N__7498\,
            in2 => \N__8469\,
            in3 => \N__8331\,
            lcout => d_i4_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDRE6H_0_3_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__7507\,
            in1 => \N__7653\,
            in2 => \N__4918\,
            in3 => \N__4938\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICDD7F_5_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5733\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__7508\,
            lcout => OPEN,
            ltout => \beamY_RNICDD7FZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRJ4CH2_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__7981\,
            in1 => \N__4960\,
            in2 => \N__4981\,
            in3 => \N__5920\,
            lcout => \font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUBM4F_7_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4978\,
            in1 => \N__8281\,
            in2 => \N__4939\,
            in3 => \N__6999\,
            lcout => \beamY_RNIUBM4FZ0Z_7\,
            ltout => \beamY_RNIUBM4FZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKUC181_5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100000110"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__5707\,
            in2 => \N__4963\,
            in3 => \N__5659\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un61_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIA9P0Q_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__4937\,
            in1 => \N__4913\,
            in2 => \N__6622\,
            in3 => \N__7001\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI52RJO_5_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7000\,
            in1 => \N__5706\,
            in2 => \N__4917\,
            in3 => \N__4936\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDRE6H_3_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000011111001"
        )
    port map (
            in0 => \N__4932\,
            in1 => \N__4909\,
            in2 => \N__7667\,
            in3 => \N__7506\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un61_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICIBSR6_2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__5835\,
            in1 => \N__5814\,
            in2 => \_gnd_net_\,
            in3 => \N__8991\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIID28F1_0_3_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__5893\,
            in1 => \N__5632\,
            in2 => \N__7677\,
            in3 => \N__5688\,
            lcout => OPEN,
            ltout => \beamY_RNIID28F1_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHMJMF3_3_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5661\,
            in2 => \N__5041\,
            in3 => \N__5026\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI4AB1_5_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__5139\,
            in1 => \N__5178\,
            in2 => \N__6912\,
            in3 => \N__5038\,
            lcout => un13_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNII5M_9_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5101\,
            in1 => \N__6903\,
            in2 => \N__5074\,
            in3 => \N__5138\,
            lcout => OPEN,
            ltout => \un18_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_5_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5037\,
            in2 => \N__5029\,
            in3 => \N__5177\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIID28F1_3_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__5689\,
            in1 => \N__7668\,
            in2 => \N__5637\,
            in3 => \N__5892\,
            lcout => \beamY_RNIID28F1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5020\,
            in2 => \_gnd_net_\,
            in3 => \N__10649\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10650\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5018\,
            in3 => \N__4984\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5275\,
            in3 => \N__5251\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9075\,
            in2 => \N__5248\,
            in3 => \N__5221\,
            lcout => un1_visiblex_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5218\,
            in3 => \N__5188\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5184\,
            in3 => \N__5146\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9076\,
            in2 => \N__5143\,
            in3 => \N__5110\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6902\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9053\,
            in2 => \N__5104\,
            in3 => \N__5077\,
            lcout => \un5_visiblex_cry_7_c_RNIVZ0Z952\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5062\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHS3_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5970\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBT9_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5305\,
            in3 => \N__5944\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9539\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_67_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9540\,
            in1 => \N__6263\,
            in2 => \N__10934\,
            in3 => \N__6191\,
            lcout => g0_0_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6254\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6186\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOV5_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5296\,
            in3 => \N__5287\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQ06_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9035\,
            in2 => \N__5341\,
            in3 => \N__5284\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9544\,
            in2 => \_gnd_net_\,
            in3 => \N__5281\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5278\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9546\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9563\,
            in3 => \_gnd_net_\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9545\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6196\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5332\,
            in2 => \_gnd_net_\,
            in3 => \N__5326\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5323\,
            in2 => \N__9052\,
            in3 => \N__5317\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9565\,
            in2 => \_gnd_net_\,
            in3 => \N__5314\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5311\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5308\,
            in3 => \_gnd_net_\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5404\,
            in2 => \N__6151\,
            in3 => \N__5398\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5358\,
            in2 => \N__5395\,
            in3 => \N__5386\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6324\,
            in1 => \N__5347\,
            in2 => \N__5383\,
            in3 => \N__5374\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5371\,
            in1 => \N__5359\,
            in2 => \N__9579\,
            in3 => \N__5365\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5362\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5357\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIM4P7_0_2_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__8888\,
            in1 => \N__7931\,
            in2 => \N__8827\,
            in3 => \N__5487\,
            lcout => OPEN,
            ltout => \beamY_fast_RNIM4P7_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIO71D_3_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8807\,
            in2 => \N__5506\,
            in3 => \N__5450\,
            lcout => \beamY_fast_RNIO71DZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIM4P7_2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110100101"
        )
    port map (
            in0 => \N__8886\,
            in1 => \N__7930\,
            in2 => \N__8826\,
            in3 => \N__5486\,
            lcout => OPEN,
            ltout => \beamY_fast_RNIM4P7Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIJP9E_3_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__8808\,
            in1 => \N__8887\,
            in2 => \N__5455\,
            in3 => \N__5449\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8340\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6727\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9A1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5599\,
            in2 => \N__9109\,
            in3 => \N__5416\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAA1_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6680\,
            in2 => \N__9110\,
            in3 => \N__5413\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5410\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5407\,
            in3 => \N__6558\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9KEQ_8_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6472\,
            in1 => \N__5614\,
            in2 => \_gnd_net_\,
            in3 => \N__7853\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIK0NV_9_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7786\,
            in1 => \N__6798\,
            in2 => \_gnd_net_\,
            in3 => \N__5608\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIK0NV_0_9_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5602\,
            in3 => \_gnd_net_\,
            lcout => \beamY_RNIK0NV_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIPE7D_6_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6820\,
            in1 => \N__7854\,
            in2 => \N__6493\,
            in3 => \N__6762\,
            lcout => OPEN,
            ltout => \un5_visibley_c7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUUSO1_9_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101000"
        )
    port map (
            in0 => \N__6729\,
            in1 => \N__5593\,
            in2 => \N__5587\,
            in3 => \N__7787\,
            lcout => \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_9_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5584\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9820\,
            ce => \N__8250\,
            sr => \_gnd_net_\
        );

    \beamY_fast_7_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8153\,
            in2 => \_gnd_net_\,
            in3 => \N__5566\,
            lcout => \beamY_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9820\,
            ce => \N__8250\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5548\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9820\,
            ce => \N__8250\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI1QVS_9_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011110001111"
        )
    port map (
            in0 => \N__7855\,
            in1 => \N__5530\,
            in2 => \N__5521\,
            in3 => \N__8764\,
            lcout => \beamY_fast_RNI1QVSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9N7M7_5_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8412\,
            in1 => \N__7027\,
            in2 => \N__7003\,
            in3 => \N__7520\,
            lcout => \beamY_RNI9N7M7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2GUN3_1_9_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010110101110"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__8409\,
            in2 => \N__8476\,
            in3 => \N__8324\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un47_sum_c5,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI3M5H7_0_3_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__8410\,
            in1 => \_gnd_net_\,
            in2 => \N__5743\,
            in3 => \N__7026\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0RA9O_5_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000111100"
        )
    port map (
            in0 => \N__7519\,
            in1 => \N__6967\,
            in2 => \N__5722\,
            in3 => \N__6637\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRRO4H1_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101100000000"
        )
    port map (
            in0 => \N__6638\,
            in1 => \N__7666\,
            in2 => \N__5719\,
            in3 => \N__5716\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKUC181_0_5_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__5633\,
            in1 => \N__5697\,
            in2 => \_gnd_net_\,
            in3 => \N__5667\,
            lcout => \beamY_RNIKUC181_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI779U3_5_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8411\,
            in1 => \N__7025\,
            in2 => \_gnd_net_\,
            in3 => \N__7518\,
            lcout => \beamY_RNI779U3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKPNA02_5_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000101111110"
        )
    port map (
            in0 => \N__5698\,
            in1 => \N__5668\,
            in2 => \N__5638\,
            in3 => \N__5894\,
            lcout => \beamY_RNIKPNA02Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5AJJ02_3_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__5918\,
            in1 => \N__5896\,
            in2 => \N__7678\,
            in3 => \N__7522\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5F8A81_3_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__7521\,
            in1 => \N__7672\,
            in2 => \_gnd_net_\,
            in3 => \N__5917\,
            lcout => OPEN,
            ltout => \beamY_RNI5F8A81Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7VNCG5_3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__8103\,
            in1 => \N__5844\,
            in2 => \N__5899\,
            in3 => \N__5895\,
            lcout => OPEN,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIAJLT9A_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__5872\,
            in1 => \N__5853\,
            in2 => \N__5866\,
            in3 => \N__5863\,
            lcout => \beamY_RNIAJLT9AZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1UL7G5_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__7673\,
            in1 => \N__8104\,
            in2 => \N__5857\,
            in3 => \N__5845\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un68_sum_c4,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQBCMCE_3_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__5790\,
            in1 => \N__5836\,
            in2 => \N__5824\,
            in3 => \N__5821\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISDALMO_2_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__5803\,
            in1 => \N__5797\,
            in2 => \N__5791\,
            in3 => \N__6853\,
            lcout => font_un42_pixel_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9718\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5982\,
            in2 => \N__5779\,
            in3 => \N__5764\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_60_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7213\,
            in2 => \N__7111\,
            in3 => \N__5761\,
            lcout => \Pixel_1_esr_RNOZ0Z_60\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7212\,
            in1 => \N__5983\,
            in2 => \N__7252\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOC_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7237\,
            in2 => \_gnd_net_\,
            in3 => \N__5974\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIO1J8_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6262\,
            in1 => \N__6193\,
            in2 => \N__10933\,
            in3 => \N__9562\,
            lcout => \G_25_i_o8_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_21_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__9719\,
            in2 => \_gnd_net_\,
            in3 => \N__9639\,
            lcout => \G_25_i_a8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_65_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6261\,
            in1 => \N__6192\,
            in2 => \N__10932\,
            in3 => \N__9561\,
            lcout => g0_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNISG94_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6252\,
            in2 => \_gnd_net_\,
            in3 => \N__6194\,
            lcout => un22_visibley_2,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2G_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5971\,
            in2 => \N__6147\,
            in3 => \N__5959\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJ_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6060\,
            in2 => \N__5956\,
            in3 => \N__5947\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI273E1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__5943\,
            in2 => \N__5932\,
            in3 => \N__5923\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6067\,
            in1 => \N__6061\,
            in2 => \N__9564\,
            in3 => \N__6052\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6049\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_8_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6046\,
            in1 => \N__6253\,
            in2 => \_gnd_net_\,
            in3 => \N__6195\,
            lcout => g0_i_o4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_20_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9726\,
            in1 => \N__11105\,
            in2 => \N__10548\,
            in3 => \N__10847\,
            lcout => un22_visibleylt9_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10941\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEM_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6040\,
            in2 => \N__6000\,
            in3 => \N__6034\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICND41_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6031\,
            in2 => \N__6019\,
            in3 => \N__6010\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNI9KOM2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6126\,
            in1 => \N__6007\,
            in2 => \N__6001\,
            in3 => \N__5986\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6208\,
            in2 => \_gnd_net_\,
            in3 => \N__6202\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6199\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6187\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIK454_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__10925\,
            in1 => \N__9640\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un22_visibley_3,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9J1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6334\,
            in2 => \N__6096\,
            in3 => \N__6130\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAM72_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6127\,
            in2 => \N__6115\,
            in3 => \N__6106\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI53BF5_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7182\,
            in1 => \N__6103\,
            in2 => \N__6097\,
            in3 => \N__6082\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6079\,
            in2 => \_gnd_net_\,
            in3 => \N__6073\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6070\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9641\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10924\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10942\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6300\,
            in2 => \N__6217\,
            in3 => \N__6328\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6325\,
            in2 => \N__6313\,
            in3 => \N__6304\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI31V25_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7322\,
            in1 => \N__6301\,
            in2 => \N__6292\,
            in3 => \N__6283\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6280\,
            in2 => \_gnd_net_\,
            in3 => \N__6274\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6271\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7516\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6419\,
            in2 => \N__6361\,
            in3 => \N__6376\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6343\,
            in2 => \N__6424\,
            in3 => \N__6373\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58S32_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6423\,
            in2 => \N__6460\,
            in3 => \N__6370\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNISMP75_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7420\,
            in1 => \N__6400\,
            in2 => \N__6448\,
            in3 => \N__6367\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6436\,
            in2 => \_gnd_net_\,
            in3 => \N__6364\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8377\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_3_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8034\,
            in1 => \N__8969\,
            in2 => \_gnd_net_\,
            in3 => \N__7958\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8402\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6514\,
            in2 => \N__6352\,
            in3 => \N__6337\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48A1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6385\,
            in2 => \N__6520\,
            in3 => \N__6451\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5Q1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6518\,
            in2 => \N__6589\,
            in3 => \N__6439\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIGK8A2_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6418\,
            in1 => \N__6499\,
            in2 => \N__6571\,
            in3 => \N__6430\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6538\,
            in1 => \N__6519\,
            in2 => \N__6559\,
            in3 => \N__6427\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6403\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9KEQ_0_8_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_RNI9KEQ_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8341\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8R_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9102\,
            in2 => \N__6394\,
            in3 => \N__6379\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555B1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6595\,
            in2 => \N__9111\,
            in3 => \N__6580\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797B1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6577\,
            in2 => \N__9112\,
            in3 => \N__6562\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6554\,
            in2 => \_gnd_net_\,
            in3 => \N__6532\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6529\,
            in2 => \_gnd_net_\,
            in3 => \N__6523\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6502\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIRPUB_6_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6489\,
            in1 => \N__6819\,
            in2 => \_gnd_net_\,
            in3 => \N__6758\,
            lcout => un5_visibley_c6_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_0_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000000100"
        )
    port map (
            in0 => \N__8048\,
            in1 => \N__8914\,
            in2 => \N__7966\,
            in3 => \N__8996\,
            lcout => OPEN,
            ltout => \un11_visibleylto9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIICI12_5_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8415\,
            in1 => \N__8339\,
            in2 => \N__6466\,
            in3 => \N__6735\,
            lcout => OPEN,
            ltout => \un11_visibleylto9_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6D913_9_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6463\,
            in3 => \N__6689\,
            lcout => un11_visibley,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_6_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6838\,
            lcout => \beamY_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__8229\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIH5V7_6_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6818\,
            in2 => \_gnd_net_\,
            in3 => \N__6757\,
            lcout => un5_visibley_c6_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_5_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6787\,
            lcout => \beamY_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9823\,
            ce => \N__8229\,
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0DB_9_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6961\,
            in1 => \N__7800\,
            in2 => \N__6610\,
            in3 => \N__7868\,
            lcout => \beamY_RNIJ0DBZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIECTA3_8_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010000111"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__6736\,
            in2 => \N__8470\,
            in3 => \N__6690\,
            lcout => \beamY_RNIECTA3Z0Z_8\,
            ltout => \beamY_RNIECTA3Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI3M5H7_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__8414\,
            in1 => \N__6995\,
            in2 => \N__6649\,
            in3 => \_gnd_net_\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICE7B5_4_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__6601\,
            in1 => \N__7024\,
            in2 => \_gnd_net_\,
            in3 => \N__7959\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_1_5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__9004\,
            in2 => \N__10345\,
            in3 => \N__8921\,
            lcout => un1_beamylto9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI4H1V1_0_9_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__8344\,
            in1 => \N__8465\,
            in2 => \_gnd_net_\,
            in3 => \N__8413\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0,
            ltout => \font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIKDT19_9_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101101001"
        )
    port map (
            in0 => \N__7023\,
            in1 => \N__6994\,
            in2 => \N__6970\,
            in3 => \_gnd_net_\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGKP3_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8065\,
            in1 => \N__8767\,
            in2 => \_gnd_net_\,
            in3 => \N__7960\,
            lcout => un1_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_46_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010100010"
        )
    port map (
            in0 => \N__6946\,
            in1 => \N__9754\,
            in2 => \N__10849\,
            in3 => \N__6955\,
            lcout => un27lt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_45_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110110100010"
        )
    port map (
            in0 => \N__6954\,
            in1 => \N__6945\,
            in2 => \N__9763\,
            in3 => \N__6937\,
            lcout => un1_visiblex_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_52_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__6872\,
            in1 => \N__6855\,
            in2 => \_gnd_net_\,
            in3 => \N__9007\,
            lcout => OPEN,
            ltout => \g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_29_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__10356\,
            in1 => \N__10034\,
            in2 => \N__6931\,
            in3 => \N__8060\,
            lcout => g1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI34L6_10_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8636\,
            in1 => \N__8584\,
            in2 => \N__6928\,
            in3 => \N__6916\,
            lcout => un1_beamx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILTIMMO_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010100101"
        )
    port map (
            in0 => \N__8059\,
            in1 => \N__6854\,
            in2 => \N__6874\,
            in3 => \N__9005\,
            lcout => font_un78_pixellto3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_50_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111010110001"
        )
    port map (
            in0 => \N__9006\,
            in1 => \N__6873\,
            in2 => \N__6859\,
            in3 => \N__8061\,
            lcout => g1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__10543\,
            in1 => \N__10722\,
            in2 => \_gnd_net_\,
            in3 => \N__10429\,
            lcout => OPEN,
            ltout => \r_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI6J1NH2_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110001001100"
        )
    port map (
            in0 => \N__10681\,
            in1 => \N__8544\,
            in2 => \N__7096\,
            in3 => \N__9121\,
            lcout => \Pixel_3_sqmuxa_1_1\,
            ltout => \Pixel_3_sqmuxa_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEC74VJ1_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001100000"
        )
    port map (
            in0 => \N__10358\,
            in1 => \N__7093\,
            in2 => \N__7087\,
            in3 => \N__10033\,
            lcout => \Pixel_7_sqmuxa_1\,
            ltout => \Pixel_7_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_9_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__7084\,
            in1 => \N__7131\,
            in2 => \N__7075\,
            in3 => \N__8512\,
            lcout => \G_25_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_28_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001000"
        )
    port map (
            in0 => \N__10544\,
            in1 => \N__10723\,
            in2 => \N__7072\,
            in3 => \N__10430\,
            lcout => OPEN,
            ltout => \g0_0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_11_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7057\,
            in1 => \N__7048\,
            in2 => \N__7051\,
            in3 => \N__7036\,
            lcout => \G_25_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_27_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011001"
        )
    port map (
            in0 => \N__10217\,
            in1 => \N__10357\,
            in2 => \_gnd_net_\,
            in3 => \N__10032\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_49_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7042\,
            in1 => \N__7159\,
            in2 => \_gnd_net_\,
            in3 => \N__7035\,
            lcout => g0_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_4_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__7120\,
            in1 => \N__7279\,
            in2 => \N__7582\,
            in3 => \N__7294\,
            lcout => \Pixel_9_u_ns_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11103\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_35_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111011111"
        )
    port map (
            in0 => \N__10563\,
            in1 => \N__10359\,
            in2 => \N__10219\,
            in3 => \N__10442\,
            lcout => g1_0_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_15_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__10443\,
            in1 => \N__10363\,
            in2 => \_gnd_net_\,
            in3 => \N__10564\,
            lcout => g1_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_24_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__10677\,
            in1 => \N__10726\,
            in2 => \N__10578\,
            in3 => \N__10444\,
            lcout => \G_25_i_a8_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_17_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__10218\,
            in1 => \N__10076\,
            in2 => \_gnd_net_\,
            in3 => \N__10676\,
            lcout => g2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_64_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001110"
        )
    port map (
            in0 => \N__10846\,
            in1 => \N__9762\,
            in2 => \N__9139\,
            in3 => \N__9657\,
            lcout => \N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_12_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7150\,
            in1 => \N__9268\,
            in2 => \N__7138\,
            in3 => \N__7119\,
            lcout => \N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9655\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7300\,
            in2 => \N__10861\,
            in3 => \N__7099\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7327\,
            in2 => \N__7264\,
            in3 => \N__7240\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIP79LC_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7211\,
            in1 => \N__7333\,
            in2 => \N__7351\,
            in3 => \N__7228\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109G5_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7225\,
            in2 => \_gnd_net_\,
            in3 => \N__7216\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_56_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__10843\,
            in2 => \_gnd_net_\,
            in3 => \N__9758\,
            lcout => un28_visibleylt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_37_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__10675\,
            in1 => \N__10571\,
            in2 => \_gnd_net_\,
            in3 => \N__10445\,
            lcout => OPEN,
            ltout => \g0_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_16_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__10074\,
            in1 => \N__10192\,
            in2 => \N__7195\,
            in3 => \N__10368\,
            lcout => g1_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9752\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17M43_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7192\,
            in2 => \N__7380\,
            in3 => \N__7186\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VL4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7183\,
            in2 => \N__7171\,
            in3 => \N__7162\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNICOQ2B_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9390\,
            in1 => \N__7387\,
            in2 => \N__7381\,
            in3 => \N__7366\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7363\,
            in2 => \_gnd_net_\,
            in3 => \N__7357\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7354\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KK4_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__7347\,
            in1 => \_gnd_net_\,
            in2 => \N__7326\,
            in3 => \_gnd_net_\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7318\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_13_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111000101"
        )
    port map (
            in0 => \N__7588\,
            in1 => \N__7275\,
            in2 => \N__7531\,
            in3 => \N__7572\,
            lcout => \Pixel_9_sn_N_7_mux_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIVFV5_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__10844\,
            in1 => \N__9760\,
            in2 => \_gnd_net_\,
            in3 => \N__11106\,
            lcout => OPEN,
            ltout => \un16_visibleylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNISDFC_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7550\,
            in2 => \N__7282\,
            in3 => \N__9580\,
            lcout => un16_visibley_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_33_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7597\,
            in1 => \N__10944\,
            in2 => \N__9586\,
            in3 => \N__7551\,
            lcout => \Pixel_7_sqmuxa_3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_55_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9761\,
            in1 => \N__11107\,
            in2 => \N__10579\,
            in3 => \N__10845\,
            lcout => OPEN,
            ltout => \un22_visibleylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_32_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__9584\,
            in1 => \N__7571\,
            in2 => \N__7555\,
            in3 => \N__7552\,
            lcout => un22_visibley,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7517\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7419\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7622\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51F3_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7421\,
            in2 => \N__7447\,
            in3 => \N__7438\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNU3_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7435\,
            in2 => \N__7426\,
            in3 => \N__7429\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKE4_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7425\,
            in2 => \N__7399\,
            in3 => \N__7390\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIC4FVA_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8505\,
            in1 => \N__7750\,
            in2 => \N__7744\,
            in3 => \N__7735\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7732\,
            in2 => \_gnd_net_\,
            in3 => \N__7726\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8092\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6V5_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8500\,
            in2 => \N__7606\,
            in3 => \N__7723\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINI399_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7720\,
            in2 => \N__8506\,
            in3 => \N__7714\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BRO9_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8504\,
            in2 => \N__7711\,
            in3 => \N__7702\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAPMAL_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9443\,
            in1 => \N__8482\,
            in2 => \N__7699\,
            in3 => \N__7690\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1B_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7687\,
            in2 => \_gnd_net_\,
            in3 => \N__7681\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7635\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8499\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI4H1V1_9_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__8475\,
            in1 => \N__8416\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => font_un42_pixel_if_generate_plus_mult1_un47_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2ROB_9_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__7965\,
            in1 => \N__7801\,
            in2 => \N__8269\,
            in3 => \N__7870\,
            lcout => un8_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001111000"
        )
    port map (
            in0 => \N__8254\,
            in1 => \N__10213\,
            in2 => \N__10346\,
            in3 => \N__8158\,
            lcout => un28lto1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8102\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8995\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8047\,
            lcout => un4_beamylt6,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_5_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8842\,
            in1 => \N__8922\,
            in2 => \N__7969\,
            in3 => \N__7961\,
            lcout => OPEN,
            ltout => \un4_beamylt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_9_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__7880\,
            in1 => \N__8765\,
            in2 => \N__7813\,
            in3 => \N__7809\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__9923\,
            in1 => \N__9095\,
            in2 => \_gnd_net_\,
            in3 => \N__8994\,
            lcout => \beamY_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMJIF_7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8923\,
            in1 => \N__8854\,
            in2 => \N__8848\,
            in3 => \N__8766\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110000"
        )
    port map (
            in0 => \N__8560\,
            in1 => \N__8583\,
            in2 => \N__8698\,
            in3 => \N__8590\,
            lcout => OPEN,
            ltout => \Pixel_1_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8701\,
            in3 => \N__9875\,
            lcout => \Pixel_1_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNINAS01_10_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8653\,
            in1 => \N__8647\,
            in2 => \N__8638\,
            in3 => \N__8596\,
            lcout => un15_beamy_2,
            ltout => \un15_beamy_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_44_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__8582\,
            in1 => \N__8559\,
            in2 => \N__8548\,
            in3 => \N__8545\,
            lcout => OPEN,
            ltout => \Pixel_9_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_22_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000010000"
        )
    port map (
            in0 => \N__8527\,
            in1 => \N__8521\,
            in2 => \N__8515\,
            in3 => \N__9949\,
            lcout => \Pixel_9_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \N__9244\,
            in2 => \N__9280\,
            in3 => \N__10585\,
            lcout => OPEN,
            ltout => \N_163_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9232\,
            in2 => \N__9226\,
            in3 => \N__9145\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9816\,
            ce => \N__9193\,
            sr => \N__9889\
        );

    \Pixel_1_esr_RNO_26_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011000000000"
        )
    port map (
            in0 => \N__9187\,
            in1 => \N__10070\,
            in2 => \N__10355\,
            in3 => \N__9181\,
            lcout => OPEN,
            ltout => \g0_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_10_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__9253\,
            in1 => \N__9175\,
            in2 => \N__9169\,
            in3 => \N__10741\,
            lcout => OPEN,
            ltout => \G_25_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9166\,
            in1 => \N__9160\,
            in2 => \N__9154\,
            in3 => \N__9151\,
            lcout => \Pixel_9_u_ns_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_69_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10549\,
            in2 => \_gnd_net_\,
            in3 => \N__11104\,
            lcout => g2_1,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OT9_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9130\,
            in2 => \N__9330\,
            in3 => \N__9124\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JF21_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11041\,
            in2 => \N__10963\,
            in3 => \N__9115\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11011\,
            in2 => \N__9331\,
            in3 => \N__10958\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QB1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__9316\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_34_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111101010000"
        )
    port map (
            in0 => \N__10550\,
            in1 => \_gnd_net_\,
            in2 => \N__9313\,
            in3 => \N__10727\,
            lcout => OPEN,
            ltout => \font_un19_pixel_0_0_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_14_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__10075\,
            in1 => \N__9310\,
            in2 => \N__9304\,
            in3 => \N__9400\,
            lcout => OPEN,
            ltout => \font_un237_pixel_6_ns_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_5_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__9301\,
            in1 => \N__9295\,
            in2 => \N__9289\,
            in3 => \N__9286\,
            lcout => font_un237_pixel_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_54_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011101101"
        )
    port map (
            in0 => \N__10574\,
            in1 => \N__9262\,
            in2 => \N__10446\,
            in3 => \N__10682\,
            lcout => OPEN,
            ltout => \g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_31_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__10214\,
            in1 => \N__10350\,
            in2 => \N__9271\,
            in3 => \N__10073\,
            lcout => font_un83_pixel_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10573\,
            in2 => \N__10729\,
            in3 => \N__10422\,
            lcout => font_un19_pixel_23,
            ltout => \font_un19_pixel_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_25_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101100100"
        )
    port map (
            in0 => \N__10072\,
            in1 => \N__10215\,
            in2 => \N__9256\,
            in3 => \N__10354\,
            lcout => font_un160_pixel_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_57_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100001001000"
        )
    port map (
            in0 => \N__10575\,
            in1 => \N__10683\,
            in2 => \N__10447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_36_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001010000"
        )
    port map (
            in0 => \N__10216\,
            in1 => \N__10351\,
            in2 => \N__9403\,
            in3 => \N__10071\,
            lcout => g3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10836\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4M96_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9667\,
            in2 => \N__9360\,
            in3 => \N__9394\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCC9_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9391\,
            in2 => \N__9379\,
            in3 => \N__9370\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNISKRFM_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11031\,
            in1 => \N__9367\,
            in2 => \N__9361\,
            in3 => \N__9346\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9343\,
            in2 => \_gnd_net_\,
            in3 => \N__9337\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0\,
            ltout => \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9334\,
            in3 => \_gnd_net_\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9753\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_7_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9661\,
            in1 => \N__10945\,
            in2 => \_gnd_net_\,
            in3 => \N__9585\,
            lcout => g0_i_o4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9924\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEB_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9484\,
            in2 => \N__9444\,
            in3 => \N__9478\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9H_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9439\,
            in2 => \N__9475\,
            in3 => \N__9466\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_62_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9463\,
            in2 => \N__9445\,
            in3 => \N__9457\,
            lcout => \Pixel_1_esr_RNOZ0Z_62\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9418\,
            in2 => \N__9454\,
            in3 => \N__9435\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJL_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9412\,
            in2 => \_gnd_net_\,
            in3 => \N__9406\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_68_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010001000"
        )
    port map (
            in0 => \N__9933\,
            in1 => \N__9942\,
            in2 => \N__9925\,
            in3 => \N__9959\,
            lcout => OPEN,
            ltout => \un28lto4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_63_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__9960\,
            in1 => \N__10261\,
            in2 => \N__9973\,
            in3 => \N__9922\,
            lcout => OPEN,
            ltout => \un28lt10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_47_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000101"
        )
    port map (
            in0 => \N__9970\,
            in1 => \N__9895\,
            in2 => \N__9964\,
            in3 => \N__9961\,
            lcout => un28_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_61_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__9943\,
            in1 => \N__9934\,
            in2 => \_gnd_net_\,
            in3 => \N__9921\,
            lcout => \un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9888\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_39_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__10305\,
            in1 => \N__10191\,
            in2 => \_gnd_net_\,
            in3 => \N__10046\,
            lcout => \Pixel_1_esr_RNOZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_58_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__10546\,
            in1 => \_gnd_net_\,
            in2 => \N__10448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_38_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010101111"
        )
    port map (
            in0 => \N__10209\,
            in1 => \N__10319\,
            in2 => \N__9775\,
            in3 => \N__10063\,
            lcout => OPEN,
            ltout => \N_1304_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_18_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010111000"
        )
    port map (
            in0 => \N__9772\,
            in1 => \N__10750\,
            in2 => \N__9766\,
            in3 => \N__10725\,
            lcout => \N_156_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_40_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10545\,
            in2 => \_gnd_net_\,
            in3 => \N__10431\,
            lcout => g1_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_48_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001010"
        )
    port map (
            in0 => \N__10547\,
            in1 => \_gnd_net_\,
            in2 => \N__10449\,
            in3 => \N__10724\,
            lcout => OPEN,
            ltout => \N_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_23_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__10210\,
            in1 => \N__10320\,
            in2 => \N__10744\,
            in3 => \N__10064\,
            lcout => \G_25_i_a8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_59_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__10577\,
            in1 => \_gnd_net_\,
            in2 => \N__10450\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \g1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_41_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011101111110"
        )
    port map (
            in0 => \N__10078\,
            in1 => \N__10212\,
            in2 => \N__10735\,
            in3 => \N__10353\,
            lcout => OPEN,
            ltout => \N_1302_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_19_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010111000"
        )
    port map (
            in0 => \N__9979\,
            in1 => \N__10375\,
            in2 => \N__10732\,
            in3 => \N__10728\,
            lcout => OPEN,
            ltout => \N_159_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_6_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10684\,
            in2 => \N__10594\,
            in3 => \N__10591\,
            lcout => font_un314_pixel_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_43_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10576\,
            in2 => \_gnd_net_\,
            in3 => \N__10438\,
            lcout => g1_3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_esr_RNO_42_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__10352\,
            in1 => \N__10211\,
            in2 => \_gnd_net_\,
            in3 => \N__10077\,
            lcout => \N_1303_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11095\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLB_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10756\,
            in2 => \N__10995\,
            in3 => \N__11035\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTH_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11032\,
            in2 => \N__11020\,
            in3 => \N__11005\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0\,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI102IB1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10962\,
            in1 => \N__11002\,
            in2 => \N__10996\,
            in3 => \N__10975\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHM_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10972\,
            in2 => \_gnd_net_\,
            in3 => \N__10966\,
            lcout => \font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10943\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10848\,
            lcout => font_un19_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
