// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 24 2015 19:04:50

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSync,
    SCLK1,
    Pixel,
    HSync,
    nCS2,
    SDATA2,
    SCLK2,
    Clock12MHz,
    nCS1,
    SDATA1);

    output VSync;
    output SCLK1;
    output Pixel;
    output HSync;
    output nCS2;
    output SDATA2;
    output SCLK2;
    input Clock12MHz;
    output nCS1;
    input SDATA1;

    wire N__26093;
    wire N__26092;
    wire N__26091;
    wire N__26082;
    wire N__26081;
    wire N__26080;
    wire N__26073;
    wire N__26072;
    wire N__26071;
    wire N__26064;
    wire N__26063;
    wire N__26062;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26046;
    wire N__26045;
    wire N__26044;
    wire N__26037;
    wire N__26036;
    wire N__26035;
    wire N__26028;
    wire N__26027;
    wire N__26026;
    wire N__26019;
    wire N__26018;
    wire N__26017;
    wire N__26010;
    wire N__26009;
    wire N__26008;
    wire N__25991;
    wire N__25990;
    wire N__25989;
    wire N__25988;
    wire N__25987;
    wire N__25986;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25976;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25968;
    wire N__25967;
    wire N__25966;
    wire N__25963;
    wire N__25962;
    wire N__25961;
    wire N__25960;
    wire N__25959;
    wire N__25958;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25937;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25921;
    wire N__25918;
    wire N__25907;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25875;
    wire N__25872;
    wire N__25871;
    wire N__25870;
    wire N__25869;
    wire N__25862;
    wire N__25855;
    wire N__25852;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25823;
    wire N__25820;
    wire N__25819;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25807;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25739;
    wire N__25738;
    wire N__25737;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25715;
    wire N__25710;
    wire N__25709;
    wire N__25708;
    wire N__25705;
    wire N__25694;
    wire N__25693;
    wire N__25692;
    wire N__25691;
    wire N__25690;
    wire N__25689;
    wire N__25688;
    wire N__25687;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25654;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25621;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25586;
    wire N__25585;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25542;
    wire N__25541;
    wire N__25540;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25518;
    wire N__25517;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25474;
    wire N__25463;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25432;
    wire N__25427;
    wire N__25418;
    wire N__25417;
    wire N__25416;
    wire N__25415;
    wire N__25410;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25398;
    wire N__25397;
    wire N__25396;
    wire N__25395;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25387;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25373;
    wire N__25370;
    wire N__25365;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25327;
    wire N__25322;
    wire N__25321;
    wire N__25314;
    wire N__25311;
    wire N__25310;
    wire N__25307;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25285;
    wire N__25280;
    wire N__25277;
    wire N__25268;
    wire N__25265;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25225;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25208;
    wire N__25207;
    wire N__25206;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25177;
    wire N__25168;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25150;
    wire N__25149;
    wire N__25146;
    wire N__25145;
    wire N__25142;
    wire N__25141;
    wire N__25140;
    wire N__25137;
    wire N__25136;
    wire N__25135;
    wire N__25134;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25105;
    wire N__25098;
    wire N__25095;
    wire N__25082;
    wire N__25081;
    wire N__25080;
    wire N__25079;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25074;
    wire N__25071;
    wire N__25070;
    wire N__25069;
    wire N__25068;
    wire N__25067;
    wire N__25066;
    wire N__25065;
    wire N__25064;
    wire N__25059;
    wire N__25058;
    wire N__25057;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25043;
    wire N__25042;
    wire N__25037;
    wire N__25036;
    wire N__25035;
    wire N__25032;
    wire N__25031;
    wire N__25030;
    wire N__25029;
    wire N__25028;
    wire N__25027;
    wire N__25026;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25016;
    wire N__25015;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25008;
    wire N__25007;
    wire N__25006;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24985;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24967;
    wire N__24964;
    wire N__24959;
    wire N__24954;
    wire N__24949;
    wire N__24938;
    wire N__24929;
    wire N__24920;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24904;
    wire N__24897;
    wire N__24890;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24860;
    wire N__24859;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24855;
    wire N__24854;
    wire N__24853;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24839;
    wire N__24838;
    wire N__24837;
    wire N__24836;
    wire N__24835;
    wire N__24834;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24828;
    wire N__24827;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24821;
    wire N__24818;
    wire N__24817;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24804;
    wire N__24801;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24786;
    wire N__24781;
    wire N__24778;
    wire N__24777;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24760;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24752;
    wire N__24749;
    wire N__24748;
    wire N__24743;
    wire N__24734;
    wire N__24729;
    wire N__24726;
    wire N__24725;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24707;
    wire N__24704;
    wire N__24695;
    wire N__24690;
    wire N__24683;
    wire N__24678;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24659;
    wire N__24656;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24629;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24598;
    wire N__24595;
    wire N__24594;
    wire N__24593;
    wire N__24588;
    wire N__24583;
    wire N__24580;
    wire N__24575;
    wire N__24572;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24556;
    wire N__24545;
    wire N__24544;
    wire N__24543;
    wire N__24542;
    wire N__24541;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24525;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24511;
    wire N__24510;
    wire N__24509;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24505;
    wire N__24504;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24485;
    wire N__24484;
    wire N__24483;
    wire N__24482;
    wire N__24481;
    wire N__24480;
    wire N__24479;
    wire N__24478;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24474;
    wire N__24473;
    wire N__24472;
    wire N__24471;
    wire N__24468;
    wire N__24463;
    wire N__24458;
    wire N__24451;
    wire N__24440;
    wire N__24437;
    wire N__24432;
    wire N__24425;
    wire N__24420;
    wire N__24413;
    wire N__24404;
    wire N__24393;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24349;
    wire N__24348;
    wire N__24347;
    wire N__24344;
    wire N__24333;
    wire N__24330;
    wire N__24325;
    wire N__24322;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24139;
    wire N__24138;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24100;
    wire N__24093;
    wire N__24090;
    wire N__24081;
    wire N__24078;
    wire N__24071;
    wire N__24068;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24005;
    wire N__24002;
    wire N__24001;
    wire N__24000;
    wire N__23999;
    wire N__23998;
    wire N__23995;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23987;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23971;
    wire N__23970;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23951;
    wire N__23944;
    wire N__23941;
    wire N__23936;
    wire N__23927;
    wire N__23922;
    wire N__23917;
    wire N__23908;
    wire N__23891;
    wire N__23888;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23884;
    wire N__23883;
    wire N__23882;
    wire N__23881;
    wire N__23880;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23861;
    wire N__23860;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23844;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23810;
    wire N__23807;
    wire N__23802;
    wire N__23799;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23789;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23774;
    wire N__23765;
    wire N__23760;
    wire N__23753;
    wire N__23748;
    wire N__23745;
    wire N__23736;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23609;
    wire N__23608;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23568;
    wire N__23565;
    wire N__23560;
    wire N__23555;
    wire N__23548;
    wire N__23545;
    wire N__23534;
    wire N__23531;
    wire N__23530;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23519;
    wire N__23514;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23489;
    wire N__23486;
    wire N__23479;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23443;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23435;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23426;
    wire N__23425;
    wire N__23424;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23418;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23399;
    wire N__23390;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23359;
    wire N__23354;
    wire N__23353;
    wire N__23350;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23322;
    wire N__23319;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23303;
    wire N__23302;
    wire N__23301;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23289;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23281;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23265;
    wire N__23264;
    wire N__23261;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23244;
    wire N__23243;
    wire N__23236;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23226;
    wire N__23217;
    wire N__23214;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23192;
    wire N__23185;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23081;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23054;
    wire N__23051;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23032;
    wire N__23031;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23020;
    wire N__23019;
    wire N__23018;
    wire N__23017;
    wire N__23016;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22987;
    wire N__22986;
    wire N__22985;
    wire N__22984;
    wire N__22979;
    wire N__22970;
    wire N__22965;
    wire N__22962;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22940;
    wire N__22935;
    wire N__22930;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22793;
    wire N__22792;
    wire N__22789;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22777;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22769;
    wire N__22766;
    wire N__22761;
    wire N__22758;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22744;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22736;
    wire N__22733;
    wire N__22732;
    wire N__22731;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22717;
    wire N__22712;
    wire N__22709;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22665;
    wire N__22664;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22611;
    wire N__22608;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22582;
    wire N__22577;
    wire N__22574;
    wire N__22569;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22525;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22492;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22477;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22462;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22413;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22314;
    wire N__22311;
    wire N__22310;
    wire N__22309;
    wire N__22306;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22246;
    wire N__22243;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22192;
    wire N__22189;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22171;
    wire N__22168;
    wire N__22163;
    wire N__22162;
    wire N__22159;
    wire N__22158;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22147;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22137;
    wire N__22132;
    wire N__22127;
    wire N__22120;
    wire N__22117;
    wire N__22112;
    wire N__22107;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22093;
    wire N__22092;
    wire N__22089;
    wire N__22088;
    wire N__22087;
    wire N__22086;
    wire N__22085;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22076;
    wire N__22075;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22068;
    wire N__22067;
    wire N__22060;
    wire N__22057;
    wire N__22048;
    wire N__22045;
    wire N__22036;
    wire N__22033;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22025;
    wire N__22024;
    wire N__22023;
    wire N__22022;
    wire N__22021;
    wire N__22020;
    wire N__22013;
    wire N__22006;
    wire N__22005;
    wire N__22004;
    wire N__22003;
    wire N__22000;
    wire N__21995;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21968;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21909;
    wire N__21908;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21900;
    wire N__21893;
    wire N__21892;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21871;
    wire N__21870;
    wire N__21867;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21852;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21833;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21789;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21742;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21625;
    wire N__21624;
    wire N__21623;
    wire N__21620;
    wire N__21615;
    wire N__21612;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21510;
    wire N__21503;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21425;
    wire N__21422;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21317;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21259;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21163;
    wire N__21160;
    wire N__21159;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21141;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21053;
    wire N__21052;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20970;
    wire N__20967;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20939;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20930;
    wire N__20925;
    wire N__20924;
    wire N__20921;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20893;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20887;
    wire N__20886;
    wire N__20885;
    wire N__20884;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20866;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20858;
    wire N__20855;
    wire N__20850;
    wire N__20847;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20791;
    wire N__20790;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20712;
    wire N__20693;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20648;
    wire N__20641;
    wire N__20638;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20603;
    wire N__20602;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20473;
    wire N__20468;
    wire N__20465;
    wire N__20464;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20350;
    wire N__20349;
    wire N__20348;
    wire N__20345;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20321;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20279;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20218;
    wire N__20217;
    wire N__20216;
    wire N__20211;
    wire N__20210;
    wire N__20209;
    wire N__20208;
    wire N__20207;
    wire N__20206;
    wire N__20205;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20199;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20178;
    wire N__20175;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20150;
    wire N__20145;
    wire N__20142;
    wire N__20137;
    wire N__20132;
    wire N__20125;
    wire N__20122;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20104;
    wire N__20099;
    wire N__20096;
    wire N__20091;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20058;
    wire N__20057;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19997;
    wire N__19994;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19982;
    wire N__19981;
    wire N__19980;
    wire N__19979;
    wire N__19978;
    wire N__19977;
    wire N__19976;
    wire N__19975;
    wire N__19974;
    wire N__19973;
    wire N__19972;
    wire N__19971;
    wire N__19970;
    wire N__19969;
    wire N__19968;
    wire N__19967;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19960;
    wire N__19957;
    wire N__19956;
    wire N__19955;
    wire N__19954;
    wire N__19953;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19819;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19753;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19717;
    wire N__19716;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19698;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19681;
    wire N__19678;
    wire N__19677;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19600;
    wire N__19599;
    wire N__19598;
    wire N__19595;
    wire N__19590;
    wire N__19587;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19511;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19451;
    wire N__19450;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19433;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19419;
    wire N__19418;
    wire N__19413;
    wire N__19412;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19369;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19352;
    wire N__19349;
    wire N__19344;
    wire N__19341;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19322;
    wire N__19321;
    wire N__19320;
    wire N__19319;
    wire N__19318;
    wire N__19315;
    wire N__19310;
    wire N__19309;
    wire N__19308;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19304;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19300;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19292;
    wire N__19291;
    wire N__19290;
    wire N__19289;
    wire N__19288;
    wire N__19285;
    wire N__19284;
    wire N__19281;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19265;
    wire N__19262;
    wire N__19257;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19243;
    wire N__19234;
    wire N__19229;
    wire N__19226;
    wire N__19221;
    wire N__19218;
    wire N__19213;
    wire N__19210;
    wire N__19203;
    wire N__19198;
    wire N__19187;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19167;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19135;
    wire N__19132;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19114;
    wire N__19113;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__19107;
    wire N__19102;
    wire N__19093;
    wire N__19086;
    wire N__19081;
    wire N__19074;
    wire N__19071;
    wire N__19066;
    wire N__19063;
    wire N__19052;
    wire N__19051;
    wire N__19048;
    wire N__19047;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19010;
    wire N__19005;
    wire N__18998;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18974;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18944;
    wire N__18941;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18726;
    wire N__18725;
    wire N__18724;
    wire N__18721;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18704;
    wire N__18701;
    wire N__18700;
    wire N__18699;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18687;
    wire N__18684;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18638;
    wire N__18637;
    wire N__18632;
    wire N__18629;
    wire N__18628;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18615;
    wire N__18614;
    wire N__18613;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18577;
    wire N__18572;
    wire N__18569;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18551;
    wire N__18548;
    wire N__18547;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18542;
    wire N__18541;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18505;
    wire N__18504;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18482;
    wire N__18481;
    wire N__18480;
    wire N__18479;
    wire N__18478;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18434;
    wire N__18431;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18402;
    wire N__18399;
    wire N__18398;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18360;
    wire N__18359;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18343;
    wire N__18338;
    wire N__18335;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18310;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18292;
    wire N__18291;
    wire N__18288;
    wire N__18287;
    wire N__18286;
    wire N__18285;
    wire N__18284;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18261;
    wire N__18260;
    wire N__18257;
    wire N__18256;
    wire N__18255;
    wire N__18254;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18242;
    wire N__18237;
    wire N__18230;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18223;
    wire N__18222;
    wire N__18213;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18186;
    wire N__18183;
    wire N__18170;
    wire N__18169;
    wire N__18168;
    wire N__18165;
    wire N__18164;
    wire N__18163;
    wire N__18162;
    wire N__18159;
    wire N__18158;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18146;
    wire N__18143;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18139;
    wire N__18138;
    wire N__18137;
    wire N__18136;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18121;
    wire N__18116;
    wire N__18109;
    wire N__18108;
    wire N__18107;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18093;
    wire N__18088;
    wire N__18085;
    wire N__18078;
    wire N__18073;
    wire N__18066;
    wire N__18063;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17989;
    wire N__17984;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17900;
    wire N__17897;
    wire N__17892;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17870;
    wire N__17867;
    wire N__17866;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17830;
    wire N__17829;
    wire N__17828;
    wire N__17825;
    wire N__17820;
    wire N__17819;
    wire N__17816;
    wire N__17811;
    wire N__17808;
    wire N__17803;
    wire N__17800;
    wire N__17795;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17772;
    wire N__17769;
    wire N__17764;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17732;
    wire N__17729;
    wire N__17728;
    wire N__17727;
    wire N__17726;
    wire N__17717;
    wire N__17714;
    wire N__17713;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17690;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17684;
    wire N__17681;
    wire N__17680;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17661;
    wire N__17658;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17633;
    wire N__17624;
    wire N__17621;
    wire N__17620;
    wire N__17619;
    wire N__17616;
    wire N__17615;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17601;
    wire N__17598;
    wire N__17597;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17545;
    wire N__17542;
    wire N__17541;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17530;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17487;
    wire N__17482;
    wire N__17471;
    wire N__17468;
    wire N__17467;
    wire N__17466;
    wire N__17463;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17445;
    wire N__17442;
    wire N__17437;
    wire N__17434;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17278;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17260;
    wire N__17255;
    wire N__17252;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17240;
    wire N__17237;
    wire N__17236;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17189;
    wire N__17186;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17168;
    wire N__17165;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17153;
    wire N__17150;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17117;
    wire N__17116;
    wire N__17115;
    wire N__17114;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17092;
    wire N__17087;
    wire N__17078;
    wire N__17077;
    wire N__17074;
    wire N__17073;
    wire N__17070;
    wire N__17069;
    wire N__17068;
    wire N__17067;
    wire N__17066;
    wire N__17065;
    wire N__17062;
    wire N__17057;
    wire N__17054;
    wire N__17045;
    wire N__17040;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16940;
    wire N__16937;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16877;
    wire N__16876;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16817;
    wire N__16816;
    wire N__16811;
    wire N__16808;
    wire N__16807;
    wire N__16806;
    wire N__16805;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16747;
    wire N__16742;
    wire N__16739;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16626;
    wire N__16621;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16585;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16577;
    wire N__16574;
    wire N__16569;
    wire N__16566;
    wire N__16559;
    wire N__16556;
    wire N__16555;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16544;
    wire N__16543;
    wire N__16538;
    wire N__16535;
    wire N__16530;
    wire N__16527;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16513;
    wire N__16512;
    wire N__16511;
    wire N__16508;
    wire N__16507;
    wire N__16500;
    wire N__16499;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16482;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16463;
    wire N__16458;
    wire N__16455;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16425;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16410;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16406;
    wire N__16403;
    wire N__16402;
    wire N__16401;
    wire N__16400;
    wire N__16399;
    wire N__16394;
    wire N__16393;
    wire N__16388;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16366;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16347;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16325;
    wire N__16316;
    wire N__16311;
    wire N__16306;
    wire N__16297;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16282;
    wire N__16279;
    wire N__16278;
    wire N__16277;
    wire N__16276;
    wire N__16275;
    wire N__16274;
    wire N__16273;
    wire N__16270;
    wire N__16269;
    wire N__16268;
    wire N__16267;
    wire N__16266;
    wire N__16265;
    wire N__16262;
    wire N__16261;
    wire N__16260;
    wire N__16259;
    wire N__16258;
    wire N__16257;
    wire N__16256;
    wire N__16255;
    wire N__16252;
    wire N__16251;
    wire N__16250;
    wire N__16249;
    wire N__16248;
    wire N__16247;
    wire N__16246;
    wire N__16245;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16241;
    wire N__16234;
    wire N__16231;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16221;
    wire N__16218;
    wire N__16217;
    wire N__16216;
    wire N__16215;
    wire N__16214;
    wire N__16213;
    wire N__16212;
    wire N__16209;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16189;
    wire N__16182;
    wire N__16181;
    wire N__16174;
    wire N__16167;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16128;
    wire N__16125;
    wire N__16118;
    wire N__16113;
    wire N__16110;
    wire N__16109;
    wire N__16106;
    wire N__16101;
    wire N__16098;
    wire N__16093;
    wire N__16090;
    wire N__16085;
    wire N__16080;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16061;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16037;
    wire N__16026;
    wire N__16023;
    wire N__15998;
    wire N__15997;
    wire N__15996;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15991;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15974;
    wire N__15971;
    wire N__15964;
    wire N__15959;
    wire N__15952;
    wire N__15947;
    wire N__15938;
    wire N__15937;
    wire N__15936;
    wire N__15935;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15918;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15876;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15851;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15838;
    wire N__15837;
    wire N__15836;
    wire N__15833;
    wire N__15832;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15817;
    wire N__15816;
    wire N__15815;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15811;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15797;
    wire N__15794;
    wire N__15787;
    wire N__15782;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15766;
    wire N__15765;
    wire N__15764;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15756;
    wire N__15755;
    wire N__15754;
    wire N__15751;
    wire N__15750;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15742;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15730;
    wire N__15723;
    wire N__15722;
    wire N__15721;
    wire N__15720;
    wire N__15719;
    wire N__15718;
    wire N__15715;
    wire N__15708;
    wire N__15703;
    wire N__15694;
    wire N__15689;
    wire N__15688;
    wire N__15685;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15665;
    wire N__15664;
    wire N__15659;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15643;
    wire N__15642;
    wire N__15641;
    wire N__15636;
    wire N__15631;
    wire N__15624;
    wire N__15615;
    wire N__15612;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15591;
    wire N__15588;
    wire N__15583;
    wire N__15572;
    wire N__15567;
    wire N__15562;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15521;
    wire N__15520;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15418;
    wire N__15413;
    wire N__15410;
    wire N__15409;
    wire N__15406;
    wire N__15405;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15391;
    wire N__15390;
    wire N__15389;
    wire N__15386;
    wire N__15381;
    wire N__15380;
    wire N__15379;
    wire N__15376;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15358;
    wire N__15353;
    wire N__15344;
    wire N__15343;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15329;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15314;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15294;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15275;
    wire N__15272;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15209;
    wire N__15206;
    wire N__15205;
    wire N__15202;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15176;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15164;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15146;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15135;
    wire N__15130;
    wire N__15129;
    wire N__15128;
    wire N__15127;
    wire N__15124;
    wire N__15121;
    wire N__15116;
    wire N__15113;
    wire N__15104;
    wire N__15101;
    wire N__15100;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15086;
    wire N__15083;
    wire N__15078;
    wire N__15075;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14991;
    wire N__14990;
    wire N__14989;
    wire N__14984;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14973;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14947;
    wire N__14942;
    wire N__14939;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14925;
    wire N__14922;
    wire N__14921;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14898;
    wire N__14893;
    wire N__14892;
    wire N__14891;
    wire N__14890;
    wire N__14889;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14846;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14838;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14813;
    wire N__14812;
    wire N__14811;
    wire N__14810;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14790;
    wire N__14789;
    wire N__14786;
    wire N__14785;
    wire N__14784;
    wire N__14783;
    wire N__14782;
    wire N__14781;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14761;
    wire N__14756;
    wire N__14751;
    wire N__14746;
    wire N__14739;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14701;
    wire N__14700;
    wire N__14697;
    wire N__14696;
    wire N__14695;
    wire N__14694;
    wire N__14691;
    wire N__14690;
    wire N__14689;
    wire N__14688;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14662;
    wire N__14661;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14623;
    wire N__14622;
    wire N__14621;
    wire N__14618;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14606;
    wire N__14601;
    wire N__14596;
    wire N__14593;
    wire N__14588;
    wire N__14585;
    wire N__14580;
    wire N__14573;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14521;
    wire N__14520;
    wire N__14519;
    wire N__14518;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14502;
    wire N__14495;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14487;
    wire N__14482;
    wire N__14481;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14473;
    wire N__14472;
    wire N__14471;
    wire N__14470;
    wire N__14469;
    wire N__14466;
    wire N__14459;
    wire N__14454;
    wire N__14451;
    wire N__14442;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14430;
    wire N__14425;
    wire N__14422;
    wire N__14421;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14403;
    wire N__14400;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14361;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14311;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14303;
    wire N__14300;
    wire N__14299;
    wire N__14298;
    wire N__14297;
    wire N__14294;
    wire N__14289;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14273;
    wire N__14270;
    wire N__14265;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14203;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14186;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14176;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14146;
    wire N__14145;
    wire N__14144;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14126;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14071;
    wire N__14070;
    wire N__14067;
    wire N__14062;
    wire N__14057;
    wire N__14056;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14038;
    wire N__14037;
    wire N__14036;
    wire N__14035;
    wire N__14034;
    wire N__14033;
    wire N__14032;
    wire N__14029;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14021;
    wire N__14020;
    wire N__14017;
    wire N__14012;
    wire N__14009;
    wire N__14004;
    wire N__14003;
    wire N__14002;
    wire N__14001;
    wire N__13998;
    wire N__13997;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13983;
    wire N__13976;
    wire N__13971;
    wire N__13966;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13952;
    wire N__13947;
    wire N__13944;
    wire N__13939;
    wire N__13928;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13922;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13907;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13884;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13864;
    wire N__13863;
    wire N__13862;
    wire N__13861;
    wire N__13860;
    wire N__13859;
    wire N__13856;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13826;
    wire N__13811;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13799;
    wire N__13796;
    wire N__13795;
    wire N__13794;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13772;
    wire N__13771;
    wire N__13768;
    wire N__13767;
    wire N__13766;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13724;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13718;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13703;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13642;
    wire N__13639;
    wire N__13636;
    wire N__13633;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13612;
    wire N__13611;
    wire N__13608;
    wire N__13603;
    wire N__13598;
    wire N__13597;
    wire N__13596;
    wire N__13595;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13581;
    wire N__13578;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13540;
    wire N__13537;
    wire N__13534;
    wire N__13527;
    wire N__13520;
    wire N__13517;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13507;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13490;
    wire N__13487;
    wire N__13486;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13412;
    wire N__13409;
    wire N__13402;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13336;
    wire N__13331;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13310;
    wire N__13309;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13302;
    wire N__13297;
    wire N__13294;
    wire N__13289;
    wire N__13286;
    wire N__13277;
    wire N__13276;
    wire N__13273;
    wire N__13272;
    wire N__13271;
    wire N__13270;
    wire N__13269;
    wire N__13268;
    wire N__13267;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13251;
    wire N__13248;
    wire N__13239;
    wire N__13232;
    wire N__13231;
    wire N__13230;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13212;
    wire N__13211;
    wire N__13208;
    wire N__13203;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13182;
    wire N__13175;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13163;
    wire N__13160;
    wire N__13159;
    wire N__13158;
    wire N__13157;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13142;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13065;
    wire N__13060;
    wire N__13055;
    wire N__13054;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13041;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13012;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__13001;
    wire N__12998;
    wire N__12993;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12978;
    wire N__12977;
    wire N__12974;
    wire N__12973;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12959;
    wire N__12954;
    wire N__12949;
    wire N__12942;
    wire N__12929;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12911;
    wire N__12908;
    wire N__12903;
    wire N__12900;
    wire N__12899;
    wire N__12898;
    wire N__12891;
    wire N__12890;
    wire N__12887;
    wire N__12886;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12866;
    wire N__12861;
    wire N__12856;
    wire N__12849;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12814;
    wire N__12813;
    wire N__12806;
    wire N__12803;
    wire N__12798;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12761;
    wire N__12758;
    wire N__12753;
    wire N__12750;
    wire N__12749;
    wire N__12746;
    wire N__12745;
    wire N__12742;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12722;
    wire N__12721;
    wire N__12720;
    wire N__12719;
    wire N__12716;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12688;
    wire N__12687;
    wire N__12682;
    wire N__12679;
    wire N__12678;
    wire N__12677;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12669;
    wire N__12668;
    wire N__12665;
    wire N__12664;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12650;
    wire N__12645;
    wire N__12640;
    wire N__12637;
    wire N__12636;
    wire N__12633;
    wire N__12632;
    wire N__12631;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12597;
    wire N__12590;
    wire N__12575;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12567;
    wire N__12560;
    wire N__12557;
    wire N__12556;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12541;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12521;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12506;
    wire N__12505;
    wire N__12502;
    wire N__12501;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12485;
    wire N__12482;
    wire N__12481;
    wire N__12480;
    wire N__12479;
    wire N__12478;
    wire N__12477;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12439;
    wire N__12432;
    wire N__12427;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12402;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12386;
    wire N__12383;
    wire N__12374;
    wire N__12367;
    wire N__12362;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12298;
    wire N__12297;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12287;
    wire N__12286;
    wire N__12283;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12241;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12226;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12193;
    wire N__12188;
    wire N__12185;
    wire N__12184;
    wire N__12179;
    wire N__12176;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12169;
    wire N__12162;
    wire N__12159;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12139;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12085;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12068;
    wire N__12065;
    wire N__12064;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12017;
    wire N__12014;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11992;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11980;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11945;
    wire N__11936;
    wire N__11933;
    wire N__11932;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11916;
    wire N__11915;
    wire N__11914;
    wire N__11913;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11898;
    wire N__11893;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11861;
    wire N__11860;
    wire N__11859;
    wire N__11858;
    wire N__11853;
    wire N__11848;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11773;
    wire N__11772;
    wire N__11771;
    wire N__11766;
    wire N__11765;
    wire N__11762;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11735;
    wire N__11726;
    wire N__11725;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11714;
    wire N__11711;
    wire N__11704;
    wire N__11699;
    wire N__11698;
    wire N__11697;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11680;
    wire N__11679;
    wire N__11678;
    wire N__11675;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11642;
    wire N__11639;
    wire N__11634;
    wire N__11631;
    wire N__11624;
    wire N__11619;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11560;
    wire N__11557;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11540;
    wire N__11539;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11529;
    wire N__11528;
    wire N__11527;
    wire N__11526;
    wire N__11523;
    wire N__11516;
    wire N__11511;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11464;
    wire N__11459;
    wire N__11456;
    wire N__11455;
    wire N__11454;
    wire N__11451;
    wire N__11450;
    wire N__11449;
    wire N__11438;
    wire N__11435;
    wire N__11434;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11413;
    wire N__11410;
    wire N__11405;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11383;
    wire N__11378;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11363;
    wire N__11360;
    wire N__11359;
    wire N__11358;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11336;
    wire N__11335;
    wire N__11334;
    wire N__11331;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11252;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11231;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11188;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11179;
    wire N__11170;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11114;
    wire N__11111;
    wire N__11106;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11029;
    wire N__11022;
    wire N__11019;
    wire N__11014;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10941;
    wire N__10936;
    wire N__10933;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10790;
    wire N__10783;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10756;
    wire N__10751;
    wire N__10748;
    wire N__10747;
    wire N__10746;
    wire N__10743;
    wire N__10738;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10726;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10714;
    wire N__10713;
    wire N__10706;
    wire N__10703;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10689;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10666;
    wire N__10663;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10598;
    wire N__10591;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10560;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10443;
    wire N__10438;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10434;
    wire N__10433;
    wire N__10432;
    wire N__10427;
    wire N__10422;
    wire N__10415;
    wire N__10412;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10360;
    wire N__10357;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10109;
    wire N__10106;
    wire N__10105;
    wire N__10104;
    wire N__10103;
    wire N__10102;
    wire N__10097;
    wire N__10090;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10074;
    wire N__10071;
    wire N__10066;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10036;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire \Clock50MHz.PixelClock ;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_1_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7;
    wire bfn_1_2_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6;
    wire bfn_1_3_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire beamY_RNITSR8_0Z0Z_8;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0;
    wire beamY_RNISI4A_0Z0Z_9;
    wire beamY_RNIE925Z0Z_6_cascade_;
    wire beamY_RNIKOP3_0Z0Z_6;
    wire un5_visibley_c2_cascade_;
    wire un5_visibley_c6_0_0_0;
    wire bfn_1_6_0_;
    wire un20_beamy_cry_1;
    wire un20_beamy_cry_2;
    wire un20_beamy_cry_3;
    wire un20_beamy_cry_4;
    wire un20_beamy_cry_5;
    wire un20_beamy_cry_6;
    wire un20_beamy_cry_7;
    wire un20_beamy_cry_8;
    wire bfn_1_7_0_;
    wire if_generate_plus_mult1_un75_sum_axbxc5_0_x1;
    wire if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_;
    wire bfn_1_9_0_;
    wire un1_voltage_0_cry_0;
    wire un1_voltage_0_cry_1;
    wire un1_voltage_0_cry_2;
    wire N_1503_cascade_;
    wire SDATA1_ibuf_RNILOUGZ0Z2;
    wire un1_voltage_1_1_axb_0_cascade_;
    wire voltage_0_1_sqmuxa_1_cascade_;
    wire voltage_3_9_iv_0_0_cascade_;
    wire N_1507;
    wire N_1507_cascade_;
    wire voltage_3_RNO_0Z0Z_0;
    wire bfn_1_12_0_;
    wire un1_voltage_3_1_cry_0;
    wire un1_voltage_3_1_cry_1;
    wire un1_voltage_3_1_cry_2;
    wire ScreenBuffer_0_0_1_sqmuxa;
    wire un4_voltage_2_0__N_13_mux_iZ0_cascade_;
    wire SDATA1_ibuf_RNI098KZ0Z2;
    wire N_35_0_i_cascade_;
    wire un4_voltage_10_9__N_4_cascade_;
    wire un4_voltage_2_0__N_5_iZ0;
    wire voltage_0_1_sqmuxa_cascade_;
    wire un1_voltage_0_cry_0_0_c_RNOZ0;
    wire N_34_0_i;
    wire N_41_i;
    wire N_41_i_cascade_;
    wire voltage_0_1_sqmuxa;
    wire ScreenBuffer_0_1_1_sqmuxa_2;
    wire un4_voltage_2_0__i2_mux;
    wire bfn_2_1_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0;
    wire un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_;
    wire un5_visibley_axbxc7_1_cascade_;
    wire chary_if_generate_plus_mult1_un33_sum_axb3_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz;
    wire chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_;
    wire beamY_RNI9425_0Z0Z_6_cascade_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_;
    wire beamY_RNI9425Z0Z_6_cascade_;
    wire if_generate_plus_mult1_un61_sum_ac0_x0;
    wire if_generate_plus_mult1_un61_sum_ac0_x1;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0_6;
    wire row_1_if_generate_plus_mult1_un61_sum_c4_d;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_;
    wire beamY_RNI75QM4Z0Z_5_cascade_;
    wire if_generate_plus_mult1_un68_sum_axbxc5_x0;
    wire if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8;
    wire if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0;
    wire if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_;
    wire beamY_RNI75QM4Z0Z_5;
    wire voltage_0_10_iv_0_2_cascade_;
    wire voltage_0_RNO_0Z0Z_2;
    wire voltage_1_9_iv_0_2_cascade_;
    wire voltage_3_RNO_0Z0Z_2;
    wire voltage_3_9_iv_0_2_cascade_;
    wire CO2_3_cascade_;
    wire N_1155_cascade_;
    wire voltage_0_10_iv_0_3;
    wire N_1519;
    wire N_1521;
    wire counter_RNI49LH1_0Z0Z_0;
    wire voltage_1_9_iv_0_0;
    wire CO1_3;
    wire voltage_2_1_sqmuxa_cascade_;
    wire N_1155;
    wire voltage_1_1_sqmuxa;
    wire voltage_1_1_sqmuxa_cascade_;
    wire voltage_1_9_iv_0_3;
    wire voltage_3_RNO_0Z0Z_3;
    wire voltage_3_9_iv_0_3;
    wire N_1510;
    wire N_1506_cascade_;
    wire counter_RNIGLLH1Z0Z_0_cascade_;
    wire N_2063;
    wire N_1522;
    wire un1_voltage_1_1_cry_0_0_c_RNOZ0;
    wire bfn_2_13_0_;
    wire counter_RNILOUG2Z0Z_3;
    wire un1_voltage_1_1_cry_0;
    wire counter_RNIT58K2Z0Z_2;
    wire voltage_1_RNO_0Z0Z_2;
    wire un1_voltage_1_1_cry_1;
    wire un1_voltage_1_1_cry_2;
    wire voltage_1_RNO_0Z0Z_3;
    wire un6_slaveselectlto9_1_cascade_;
    wire un6_slaveselect_0_cascade_;
    wire un3_slaveselectlt9;
    wire bfn_2_14_0_;
    wire voltage_2_RNIKG123Z0Z_1;
    wire un1_voltage_2_1_cry_0;
    wire counter_RNI2RBA2Z0Z_3;
    wire un1_voltage_2_1_cry_1;
    wire un1_voltage_2_1_axb_3;
    wire voltage_2_9_iv_0_3;
    wire un1_voltage_2_1_cry_2;
    wire N_46_1;
    wire un1_sclk17_2_1_cascade_;
    wire un1_sclk17_1_1_cascade_;
    wire bfn_4_1_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7;
    wire bfn_4_2_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7;
    wire bfn_4_3_0_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0;
    wire un5_visibley_c2;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_;
    wire beamY_RNIEDF31Z0Z_6;
    wire chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_c4_3_1;
    wire chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_6_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0;
    wire row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0;
    wire row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0;
    wire beamY_RNIFS4TZ0Z_7;
    wire beamY_RNIFS4TZ0Z_7_cascade_;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_;
    wire beamY_RNIQTGS2Z0Z_8_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb3_cascade_;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0;
    wire beamY_RNIQTGS2Z0Z_8;
    wire chary_if_generate_plus_mult1_un54_sum_c4;
    wire beamY_RNI0K169Z0Z_6_cascade_;
    wire un5_visibley_0_29;
    wire chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_;
    wire if_m1_x1_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_c5;
    wire row_1_if_generate_plus_mult1_un61_sum_axb4_i;
    wire if_m1_x0;
    wire un113_pixel_3_0_11__g1_0;
    wire chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_;
    wire GB_BUFFER_Clock12MHz_c_g_THRU_CO;
    wire N_1159_i;
    wire N_1154;
    wire N_1159_i_cascade_;
    wire voltage_2_1_sqmuxa;
    wire voltage_0_0_sqmuxa_1;
    wire slaveselect_RNILOQC2Z0Z_1;
    wire slaveselect_RNILOQC2Z0Z_1_cascade_;
    wire counter_RNICHLH1Z0Z_0;
    wire un1_voltage_012_0_cascade_;
    wire un74_voltage_0;
    wire N_1153;
    wire voltage_0_1_sqmuxa_1;
    wire N_1153_cascade_;
    wire voltage_3_1_sqmuxa;
    wire voltage_3_RNO_0Z0Z_1;
    wire voltage_3_9_iv_0_1_cascade_;
    wire un1_voltage_012_0;
    wire voltage_1_9_iv_0_1;
    wire voltage_1_RNO_0Z0Z_1;
    wire N_1504_cascade_;
    wire N_1504;
    wire counter_RNI8DLH1Z0Z_0;
    wire N_1508;
    wire slaveselect_RNILOQC2Z0Z_2;
    wire bfn_4_13_0_;
    wire counter_cry_1;
    wire counter_cry_2;
    wire counter_cry_3;
    wire counter_cry_4;
    wire counter_cry_5;
    wire counter_cry_6;
    wire counter_cry_7;
    wire counter_cry_8;
    wire bfn_4_14_0_;
    wire un1_counter_i_0;
    wire bfn_5_3_0_;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_;
    wire chessboardpixel_un173_pixellt10;
    wire chessboardpixel_un151_pixel_27;
    wire chessboardpixel_un177_pixel_26_cascade_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0;
    wire beamY_i_2;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0;
    wire un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_;
    wire chessboardpixel_un199_pixellt10;
    wire un113_pixel_4_0_15__un1_beamylto9_3;
    wire VSync_c;
    wire un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_;
    wire beamY_RNII8O41Z0Z_9;
    wire un113_pixel_4_0_15__g0_i_a3_0Z0Z_4;
    wire if_m1_5;
    wire if_generate_plus_mult1_un54_sum_axbxc5_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_cZ0Z4;
    wire if_generate_plus_mult1_un75_sum_ac0_5_x1;
    wire row_1_if_i2_mux_0_cascade_;
    wire if_generate_plus_mult1_un75_sum_ac0_5_x0;
    wire row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_;
    wire un5_visibley_c5;
    wire beamY_RNIJNLCZ0Z_9;
    wire beamY_RNIJNLCZ0Z_9_cascade_;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum;
    wire beamY_RNIVGU01Z0Z_9;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0;
    wire row_1_if_generate_plus_mult1_un75_sum_ac0_5;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum;
    wire if_generate_plus_mult1_un75_sum_c5_x0;
    wire if_generate_plus_mult1_un75_sum_c5_x1_cascade_;
    wire beamY_RNIPNEA3_0Z0Z_6;
    wire beamY_RNI0K169Z0Z_6;
    wire chary_if_generate_plus_mult1_un61_sum_c4;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9;
    wire chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_;
    wire beamYZ0Z_6;
    wire beamYZ0Z_5;
    wire chary_if_generate_plus_mult1_un75_sum_c5_N_9;
    wire beamY_RNIPLAE31Z0Z_4_cascade_;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0;
    wire beamY_RNIV42D31_0Z0Z_6;
    wire un113_pixel_3_0_11__N_4_i_0;
    wire g1_0_0;
    wire chary_if_generate_plus_mult1_un61_sum_axb3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum;
    wire beamY_RNIV42D31Z0Z_6;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_axbxc5_0;
    wire un113_pixel_3_0_11__g0_0_x2_0Z0Z_0;
    wire un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0;
    wire N_1520;
    wire un1_voltage_2_1_cry_0_c_RNOZ0;
    wire voltage_2_9_iv_0_0;
    wire un1_voltage_2_1_axb_0_cascade_;
    wire voltage_2_9_iv_0_2;
    wire voltage_2_RNO_0Z0Z_2;
    wire un1_voltage_012_3_0;
    wire voltage_2_9_iv_0_1;
    wire voltage_2_RNO_0Z0Z_1;
    wire un42_cry_1_c_RNOZ0;
    wire bfn_5_11_0_;
    wire un42_cry_1;
    wire counter_RNIGLLH1Z0Z_0;
    wire un42_cry_2;
    wire voltage_011_0;
    wire un42_cry_3;
    wire voltage_011;
    wire ScreenBuffer_1_122_1_cascade_;
    wire ScreenBuffer_1_3_1_sqmuxa;
    wire ScreenBuffer_1_0_1_sqmuxa;
    wire Z_decfrac4;
    wire un1_sclk17_0_0_cascade_;
    wire un39_0_3;
    wire un39_0_3_cascade_;
    wire un5_slaveselect_1;
    wire un5_slaveselect_1_cascade_;
    wire ScreenBuffer_1_122_1;
    wire un39_0_6;
    wire ScreenBuffer_1_2_1_sqmuxa;
    wire ScreenBuffer_1_2_1_sqmuxa_cascade_;
    wire un10_slaveselect;
    wire slaveselect_RNILOQC2Z0Z_0_cascade_;
    wire Z_decfrac4_2;
    wire counterZ0Z_9;
    wire counterZ0Z_7;
    wire un1_counter_1lto9_2_cascade_;
    wire un10_slaveselectlt4;
    wire counterZ0Z_4;
    wire un1_counter_1lt9;
    wire counterZ0Z_6;
    wire counterZ0Z_5;
    wire counterZ0Z_8;
    wire slaveselect_1lto9_4;
    wire slaveselect_1lto9_3;
    wire SCLK1_0_i;
    wire bfn_6_2_0_;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum;
    wire un113_pixel_4_0_15__un5_beamx_2Z0Z_0;
    wire un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_;
    wire un5_beamx_0;
    wire un5_beamx_0_cascade_;
    wire un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_;
    wire un13_beamylt6_0;
    wire un13_beamylt6_0_cascade_;
    wire un18_beamylt4;
    wire un113_pixel_4_0_15__un4_rowZ0Z_2;
    wire if_generate_plus_mult1_un54_sum_axbxc5;
    wire r_N_6;
    wire un113_pixel_4_0_15__un3_beamxZ0Z_7;
    wire un1_beamxlt10_0_cascade_;
    wire HSync_c;
    wire un18_beamylt10_0;
    wire if_generate_plus_mult1_un82_sum_axbxc5_0_x1;
    wire if_generate_plus_mult1_un82_sum_axbxc5_0_x0;
    wire un1_beamy_4;
    wire row_1_if_generate_plus_mult1_un68_sum_i_5;
    wire un113_pixel_4_0_15__un4_rowZ0Z_5;
    wire un13_beamy_0;
    wire chessboardpixel_un174_pixel;
    wire un4_row_cascade_;
    wire beamYZ0Z_9;
    wire beamYZ0Z_8;
    wire beamYZ0Z_7;
    wire un4_beamylt8_0;
    wire un4_beamy_0;
    wire un113_pixel_4_0_15__un8_beamylto9Z0Z_1;
    wire beamYZ0Z_4;
    wire un8_beamy;
    wire N_6_i;
    wire N_6_i_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3;
    wire beamYZ0Z_3;
    wire un4_beamylt6;
    wire if_m1_ns;
    wire if_m2_2_cascade_;
    wire row_1_if_generate_plus_mult1_un82_sum_axbxc5_0;
    wire bfn_6_9_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4;
    wire bfn_6_10_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_i;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803;
    wire voltage_2Z0Z_0;
    wire voltage_1Z0Z_0;
    wire voltage_2Z0Z_2;
    wire voltage_1Z0Z_2;
    wire voltage_2Z0Z_3;
    wire voltage_1Z0Z_3;
    wire voltage_2Z0Z_1;
    wire voltage_1Z0Z_1;
    wire un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0;
    wire N_1505;
    wire N_1509;
    wire un42_cry_2_c_RNOZ0;
    wire un1_sclk17_6_1_cascade_;
    wire un1_sclk17_3_1_cascade_;
    wire ScreenBuffer_0_0_1_sqmuxa_0;
    wire slaveselect_RNILOQCZ0Z2;
    wire un1_sclk17_8_0_0_cascade_;
    wire voltage_3Z0Z_2;
    wire voltage_0Z0Z_2;
    wire un1_sclk17_7_1;
    wire un5_slaveselect;
    wire SDATA2_c;
    wire un1_sclk17_9_1_cascade_;
    wire counterZ0Z_3;
    wire counterZ0Z_0;
    wire counterZ0Z_2;
    wire counterZ0Z_1;
    wire un1_sclk17_4_1;
    wire bfn_7_2_0_;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i;
    wire bfn_7_4_0_;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_0;
    wire bfn_7_5_0_;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538;
    wire charx_if_generate_plus_mult1_un33_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_;
    wire charx_if_generate_plus_mult1_un26_sum_i_5;
    wire bfn_7_6_0_;
    wire charx_if_generate_plus_mult1_un33_sum_i;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_3;
    wire charx_if_generate_plus_mult1_un40_sum_axb_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4;
    wire un113_pixel_4_0_15__un18_beamylto9Z0Z_2;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0;
    wire charx_if_generate_plus_mult1_un33_sum_i_5;
    wire un1_beamx_2;
    wire charx_i_24;
    wire charx_if_generate_plus_mult1_un1_sum_axb1_cascade_;
    wire font_un3_pixel_28_cascade_;
    wire un113_pixel_4_0_15__un15_beamyZ0Z_2;
    wire un13_beamy;
    wire font_un61_pixel_cascade_;
    wire un4_row;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf;
    wire charx_23;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3;
    wire charx_if_generate_plus_mult1_un1_sum_axb1;
    wire N_9_i_cascade_;
    wire N_13_0;
    wire ScreenBuffer_0_8Z0Z_0;
    wire ScreenBuffer_1_0Z0Z_0;
    wire currentchar_1_9_ns_1_0_cascade_;
    wire ScreenBuffer_1_1Z0Z_0;
    wire currentchar_1_6_ns_1_0_cascade_;
    wire ScreenBuffer_0_1Z0Z_0;
    wire ScreenBuffer_1_0Z0Z_4;
    wire ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_;
    wire ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_;
    wire row_1_if_generate_plus_mult1_un75_sum_c5;
    wire row_1_if_generate_plus_mult1_un68_sum_cZ0Z4;
    wire row_1_if_generate_plus_mult1_un75_sum_axbxc5_0;
    wire ScreenBuffer_1_2Z0Z_0;
    wire un3_rowlto1_cascade_;
    wire ScreenBuffer_0_2Z0Z_0;
    wire ScreenBuffer_1_1_1_sqmuxa;
    wire ScreenBuffer_0_0Z0Z_0;
    wire ScreenBuffer_1_1Z0Z_4;
    wire ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_;
    wire currentchar_1_11_ns_1_4;
    wire ScreenBuffer_1_2_RNIUP6F2FZ0Z_4;
    wire ScreenBuffer_1_3Z0Z_4;
    wire ScreenBuffer_1_3_RNIVS9G2FZ0Z_4;
    wire g1Z0Z_1_cascade_;
    wire N_1428_0_cascade_;
    wire un113_pixel_4_0_15__g1_1_cascade_;
    wire N_1300_0;
    wire un112_pixel_0_2_cascade_;
    wire N_1293_0;
    wire slaveselect_RNILOQC2Z0Z_0;
    wire ScreenBuffer_1_2Z0Z_4;
    wire ScreenBuffer_1_3Z0Z_2;
    wire ScreenBuffer_1_0Z0Z_2;
    wire un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_;
    wire un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_;
    wire m10_0_x1;
    wire un112_pixel_2_2_cascade_;
    wire un113_pixel_3_0_11__g0_0Z0Z_0;
    wire ScreenBuffer_0_7_RNIHMH43T2Z0Z_0;
    wire beamY_RNIDQUNU91Z0Z_0_cascade_;
    wire un115_pixel_2_sn_5_cascade_;
    wire un112_pixel_7_cascade_;
    wire beamY_RNIINK7J73Z0Z_0;
    wire bfn_8_1_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_8_2_0_;
    wire un3_beamx_0;
    wire un8_beamx_cry_9;
    wire beamXZ0Z_10;
    wire bfn_8_3_0_;
    wire beamXZ0Z_1;
    wire un5_visiblex_cry_0;
    wire beamXZ0Z_2;
    wire un5_visiblex_cry_1;
    wire beamXZ0Z_3;
    wire un5_visiblex_cry_2;
    wire beamXZ0Z_4;
    wire un5_visiblex_cry_3;
    wire beamXZ0Z_5;
    wire un5_visiblex_cry_4;
    wire beamXZ0Z_6;
    wire un5_visiblex_cry_5;
    wire beamXZ0Z_7;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire beamXZ0Z_8;
    wire bfn_8_4_0_;
    wire beamXZ0Z_9;
    wire un5_visiblex_cry_8;
    wire CO3_0_cascade_;
    wire charx_if_generate_plus_mult1_un26_sum_s_2_sf;
    wire chary_if_generate_plus_mult1_un33_sum_axb3;
    wire chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3;
    wire N_13;
    wire un113_pixel_4_0_15__un4_rowZ0Z_1;
    wire un1_voltage_0_axb_0;
    wire voltage_0_10_iv_0_0;
    wire un1_voltage_012_2_0;
    wire voltage_0_10_iv_0_1;
    wire voltage_0_RNO_0Z0Z_1;
    wire nCS1_c;
    wire un1_counter_1_0;
    wire voltage_0_0_sqmuxa_1_g;
    wire voltage_3Z0Z_0;
    wire voltage_0Z0Z_0;
    wire un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0;
    wire bfn_8_7_0_;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2;
    wire charx_if_generate_plus_mult1_un68_sum_i_5;
    wire charx_if_generate_plus_mult1_un75_sum_cry_3;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1;
    wire charx_if_generate_plus_mult1_un68_sum_i;
    wire bfn_8_8_0_;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_1;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_4;
    wire column_1_if_generate_plus_mult1_un61_sum_iZ0;
    wire chary_24;
    wire un113_pixel_4_0_15__gZ0Z2;
    wire font_un3_pixel_30;
    wire un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1;
    wire font_un57_pixel_cascade_;
    wire currentchar_1_5;
    wire font_un67_pixel_ac0_5;
    wire font_un64_pixel_ac0_5;
    wire un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_;
    wire N_12;
    wire un113_pixel_4_0_15__g0_iZ0Z_2;
    wire un113_pixel_4_0_15__g0_iZ0Z_5_cascade_;
    wire beamXZ0Z_0;
    wire un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6;
    wire beamY_RNIOEPPEK1Z0Z_0_cascade_;
    wire un112_pixel_1_2;
    wire N_3461_0_cascade_;
    wire N_4568_0_cascade_;
    wire N_1305_0;
    wire un113_pixel_4_0_15__g0_0Z0Z_2;
    wire Pixel_3_sqmuxa_0;
    wire g0_1_1;
    wire N_1_0_cascade_;
    wire ScreenBuffer_1_3Z0Z_3;
    wire ScreenBuffer_1_1Z0Z_3;
    wire ScreenBuffer_1_2Z0Z_3;
    wire un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_;
    wire un113_pixel_3_0_11__currentchar_N_13_cascade_;
    wire voltage_3Z0Z_3;
    wire voltage_0Z0Z_3;
    wire ScreenBuffer_1_0Z0Z_3;
    wire un113_pixel_4_0_15__g0_1Z0Z_0;
    wire un113_pixel_4_0_15__g0_3_0;
    wire voltage_3Z0Z_1;
    wire slaveselectZ0;
    wire voltage_0Z0Z_1;
    wire un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0;
    wire ScreenBuffer_0_12Z0Z_0;
    wire ScreenBuffer_0_4Z0Z_0;
    wire ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_;
    wire ScreenBuffer_0_6Z0Z_0;
    wire ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_;
    wire currentchar_m7_0_cascade_;
    wire ScreenBuffer_0_7Z0Z_0;
    wire ScreenBuffer_0_5Z0Z_0;
    wire un113_pixel_3_0_11__currentchar_N_13;
    wire un112_pixel_1_2_x1;
    wire un112_pixel_2_8_cascade_;
    wire un115_pixel_4_am_7;
    wire N_1287_cascade_;
    wire currentchar_1_0_cascade_;
    wire un115_pixel_4_bm_7;
    wire ScreenBuffer_0_7_RNII0GVLQZ0Z_0;
    wire un113_pixel_1_0_3__N_10_mux_cascade_;
    wire N_1285_0_0_0_cascade_;
    wire un113_pixel_3_0_11__g1_0_0_0;
    wire m14;
    wire m14_cascade_;
    wire beamY_RNI7RM4IFZ0Z_0;
    wire un113_pixel_3_0_11__g1_1_0;
    wire beamY_RNIPQEDM42Z0Z_0;
    wire N_1293;
    wire N_1306_cascade_;
    wire N_1327_0;
    wire m11_cascade_;
    wire un113_pixel_4_0_15__N_17;
    wire un115_pixel_6_bm_2_cascade_;
    wire N_1330;
    wire un115_pixel_6_am_2;
    wire bfn_9_1_0_;
    wire un5_visiblex_i_24;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12;
    wire bfn_9_2_0_;
    wire if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_1;
    wire if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx;
    wire if_generate_plus_mult1_un47_sum_0_cry_3_ma;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_2;
    wire N_1184_0_i;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_3;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_4;
    wire un5_visiblex_i_25;
    wire N_2110_i_cascade_;
    wire column_1_if_generate_plus_mult1_un47_sum0_5;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2;
    wire column_1_if_generate_plus_mult1_un47_sum0_3;
    wire if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum0_2;
    wire SDATA1_c;
    wire un1_sclk17_9_0_3;
    wire un1_sclk17_5_1_0;
    wire ScreenBuffer_0_9Z0Z_0;
    wire Clock12MHz_c_g;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4;
    wire column_1_if_generate_plus_mult1_un47_sum0_4;
    wire bfn_9_5_0_;
    wire if_generate_plus_mult1_un54_sum_axb_2_l_fx;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_1;
    wire if_generate_plus_mult1_un47_sum_m_5;
    wire if_generate_plus_mult1_un54_sum_axb_3_l_fx;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_2;
    wire if_generate_plus_mult1_un54_sum_axb_4_l_fx;
    wire N_2110_i;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_4;
    wire if_generate_plus_mult1_un54_sum_s_5_cascade_;
    wire bfn_9_6_0_;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2;
    wire charx_if_generate_plus_mult1_un54_sum_i_5;
    wire charx_if_generate_plus_mult1_un61_sum_cry_3;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum_i;
    wire bfn_9_7_0_;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0;
    wire charx_if_generate_plus_mult1_un75_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_3;
    wire charx_if_generate_plus_mult1_un68_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0;
    wire charx_if_generate_plus_mult1_un61_sum_i;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0;
    wire charx_if_generate_plus_mult1_un61_sum_i_5;
    wire bfn_9_8_0_;
    wire N_2096_i;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_s_5;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un54_sum_i_5;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_4;
    wire column_1_i_i_3;
    wire N_11;
    wire un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0;
    wire un113_pixel_4_0_15__g0_i_a3_2;
    wire Pixel_c;
    wire PixelClock_g;
    wire un113_pixel_7_1_7__g0_6Z0Z_0;
    wire N_3078_0;
    wire N_1297_0_cascade_;
    wire font_un67_pixel_ac0_5_0;
    wire chary_if_generate_plus_mult1_un68_sum_c5;
    wire chary_if_generate_plus_mult1_un1_sum_axbxc3_2;
    wire un113_pixel_4_0_15__g0_4_0Z0Z_0;
    wire beamYZ0Z_2;
    wire chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i;
    wire un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_;
    wire font_un3_pixel_28;
    wire N_1342;
    wire un113_pixel_4_0_15__g0_5Z0Z_1;
    wire font_un71_pixellt7_0_1;
    wire font_un64_pixel_ac0_5_0;
    wire un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3;
    wire font_un3_pixel_0_29;
    wire un113_pixel_4_0_15__g0_5Z0Z_4_cascade_;
    wire N_9;
    wire un113_pixel_4_0_15__g2Z0Z_0_cascade_;
    wire N_4566_0;
    wire un115_pixel_4;
    wire N_4564_0;
    wire N_5_0;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1;
    wire N_4561_0;
    wire g1_0;
    wire N_2075;
    wire un115_pixel_2_s_6_cascade_;
    wire un115_pixel_2_d_0_6_cascade_;
    wire un115_pixel_3_bm_6;
    wire ScreenBuffer_1_2Z0Z_1;
    wire ScreenBuffer_1_0Z0Z_1;
    wire N_1_7_0;
    wire ScreenBuffer_1_3Z0Z_1;
    wire ScreenBuffer_1_1Z0Z_1;
    wire m8;
    wire ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1;
    wire ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1;
    wire ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1;
    wire ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_;
    wire un113_pixel_3_0_11__gZ0Z1;
    wire un115_pixel_5_s_7;
    wire un115_pixel_5_am_7_cascade_;
    wire un115_pixel_5_bm_7;
    wire N_1288;
    wire un113_pixel_3_0_11__currentchar_1_4Z0Z_2;
    wire un113_pixel_4_0_15__g1Z0Z_0;
    wire m9;
    wire m9_cascade_;
    wire m6;
    wire m6_cascade_;
    wire beamY_RNICJUESD2Z0Z_0;
    wire N_1286_0_0_0;
    wire N_1289;
    wire font_un3_pixel_29;
    wire N_4562_0_0_0_cascade_;
    wire N_1340_0;
    wire beamY_RNICJUESD2_0Z0Z_0;
    wire beamY_RNI1H36941Z0Z_0;
    wire font_un125_pixel_1_bm;
    wire un113_pixel_6_1_5__N_11_cascade_;
    wire un113_pixel_2_0_3__N_8;
    wire beamY_RNICJUESD2_2Z0Z_0;
    wire m17;
    wire m12;
    wire un115_pixel_5_ns_x1_0;
    wire un115_pixel_5_ns_x0_0;
    wire N_1325_cascade_;
    wire un115_pixel_7_bm_0;
    wire N_1315_cascade_;
    wire N_1322;
    wire N_1329;
    wire N_1294_cascade_;
    wire beamY_RNICJUESD2_1Z0Z_0;
    wire N_1308;
    wire un115_pixel_5_d_2;
    wire un113_pixel_1_0_3__N_10_mux;
    wire beamY_RNIMR86ES2Z0Z_0;
    wire bfn_11_1_0_;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire CONSTANT_ONE_NET;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO;
    wire chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_2;
    wire bfn_11_3_0_;
    wire column_1_if_generate_plus_mult1_un47_sum1_2;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_1;
    wire column_1_if_generate_plus_mult1_un47_sum1_3;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_2;
    wire if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum1_4;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_3;
    wire un5_visiblex_cry_7_c_RNIVZ0Z952;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_4;
    wire column_1_if_generate_plus_mult1_un47_sum1_5;
    wire charx_if_generate_plus_mult1_un33_sum;
    wire un5_visiblex_i_0_25;
    wire N_56;
    wire N_32_i;
    wire if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx;
    wire CO3_0;
    wire charx_if_generate_plus_mult1_un26_sum_axb_3_i;
    wire charx_if_generate_plus_mult1_un54_sum;
    wire bfn_11_5_0_;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2;
    wire charx_if_generate_plus_mult1_un47_sum_i_5;
    wire charx_if_generate_plus_mult1_un61_sum_axb_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_3;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8;
    wire charx_if_generate_plus_mult1_un47_sum_i;
    wire charx_if_generate_plus_mult1_un47_sum;
    wire bfn_11_6_0_;
    wire charx_if_generate_plus_mult1_un40_sum_i_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2;
    wire charx_if_generate_plus_mult1_un54_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_3;
    wire charx_if_generate_plus_mult1_un47_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73;
    wire charx_if_generate_plus_mult1_un40_sum;
    wire charx_if_generate_plus_mult1_un40_sum_i;
    wire charx_if_generate_plus_mult1_un68_sum;
    wire bfn_11_9_0_;
    wire column_1_i_i_2;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_2;
    wire if_generate_plus_mult1_un75_sum_axb_4_l_fx;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_4;
    wire un6_rowlt7_0;
    wire chessboardpixel_un151_pixel_24;
    wire column_1_if_generate_plus_mult1_un68_sum_iZ0;
    wire un3_rowlto0;
    wire un113_pixel_3_0_11__currentchar_m7_0Z0Z_1;
    wire d_N_3_mux_cascade_;
    wire ScreenBuffer_1_2Z0Z_2;
    wire ScreenBuffer_1_1Z0Z_2;
    wire un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2;
    wire ScreenBuffer_0_10Z0Z_0;
    wire ScreenBuffer_0_11Z0Z_0;
    wire ScreenBuffer_1_3Z0Z_0;
    wire currentchar_1_5_ns_1_0_cascade_;
    wire ScreenBuffer_0_3Z0Z_0;
    wire beamY_RNIVDIFFI1Z0Z_0;
    wire beamY_RNI2RNL4M2Z0Z_0;
    wire un3_rowlto1;
    wire row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1;
    wire N_52;
    wire un112_pixel_2_8;
    wire N_4581_0_cascade_;
    wire N_1296_0_cascade_;
    wire N_1296_0;
    wire beamYZ0Z_1;
    wire N_1303_0;
    wire g0_16_x0_cascade_;
    wire g0_16_x1;
    wire N_4560_0;
    wire N_1309_0;
    wire un113_pixel_4_0_15__N_2;
    wire un113_pixel_7_1_7__N_9;
    wire beamY_RNIJIDRG11Z0Z_0_cascade_;
    wire beamY_RNIJIDRG11_0Z0Z_0;
    wire beamY_RNIRG0LHO1Z0Z_0_cascade_;
    wire ScreenBuffer_0_7_RNIB3R6U63Z0Z_0;
    wire font_un28_pixel_29;
    wire beamY_RNIRG0LHO1Z0Z_0;
    wire ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0;
    wire g0_2_x1_cascade_;
    wire g0_2_x0;
    wire N_1331_0;
    wire currentchar_1_2;
    wire currentchar_m7_0;
    wire un113_pixel_3_0_11__N_16_cascade_;
    wire un113_pixel_7_1_7__N_11;
    wire N_4573_0;
    wire un112_pixel_2_2;
    wire currentchar_1_1;
    wire beamYZ0Z_0;
    wire currentchar_1_0;
    wire un115_pixel_3_am_2;
    wire charx_if_generate_plus_mult1_un75_sum;
    wire bfn_12_9_0_;
    wire column_1_if_generate_plus_mult1_un75_sum_iZ0;
    wire G_673;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_1;
    wire if_generate_plus_mult1_un75_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_2;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire G_674;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_4;
    wire column_1_i_3;
    wire ScreenBuffer_0_10_RNIGDGIE9Z0Z_0;
    wire ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0;
    wire ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0;
    wire ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_;
    wire ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0;
    wire ScreenBuffer_0_6_RNIVTBDB12Z0Z_0;
    wire ScreenBuffer_0_6_RNITJ4B17Z0Z_0;
    wire un6_rowlto1;
    wire ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0;
    wire ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0;
    wire ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0;
    wire ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_;
    wire ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0;
    wire ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0;
    wire un6_rowlto0;
    wire column_1_i_2;
    wire ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_;
    wire ScreenBuffer_0_7_RNIN5F98I1Z0Z_0;
    wire un115_pixel_5_am_sx_1;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__11489),
            .RESETB(N__21892),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF Clock12MHz_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__26091),
            .GLOBALBUFFEROUTPUT(Clock12MHz_c_g));
    defparam Clock12MHz_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_gb_io_iopad (
            .OE(N__26093),
            .DIN(N__26092),
            .DOUT(N__26091),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_gb_io_preio (
            .PADOEN(N__26093),
            .PADOUT(N__26092),
            .PADIN(N__26091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__26082),
            .DIN(N__26081),
            .DOUT(N__26080),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__26082),
            .PADOUT(N__26081),
            .PADIN(N__26080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12338),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__26073),
            .DIN(N__26072),
            .DOUT(N__26071),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__26073),
            .PADOUT(N__26072),
            .PADIN(N__26071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SDATA2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SDATA2_obuf_iopad (
            .OE(N__26064),
            .DIN(N__26063),
            .DOUT(N__26062),
            .PACKAGEPIN(SDATA2));
    defparam SDATA2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SDATA2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SDATA2_obuf_preio (
            .PADOEN(N__26064),
            .PADOUT(N__26063),
            .PADIN(N__26062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16448),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK1_obuf_iopad (
            .OE(N__26055),
            .DIN(N__26054),
            .DOUT(N__26053),
            .PACKAGEPIN(SCLK1));
    defparam SCLK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCLK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCLK1_obuf_preio (
            .PADOEN(N__26055),
            .PADOUT(N__26054),
            .PADIN(N__26053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13679),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS2_obuf_iopad (
            .OE(N__26046),
            .DIN(N__26045),
            .DOUT(N__26044),
            .PACKAGEPIN(nCS2));
    defparam nCS2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS2_obuf_preio (
            .PADOEN(N__26046),
            .PADOUT(N__26045),
            .PADIN(N__26044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SDATA1_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SDATA1_ibuf_iopad (
            .OE(N__26037),
            .DIN(N__26036),
            .DOUT(N__26035),
            .PACKAGEPIN(SDATA1));
    defparam SDATA1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SDATA1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SDATA1_ibuf_preio (
            .PADOEN(N__26037),
            .PADOUT(N__26036),
            .PADIN(N__26035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SDATA1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS1_obuf_iopad (
            .OE(N__26028),
            .DIN(N__26027),
            .DOUT(N__26026),
            .PACKAGEPIN(nCS1));
    defparam nCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS1_obuf_preio (
            .PADOEN(N__26028),
            .PADOUT(N__26027),
            .PADIN(N__26026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__26019),
            .DIN(N__26018),
            .DOUT(N__26017),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__26019),
            .PADOUT(N__26018),
            .PADIN(N__26017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK2_obuf_iopad (
            .OE(N__26010),
            .DIN(N__26009),
            .DOUT(N__26008),
            .PACKAGEPIN(SCLK2));
    defparam SCLK2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCLK2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCLK2_obuf_preio (
            .PADOEN(N__26010),
            .PADOUT(N__26009),
            .PADIN(N__26008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13678),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__6199 (
            .O(N__25991),
            .I(N__25976));
    InMux I__6198 (
            .O(N__25990),
            .I(N__25976));
    InMux I__6197 (
            .O(N__25989),
            .I(N__25976));
    CascadeMux I__6196 (
            .O(N__25988),
            .I(N__25973));
    CascadeMux I__6195 (
            .O(N__25987),
            .I(N__25963));
    InMux I__6194 (
            .O(N__25986),
            .I(N__25953));
    InMux I__6193 (
            .O(N__25985),
            .I(N__25953));
    InMux I__6192 (
            .O(N__25984),
            .I(N__25950));
    InMux I__6191 (
            .O(N__25983),
            .I(N__25947));
    LocalMux I__6190 (
            .O(N__25976),
            .I(N__25944));
    InMux I__6189 (
            .O(N__25973),
            .I(N__25941));
    CascadeMux I__6188 (
            .O(N__25972),
            .I(N__25938));
    InMux I__6187 (
            .O(N__25971),
            .I(N__25932));
    InMux I__6186 (
            .O(N__25970),
            .I(N__25932));
    InMux I__6185 (
            .O(N__25969),
            .I(N__25929));
    InMux I__6184 (
            .O(N__25968),
            .I(N__25926));
    InMux I__6183 (
            .O(N__25967),
            .I(N__25921));
    InMux I__6182 (
            .O(N__25966),
            .I(N__25921));
    InMux I__6181 (
            .O(N__25963),
            .I(N__25918));
    InMux I__6180 (
            .O(N__25962),
            .I(N__25907));
    InMux I__6179 (
            .O(N__25961),
            .I(N__25907));
    InMux I__6178 (
            .O(N__25960),
            .I(N__25907));
    InMux I__6177 (
            .O(N__25959),
            .I(N__25907));
    InMux I__6176 (
            .O(N__25958),
            .I(N__25907));
    LocalMux I__6175 (
            .O(N__25953),
            .I(N__25902));
    LocalMux I__6174 (
            .O(N__25950),
            .I(N__25902));
    LocalMux I__6173 (
            .O(N__25947),
            .I(N__25899));
    Span4Mux_v I__6172 (
            .O(N__25944),
            .I(N__25896));
    LocalMux I__6171 (
            .O(N__25941),
            .I(N__25893));
    InMux I__6170 (
            .O(N__25938),
            .I(N__25888));
    InMux I__6169 (
            .O(N__25937),
            .I(N__25888));
    LocalMux I__6168 (
            .O(N__25932),
            .I(N__25885));
    LocalMux I__6167 (
            .O(N__25929),
            .I(N__25882));
    LocalMux I__6166 (
            .O(N__25926),
            .I(N__25875));
    LocalMux I__6165 (
            .O(N__25921),
            .I(N__25875));
    LocalMux I__6164 (
            .O(N__25918),
            .I(N__25875));
    LocalMux I__6163 (
            .O(N__25907),
            .I(N__25872));
    Span4Mux_v I__6162 (
            .O(N__25902),
            .I(N__25862));
    Span4Mux_v I__6161 (
            .O(N__25899),
            .I(N__25862));
    Span4Mux_v I__6160 (
            .O(N__25896),
            .I(N__25862));
    Span4Mux_h I__6159 (
            .O(N__25893),
            .I(N__25855));
    LocalMux I__6158 (
            .O(N__25888),
            .I(N__25855));
    Span4Mux_v I__6157 (
            .O(N__25885),
            .I(N__25855));
    Span4Mux_s2_h I__6156 (
            .O(N__25882),
            .I(N__25852));
    Span4Mux_s3_h I__6155 (
            .O(N__25875),
            .I(N__25847));
    Span4Mux_h I__6154 (
            .O(N__25872),
            .I(N__25847));
    InMux I__6153 (
            .O(N__25871),
            .I(N__25844));
    InMux I__6152 (
            .O(N__25870),
            .I(N__25841));
    InMux I__6151 (
            .O(N__25869),
            .I(N__25838));
    Odrv4 I__6150 (
            .O(N__25862),
            .I(column_1_i_3));
    Odrv4 I__6149 (
            .O(N__25855),
            .I(column_1_i_3));
    Odrv4 I__6148 (
            .O(N__25852),
            .I(column_1_i_3));
    Odrv4 I__6147 (
            .O(N__25847),
            .I(column_1_i_3));
    LocalMux I__6146 (
            .O(N__25844),
            .I(column_1_i_3));
    LocalMux I__6145 (
            .O(N__25841),
            .I(column_1_i_3));
    LocalMux I__6144 (
            .O(N__25838),
            .I(column_1_i_3));
    CascadeMux I__6143 (
            .O(N__25823),
            .I(N__25820));
    InMux I__6142 (
            .O(N__25820),
            .I(N__25814));
    InMux I__6141 (
            .O(N__25819),
            .I(N__25814));
    LocalMux I__6140 (
            .O(N__25814),
            .I(ScreenBuffer_0_10_RNIGDGIE9Z0Z_0));
    CascadeMux I__6139 (
            .O(N__25811),
            .I(N__25808));
    InMux I__6138 (
            .O(N__25808),
            .I(N__25802));
    InMux I__6137 (
            .O(N__25807),
            .I(N__25802));
    LocalMux I__6136 (
            .O(N__25802),
            .I(N__25799));
    Span4Mux_s0_h I__6135 (
            .O(N__25799),
            .I(N__25796));
    Span4Mux_h I__6134 (
            .O(N__25796),
            .I(N__25793));
    Odrv4 I__6133 (
            .O(N__25793),
            .I(ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0));
    InMux I__6132 (
            .O(N__25790),
            .I(N__25787));
    LocalMux I__6131 (
            .O(N__25787),
            .I(N__25784));
    Odrv12 I__6130 (
            .O(N__25784),
            .I(ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0));
    CascadeMux I__6129 (
            .O(N__25781),
            .I(ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_));
    InMux I__6128 (
            .O(N__25778),
            .I(N__25775));
    LocalMux I__6127 (
            .O(N__25775),
            .I(ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0));
    InMux I__6126 (
            .O(N__25772),
            .I(N__25769));
    LocalMux I__6125 (
            .O(N__25769),
            .I(N__25766));
    Span4Mux_s3_h I__6124 (
            .O(N__25766),
            .I(N__25763));
    Odrv4 I__6123 (
            .O(N__25763),
            .I(ScreenBuffer_0_6_RNIVTBDB12Z0Z_0));
    InMux I__6122 (
            .O(N__25760),
            .I(N__25756));
    InMux I__6121 (
            .O(N__25759),
            .I(N__25753));
    LocalMux I__6120 (
            .O(N__25756),
            .I(N__25750));
    LocalMux I__6119 (
            .O(N__25753),
            .I(N__25747));
    Odrv4 I__6118 (
            .O(N__25750),
            .I(ScreenBuffer_0_6_RNITJ4B17Z0Z_0));
    Odrv4 I__6117 (
            .O(N__25747),
            .I(ScreenBuffer_0_6_RNITJ4B17Z0Z_0));
    InMux I__6116 (
            .O(N__25742),
            .I(N__25729));
    InMux I__6115 (
            .O(N__25741),
            .I(N__25729));
    InMux I__6114 (
            .O(N__25740),
            .I(N__25726));
    InMux I__6113 (
            .O(N__25739),
            .I(N__25723));
    InMux I__6112 (
            .O(N__25738),
            .I(N__25720));
    InMux I__6111 (
            .O(N__25737),
            .I(N__25715));
    InMux I__6110 (
            .O(N__25736),
            .I(N__25715));
    InMux I__6109 (
            .O(N__25735),
            .I(N__25710));
    InMux I__6108 (
            .O(N__25734),
            .I(N__25710));
    LocalMux I__6107 (
            .O(N__25729),
            .I(N__25705));
    LocalMux I__6106 (
            .O(N__25726),
            .I(N__25694));
    LocalMux I__6105 (
            .O(N__25723),
            .I(N__25694));
    LocalMux I__6104 (
            .O(N__25720),
            .I(N__25694));
    LocalMux I__6103 (
            .O(N__25715),
            .I(N__25694));
    LocalMux I__6102 (
            .O(N__25710),
            .I(N__25694));
    InMux I__6101 (
            .O(N__25709),
            .I(N__25683));
    InMux I__6100 (
            .O(N__25708),
            .I(N__25680));
    Span4Mux_h I__6099 (
            .O(N__25705),
            .I(N__25677));
    Span4Mux_v I__6098 (
            .O(N__25694),
            .I(N__25674));
    InMux I__6097 (
            .O(N__25693),
            .I(N__25665));
    InMux I__6096 (
            .O(N__25692),
            .I(N__25665));
    InMux I__6095 (
            .O(N__25691),
            .I(N__25665));
    InMux I__6094 (
            .O(N__25690),
            .I(N__25665));
    InMux I__6093 (
            .O(N__25689),
            .I(N__25662));
    InMux I__6092 (
            .O(N__25688),
            .I(N__25659));
    InMux I__6091 (
            .O(N__25687),
            .I(N__25654));
    InMux I__6090 (
            .O(N__25686),
            .I(N__25654));
    LocalMux I__6089 (
            .O(N__25683),
            .I(un6_rowlto1));
    LocalMux I__6088 (
            .O(N__25680),
            .I(un6_rowlto1));
    Odrv4 I__6087 (
            .O(N__25677),
            .I(un6_rowlto1));
    Odrv4 I__6086 (
            .O(N__25674),
            .I(un6_rowlto1));
    LocalMux I__6085 (
            .O(N__25665),
            .I(un6_rowlto1));
    LocalMux I__6084 (
            .O(N__25662),
            .I(un6_rowlto1));
    LocalMux I__6083 (
            .O(N__25659),
            .I(un6_rowlto1));
    LocalMux I__6082 (
            .O(N__25654),
            .I(un6_rowlto1));
    CascadeMux I__6081 (
            .O(N__25637),
            .I(N__25634));
    InMux I__6080 (
            .O(N__25634),
            .I(N__25628));
    InMux I__6079 (
            .O(N__25633),
            .I(N__25628));
    LocalMux I__6078 (
            .O(N__25628),
            .I(ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0));
    CascadeMux I__6077 (
            .O(N__25625),
            .I(N__25622));
    InMux I__6076 (
            .O(N__25622),
            .I(N__25616));
    InMux I__6075 (
            .O(N__25621),
            .I(N__25616));
    LocalMux I__6074 (
            .O(N__25616),
            .I(N__25613));
    Span4Mux_s1_h I__6073 (
            .O(N__25613),
            .I(N__25610));
    Odrv4 I__6072 (
            .O(N__25610),
            .I(ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0));
    InMux I__6071 (
            .O(N__25607),
            .I(N__25604));
    LocalMux I__6070 (
            .O(N__25604),
            .I(ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0));
    CascadeMux I__6069 (
            .O(N__25601),
            .I(ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_));
    InMux I__6068 (
            .O(N__25598),
            .I(N__25595));
    LocalMux I__6067 (
            .O(N__25595),
            .I(ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0));
    InMux I__6066 (
            .O(N__25592),
            .I(N__25587));
    InMux I__6065 (
            .O(N__25591),
            .I(N__25580));
    InMux I__6064 (
            .O(N__25590),
            .I(N__25580));
    LocalMux I__6063 (
            .O(N__25587),
            .I(N__25577));
    InMux I__6062 (
            .O(N__25586),
            .I(N__25574));
    InMux I__6061 (
            .O(N__25585),
            .I(N__25571));
    LocalMux I__6060 (
            .O(N__25580),
            .I(N__25568));
    Span4Mux_v I__6059 (
            .O(N__25577),
            .I(N__25563));
    LocalMux I__6058 (
            .O(N__25574),
            .I(N__25563));
    LocalMux I__6057 (
            .O(N__25571),
            .I(N__25560));
    Span4Mux_h I__6056 (
            .O(N__25568),
            .I(N__25557));
    Span4Mux_h I__6055 (
            .O(N__25563),
            .I(N__25554));
    Odrv12 I__6054 (
            .O(N__25560),
            .I(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0));
    Odrv4 I__6053 (
            .O(N__25557),
            .I(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0));
    Odrv4 I__6052 (
            .O(N__25554),
            .I(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0));
    CascadeMux I__6051 (
            .O(N__25547),
            .I(N__25542));
    InMux I__6050 (
            .O(N__25546),
            .I(N__25535));
    InMux I__6049 (
            .O(N__25545),
            .I(N__25532));
    InMux I__6048 (
            .O(N__25542),
            .I(N__25529));
    InMux I__6047 (
            .O(N__25541),
            .I(N__25526));
    CascadeMux I__6046 (
            .O(N__25540),
            .I(N__25522));
    InMux I__6045 (
            .O(N__25539),
            .I(N__25519));
    CascadeMux I__6044 (
            .O(N__25538),
            .I(N__25514));
    LocalMux I__6043 (
            .O(N__25535),
            .I(N__25509));
    LocalMux I__6042 (
            .O(N__25532),
            .I(N__25506));
    LocalMux I__6041 (
            .O(N__25529),
            .I(N__25501));
    LocalMux I__6040 (
            .O(N__25526),
            .I(N__25501));
    InMux I__6039 (
            .O(N__25525),
            .I(N__25498));
    InMux I__6038 (
            .O(N__25522),
            .I(N__25495));
    LocalMux I__6037 (
            .O(N__25519),
            .I(N__25492));
    InMux I__6036 (
            .O(N__25518),
            .I(N__25489));
    CascadeMux I__6035 (
            .O(N__25517),
            .I(N__25486));
    InMux I__6034 (
            .O(N__25514),
            .I(N__25483));
    CascadeMux I__6033 (
            .O(N__25513),
            .I(N__25480));
    CascadeMux I__6032 (
            .O(N__25512),
            .I(N__25474));
    Span4Mux_v I__6031 (
            .O(N__25509),
            .I(N__25463));
    Span4Mux_h I__6030 (
            .O(N__25506),
            .I(N__25463));
    Span4Mux_v I__6029 (
            .O(N__25501),
            .I(N__25463));
    LocalMux I__6028 (
            .O(N__25498),
            .I(N__25463));
    LocalMux I__6027 (
            .O(N__25495),
            .I(N__25463));
    Span4Mux_v I__6026 (
            .O(N__25492),
            .I(N__25458));
    LocalMux I__6025 (
            .O(N__25489),
            .I(N__25458));
    InMux I__6024 (
            .O(N__25486),
            .I(N__25455));
    LocalMux I__6023 (
            .O(N__25483),
            .I(N__25452));
    InMux I__6022 (
            .O(N__25480),
            .I(N__25443));
    InMux I__6021 (
            .O(N__25479),
            .I(N__25443));
    InMux I__6020 (
            .O(N__25478),
            .I(N__25443));
    InMux I__6019 (
            .O(N__25477),
            .I(N__25443));
    InMux I__6018 (
            .O(N__25474),
            .I(N__25440));
    Span4Mux_h I__6017 (
            .O(N__25463),
            .I(N__25437));
    Span4Mux_h I__6016 (
            .O(N__25458),
            .I(N__25432));
    LocalMux I__6015 (
            .O(N__25455),
            .I(N__25432));
    Span12Mux_s11_h I__6014 (
            .O(N__25452),
            .I(N__25427));
    LocalMux I__6013 (
            .O(N__25443),
            .I(N__25427));
    LocalMux I__6012 (
            .O(N__25440),
            .I(un6_rowlto0));
    Odrv4 I__6011 (
            .O(N__25437),
            .I(un6_rowlto0));
    Odrv4 I__6010 (
            .O(N__25432),
            .I(un6_rowlto0));
    Odrv12 I__6009 (
            .O(N__25427),
            .I(un6_rowlto0));
    InMux I__6008 (
            .O(N__25418),
            .I(N__25410));
    InMux I__6007 (
            .O(N__25417),
            .I(N__25410));
    CascadeMux I__6006 (
            .O(N__25416),
            .I(N__25407));
    InMux I__6005 (
            .O(N__25415),
            .I(N__25391));
    LocalMux I__6004 (
            .O(N__25410),
            .I(N__25388));
    InMux I__6003 (
            .O(N__25407),
            .I(N__25383));
    InMux I__6002 (
            .O(N__25406),
            .I(N__25380));
    InMux I__6001 (
            .O(N__25405),
            .I(N__25373));
    InMux I__6000 (
            .O(N__25404),
            .I(N__25373));
    InMux I__5999 (
            .O(N__25403),
            .I(N__25373));
    InMux I__5998 (
            .O(N__25402),
            .I(N__25370));
    InMux I__5997 (
            .O(N__25401),
            .I(N__25365));
    InMux I__5996 (
            .O(N__25400),
            .I(N__25365));
    CascadeMux I__5995 (
            .O(N__25399),
            .I(N__25361));
    InMux I__5994 (
            .O(N__25398),
            .I(N__25357));
    InMux I__5993 (
            .O(N__25397),
            .I(N__25354));
    InMux I__5992 (
            .O(N__25396),
            .I(N__25351));
    InMux I__5991 (
            .O(N__25395),
            .I(N__25348));
    InMux I__5990 (
            .O(N__25394),
            .I(N__25345));
    LocalMux I__5989 (
            .O(N__25391),
            .I(N__25340));
    Span4Mux_v I__5988 (
            .O(N__25388),
            .I(N__25340));
    InMux I__5987 (
            .O(N__25387),
            .I(N__25337));
    InMux I__5986 (
            .O(N__25386),
            .I(N__25334));
    LocalMux I__5985 (
            .O(N__25383),
            .I(N__25327));
    LocalMux I__5984 (
            .O(N__25380),
            .I(N__25327));
    LocalMux I__5983 (
            .O(N__25373),
            .I(N__25327));
    LocalMux I__5982 (
            .O(N__25370),
            .I(N__25322));
    LocalMux I__5981 (
            .O(N__25365),
            .I(N__25322));
    InMux I__5980 (
            .O(N__25364),
            .I(N__25314));
    InMux I__5979 (
            .O(N__25361),
            .I(N__25314));
    InMux I__5978 (
            .O(N__25360),
            .I(N__25314));
    LocalMux I__5977 (
            .O(N__25357),
            .I(N__25311));
    LocalMux I__5976 (
            .O(N__25354),
            .I(N__25307));
    LocalMux I__5975 (
            .O(N__25351),
            .I(N__25292));
    LocalMux I__5974 (
            .O(N__25348),
            .I(N__25292));
    LocalMux I__5973 (
            .O(N__25345),
            .I(N__25292));
    Span4Mux_h I__5972 (
            .O(N__25340),
            .I(N__25292));
    LocalMux I__5971 (
            .O(N__25337),
            .I(N__25292));
    LocalMux I__5970 (
            .O(N__25334),
            .I(N__25292));
    Span4Mux_v I__5969 (
            .O(N__25327),
            .I(N__25292));
    Span4Mux_v I__5968 (
            .O(N__25322),
            .I(N__25289));
    InMux I__5967 (
            .O(N__25321),
            .I(N__25286));
    LocalMux I__5966 (
            .O(N__25314),
            .I(N__25280));
    Span4Mux_h I__5965 (
            .O(N__25311),
            .I(N__25280));
    InMux I__5964 (
            .O(N__25310),
            .I(N__25277));
    Span4Mux_v I__5963 (
            .O(N__25307),
            .I(N__25268));
    Span4Mux_v I__5962 (
            .O(N__25292),
            .I(N__25268));
    Span4Mux_s0_h I__5961 (
            .O(N__25289),
            .I(N__25268));
    LocalMux I__5960 (
            .O(N__25286),
            .I(N__25268));
    InMux I__5959 (
            .O(N__25285),
            .I(N__25265));
    Odrv4 I__5958 (
            .O(N__25280),
            .I(column_1_i_2));
    LocalMux I__5957 (
            .O(N__25277),
            .I(column_1_i_2));
    Odrv4 I__5956 (
            .O(N__25268),
            .I(column_1_i_2));
    LocalMux I__5955 (
            .O(N__25265),
            .I(column_1_i_2));
    CascadeMux I__5954 (
            .O(N__25256),
            .I(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_));
    InMux I__5953 (
            .O(N__25253),
            .I(N__25250));
    LocalMux I__5952 (
            .O(N__25250),
            .I(N__25247));
    Span4Mux_s3_h I__5951 (
            .O(N__25247),
            .I(N__25243));
    InMux I__5950 (
            .O(N__25246),
            .I(N__25240));
    Odrv4 I__5949 (
            .O(N__25243),
            .I(ScreenBuffer_0_7_RNIN5F98I1Z0Z_0));
    LocalMux I__5948 (
            .O(N__25240),
            .I(ScreenBuffer_0_7_RNIN5F98I1Z0Z_0));
    InMux I__5947 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__5946 (
            .O(N__25232),
            .I(un115_pixel_5_am_sx_1));
    CascadeMux I__5945 (
            .O(N__25229),
            .I(un113_pixel_3_0_11__N_16_cascade_));
    InMux I__5944 (
            .O(N__25226),
            .I(N__25221));
    InMux I__5943 (
            .O(N__25225),
            .I(N__25218));
    InMux I__5942 (
            .O(N__25224),
            .I(N__25215));
    LocalMux I__5941 (
            .O(N__25221),
            .I(N__25208));
    LocalMux I__5940 (
            .O(N__25218),
            .I(N__25202));
    LocalMux I__5939 (
            .O(N__25215),
            .I(N__25199));
    InMux I__5938 (
            .O(N__25214),
            .I(N__25196));
    InMux I__5937 (
            .O(N__25213),
            .I(N__25191));
    InMux I__5936 (
            .O(N__25212),
            .I(N__25191));
    InMux I__5935 (
            .O(N__25211),
            .I(N__25188));
    Span4Mux_s3_h I__5934 (
            .O(N__25208),
            .I(N__25185));
    InMux I__5933 (
            .O(N__25207),
            .I(N__25182));
    InMux I__5932 (
            .O(N__25206),
            .I(N__25177));
    InMux I__5931 (
            .O(N__25205),
            .I(N__25177));
    Span4Mux_v I__5930 (
            .O(N__25202),
            .I(N__25168));
    Span4Mux_s3_h I__5929 (
            .O(N__25199),
            .I(N__25168));
    LocalMux I__5928 (
            .O(N__25196),
            .I(N__25168));
    LocalMux I__5927 (
            .O(N__25191),
            .I(N__25168));
    LocalMux I__5926 (
            .O(N__25188),
            .I(un113_pixel_7_1_7__N_11));
    Odrv4 I__5925 (
            .O(N__25185),
            .I(un113_pixel_7_1_7__N_11));
    LocalMux I__5924 (
            .O(N__25182),
            .I(un113_pixel_7_1_7__N_11));
    LocalMux I__5923 (
            .O(N__25177),
            .I(un113_pixel_7_1_7__N_11));
    Odrv4 I__5922 (
            .O(N__25168),
            .I(un113_pixel_7_1_7__N_11));
    InMux I__5921 (
            .O(N__25157),
            .I(N__25154));
    LocalMux I__5920 (
            .O(N__25154),
            .I(N_4573_0));
    InMux I__5919 (
            .O(N__25151),
            .I(N__25146));
    InMux I__5918 (
            .O(N__25150),
            .I(N__25142));
    InMux I__5917 (
            .O(N__25149),
            .I(N__25137));
    LocalMux I__5916 (
            .O(N__25146),
            .I(N__25130));
    InMux I__5915 (
            .O(N__25145),
            .I(N__25127));
    LocalMux I__5914 (
            .O(N__25142),
            .I(N__25124));
    InMux I__5913 (
            .O(N__25141),
            .I(N__25119));
    InMux I__5912 (
            .O(N__25140),
            .I(N__25119));
    LocalMux I__5911 (
            .O(N__25137),
            .I(N__25116));
    InMux I__5910 (
            .O(N__25136),
            .I(N__25113));
    InMux I__5909 (
            .O(N__25135),
            .I(N__25110));
    InMux I__5908 (
            .O(N__25134),
            .I(N__25105));
    InMux I__5907 (
            .O(N__25133),
            .I(N__25105));
    Span4Mux_h I__5906 (
            .O(N__25130),
            .I(N__25098));
    LocalMux I__5905 (
            .O(N__25127),
            .I(N__25098));
    Span4Mux_h I__5904 (
            .O(N__25124),
            .I(N__25098));
    LocalMux I__5903 (
            .O(N__25119),
            .I(N__25095));
    Odrv12 I__5902 (
            .O(N__25116),
            .I(un112_pixel_2_2));
    LocalMux I__5901 (
            .O(N__25113),
            .I(un112_pixel_2_2));
    LocalMux I__5900 (
            .O(N__25110),
            .I(un112_pixel_2_2));
    LocalMux I__5899 (
            .O(N__25105),
            .I(un112_pixel_2_2));
    Odrv4 I__5898 (
            .O(N__25098),
            .I(un112_pixel_2_2));
    Odrv4 I__5897 (
            .O(N__25095),
            .I(un112_pixel_2_2));
    CascadeMux I__5896 (
            .O(N__25082),
            .I(N__25071));
    InMux I__5895 (
            .O(N__25081),
            .I(N__25059));
    InMux I__5894 (
            .O(N__25080),
            .I(N__25059));
    InMux I__5893 (
            .O(N__25079),
            .I(N__25053));
    InMux I__5892 (
            .O(N__25078),
            .I(N__25050));
    InMux I__5891 (
            .O(N__25077),
            .I(N__25043));
    InMux I__5890 (
            .O(N__25076),
            .I(N__25043));
    InMux I__5889 (
            .O(N__25075),
            .I(N__25043));
    InMux I__5888 (
            .O(N__25074),
            .I(N__25037));
    InMux I__5887 (
            .O(N__25071),
            .I(N__25037));
    InMux I__5886 (
            .O(N__25070),
            .I(N__25032));
    CascadeMux I__5885 (
            .O(N__25069),
            .I(N__25022));
    CascadeMux I__5884 (
            .O(N__25068),
            .I(N__25008));
    InMux I__5883 (
            .O(N__25067),
            .I(N__24997));
    InMux I__5882 (
            .O(N__25066),
            .I(N__24997));
    InMux I__5881 (
            .O(N__25065),
            .I(N__24997));
    InMux I__5880 (
            .O(N__25064),
            .I(N__24997));
    LocalMux I__5879 (
            .O(N__25059),
            .I(N__24992));
    InMux I__5878 (
            .O(N__25058),
            .I(N__24985));
    InMux I__5877 (
            .O(N__25057),
            .I(N__24985));
    InMux I__5876 (
            .O(N__25056),
            .I(N__24985));
    LocalMux I__5875 (
            .O(N__25053),
            .I(N__24978));
    LocalMux I__5874 (
            .O(N__25050),
            .I(N__24978));
    LocalMux I__5873 (
            .O(N__25043),
            .I(N__24978));
    InMux I__5872 (
            .O(N__25042),
            .I(N__24975));
    LocalMux I__5871 (
            .O(N__25037),
            .I(N__24972));
    InMux I__5870 (
            .O(N__25036),
            .I(N__24967));
    InMux I__5869 (
            .O(N__25035),
            .I(N__24967));
    LocalMux I__5868 (
            .O(N__25032),
            .I(N__24964));
    InMux I__5867 (
            .O(N__25031),
            .I(N__24959));
    InMux I__5866 (
            .O(N__25030),
            .I(N__24959));
    InMux I__5865 (
            .O(N__25029),
            .I(N__24954));
    InMux I__5864 (
            .O(N__25028),
            .I(N__24954));
    InMux I__5863 (
            .O(N__25027),
            .I(N__24949));
    InMux I__5862 (
            .O(N__25026),
            .I(N__24949));
    InMux I__5861 (
            .O(N__25025),
            .I(N__24938));
    InMux I__5860 (
            .O(N__25022),
            .I(N__24938));
    InMux I__5859 (
            .O(N__25021),
            .I(N__24938));
    InMux I__5858 (
            .O(N__25020),
            .I(N__24938));
    InMux I__5857 (
            .O(N__25019),
            .I(N__24938));
    InMux I__5856 (
            .O(N__25018),
            .I(N__24929));
    InMux I__5855 (
            .O(N__25017),
            .I(N__24929));
    InMux I__5854 (
            .O(N__25016),
            .I(N__24929));
    InMux I__5853 (
            .O(N__25015),
            .I(N__24929));
    InMux I__5852 (
            .O(N__25014),
            .I(N__24920));
    InMux I__5851 (
            .O(N__25013),
            .I(N__24920));
    InMux I__5850 (
            .O(N__25012),
            .I(N__24920));
    InMux I__5849 (
            .O(N__25011),
            .I(N__24920));
    InMux I__5848 (
            .O(N__25008),
            .I(N__24915));
    InMux I__5847 (
            .O(N__25007),
            .I(N__24915));
    InMux I__5846 (
            .O(N__25006),
            .I(N__24912));
    LocalMux I__5845 (
            .O(N__24997),
            .I(N__24909));
    InMux I__5844 (
            .O(N__24996),
            .I(N__24904));
    InMux I__5843 (
            .O(N__24995),
            .I(N__24904));
    Span4Mux_v I__5842 (
            .O(N__24992),
            .I(N__24897));
    LocalMux I__5841 (
            .O(N__24985),
            .I(N__24897));
    Span4Mux_v I__5840 (
            .O(N__24978),
            .I(N__24897));
    LocalMux I__5839 (
            .O(N__24975),
            .I(N__24890));
    Span4Mux_s3_v I__5838 (
            .O(N__24972),
            .I(N__24890));
    LocalMux I__5837 (
            .O(N__24967),
            .I(N__24890));
    Odrv4 I__5836 (
            .O(N__24964),
            .I(currentchar_1_1));
    LocalMux I__5835 (
            .O(N__24959),
            .I(currentchar_1_1));
    LocalMux I__5834 (
            .O(N__24954),
            .I(currentchar_1_1));
    LocalMux I__5833 (
            .O(N__24949),
            .I(currentchar_1_1));
    LocalMux I__5832 (
            .O(N__24938),
            .I(currentchar_1_1));
    LocalMux I__5831 (
            .O(N__24929),
            .I(currentchar_1_1));
    LocalMux I__5830 (
            .O(N__24920),
            .I(currentchar_1_1));
    LocalMux I__5829 (
            .O(N__24915),
            .I(currentchar_1_1));
    LocalMux I__5828 (
            .O(N__24912),
            .I(currentchar_1_1));
    Odrv4 I__5827 (
            .O(N__24909),
            .I(currentchar_1_1));
    LocalMux I__5826 (
            .O(N__24904),
            .I(currentchar_1_1));
    Odrv4 I__5825 (
            .O(N__24897),
            .I(currentchar_1_1));
    Odrv4 I__5824 (
            .O(N__24890),
            .I(currentchar_1_1));
    CascadeMux I__5823 (
            .O(N__24863),
            .I(N__24849));
    CascadeMux I__5822 (
            .O(N__24862),
            .I(N__24846));
    CascadeMux I__5821 (
            .O(N__24861),
            .I(N__24843));
    CascadeMux I__5820 (
            .O(N__24860),
            .I(N__24840));
    CascadeMux I__5819 (
            .O(N__24859),
            .I(N__24829));
    CascadeMux I__5818 (
            .O(N__24858),
            .I(N__24822));
    CascadeMux I__5817 (
            .O(N__24857),
            .I(N__24818));
    CascadeMux I__5816 (
            .O(N__24856),
            .I(N__24813));
    CascadeMux I__5815 (
            .O(N__24855),
            .I(N__24810));
    CascadeMux I__5814 (
            .O(N__24854),
            .I(N__24805));
    CascadeMux I__5813 (
            .O(N__24853),
            .I(N__24801));
    CascadeMux I__5812 (
            .O(N__24852),
            .I(N__24797));
    InMux I__5811 (
            .O(N__24849),
            .I(N__24794));
    InMux I__5810 (
            .O(N__24846),
            .I(N__24791));
    InMux I__5809 (
            .O(N__24843),
            .I(N__24786));
    InMux I__5808 (
            .O(N__24840),
            .I(N__24786));
    InMux I__5807 (
            .O(N__24839),
            .I(N__24781));
    InMux I__5806 (
            .O(N__24838),
            .I(N__24781));
    InMux I__5805 (
            .O(N__24837),
            .I(N__24778));
    InMux I__5804 (
            .O(N__24836),
            .I(N__24773));
    InMux I__5803 (
            .O(N__24835),
            .I(N__24770));
    InMux I__5802 (
            .O(N__24834),
            .I(N__24767));
    CascadeMux I__5801 (
            .O(N__24833),
            .I(N__24764));
    CascadeMux I__5800 (
            .O(N__24832),
            .I(N__24761));
    InMux I__5799 (
            .O(N__24829),
            .I(N__24756));
    InMux I__5798 (
            .O(N__24828),
            .I(N__24753));
    CascadeMux I__5797 (
            .O(N__24827),
            .I(N__24749));
    InMux I__5796 (
            .O(N__24826),
            .I(N__24743));
    InMux I__5795 (
            .O(N__24825),
            .I(N__24743));
    InMux I__5794 (
            .O(N__24822),
            .I(N__24734));
    InMux I__5793 (
            .O(N__24821),
            .I(N__24734));
    InMux I__5792 (
            .O(N__24818),
            .I(N__24734));
    InMux I__5791 (
            .O(N__24817),
            .I(N__24734));
    InMux I__5790 (
            .O(N__24816),
            .I(N__24729));
    InMux I__5789 (
            .O(N__24813),
            .I(N__24729));
    InMux I__5788 (
            .O(N__24810),
            .I(N__24726));
    InMux I__5787 (
            .O(N__24809),
            .I(N__24718));
    InMux I__5786 (
            .O(N__24808),
            .I(N__24718));
    InMux I__5785 (
            .O(N__24805),
            .I(N__24718));
    CascadeMux I__5784 (
            .O(N__24804),
            .I(N__24715));
    InMux I__5783 (
            .O(N__24801),
            .I(N__24712));
    InMux I__5782 (
            .O(N__24800),
            .I(N__24707));
    InMux I__5781 (
            .O(N__24797),
            .I(N__24707));
    LocalMux I__5780 (
            .O(N__24794),
            .I(N__24704));
    LocalMux I__5779 (
            .O(N__24791),
            .I(N__24695));
    LocalMux I__5778 (
            .O(N__24786),
            .I(N__24695));
    LocalMux I__5777 (
            .O(N__24781),
            .I(N__24695));
    LocalMux I__5776 (
            .O(N__24778),
            .I(N__24695));
    InMux I__5775 (
            .O(N__24777),
            .I(N__24690));
    InMux I__5774 (
            .O(N__24776),
            .I(N__24690));
    LocalMux I__5773 (
            .O(N__24773),
            .I(N__24683));
    LocalMux I__5772 (
            .O(N__24770),
            .I(N__24683));
    LocalMux I__5771 (
            .O(N__24767),
            .I(N__24683));
    InMux I__5770 (
            .O(N__24764),
            .I(N__24678));
    InMux I__5769 (
            .O(N__24761),
            .I(N__24678));
    InMux I__5768 (
            .O(N__24760),
            .I(N__24673));
    InMux I__5767 (
            .O(N__24759),
            .I(N__24673));
    LocalMux I__5766 (
            .O(N__24756),
            .I(N__24670));
    LocalMux I__5765 (
            .O(N__24753),
            .I(N__24667));
    InMux I__5764 (
            .O(N__24752),
            .I(N__24664));
    InMux I__5763 (
            .O(N__24749),
            .I(N__24659));
    InMux I__5762 (
            .O(N__24748),
            .I(N__24659));
    LocalMux I__5761 (
            .O(N__24743),
            .I(N__24656));
    LocalMux I__5760 (
            .O(N__24734),
            .I(N__24649));
    LocalMux I__5759 (
            .O(N__24729),
            .I(N__24649));
    LocalMux I__5758 (
            .O(N__24726),
            .I(N__24649));
    InMux I__5757 (
            .O(N__24725),
            .I(N__24646));
    LocalMux I__5756 (
            .O(N__24718),
            .I(N__24643));
    InMux I__5755 (
            .O(N__24715),
            .I(N__24640));
    LocalMux I__5754 (
            .O(N__24712),
            .I(N__24636));
    LocalMux I__5753 (
            .O(N__24707),
            .I(N__24629));
    Span4Mux_h I__5752 (
            .O(N__24704),
            .I(N__24629));
    Span4Mux_s3_v I__5751 (
            .O(N__24695),
            .I(N__24629));
    LocalMux I__5750 (
            .O(N__24690),
            .I(N__24622));
    Span4Mux_v I__5749 (
            .O(N__24683),
            .I(N__24622));
    LocalMux I__5748 (
            .O(N__24678),
            .I(N__24622));
    LocalMux I__5747 (
            .O(N__24673),
            .I(N__24619));
    Span4Mux_v I__5746 (
            .O(N__24670),
            .I(N__24616));
    Span4Mux_v I__5745 (
            .O(N__24667),
            .I(N__24613));
    LocalMux I__5744 (
            .O(N__24664),
            .I(N__24598));
    LocalMux I__5743 (
            .O(N__24659),
            .I(N__24598));
    Span4Mux_v I__5742 (
            .O(N__24656),
            .I(N__24598));
    Span4Mux_v I__5741 (
            .O(N__24649),
            .I(N__24598));
    LocalMux I__5740 (
            .O(N__24646),
            .I(N__24598));
    Span4Mux_s2_h I__5739 (
            .O(N__24643),
            .I(N__24598));
    LocalMux I__5738 (
            .O(N__24640),
            .I(N__24598));
    CascadeMux I__5737 (
            .O(N__24639),
            .I(N__24595));
    Span4Mux_h I__5736 (
            .O(N__24636),
            .I(N__24588));
    Span4Mux_v I__5735 (
            .O(N__24629),
            .I(N__24588));
    Span4Mux_h I__5734 (
            .O(N__24622),
            .I(N__24583));
    Span4Mux_v I__5733 (
            .O(N__24619),
            .I(N__24583));
    Span4Mux_s1_h I__5732 (
            .O(N__24616),
            .I(N__24580));
    Span4Mux_v I__5731 (
            .O(N__24613),
            .I(N__24575));
    Span4Mux_v I__5730 (
            .O(N__24598),
            .I(N__24575));
    InMux I__5729 (
            .O(N__24595),
            .I(N__24572));
    InMux I__5728 (
            .O(N__24594),
            .I(N__24567));
    InMux I__5727 (
            .O(N__24593),
            .I(N__24567));
    Span4Mux_v I__5726 (
            .O(N__24588),
            .I(N__24564));
    Span4Mux_v I__5725 (
            .O(N__24583),
            .I(N__24561));
    Span4Mux_h I__5724 (
            .O(N__24580),
            .I(N__24556));
    Span4Mux_h I__5723 (
            .O(N__24575),
            .I(N__24556));
    LocalMux I__5722 (
            .O(N__24572),
            .I(beamYZ0Z_0));
    LocalMux I__5721 (
            .O(N__24567),
            .I(beamYZ0Z_0));
    Odrv4 I__5720 (
            .O(N__24564),
            .I(beamYZ0Z_0));
    Odrv4 I__5719 (
            .O(N__24561),
            .I(beamYZ0Z_0));
    Odrv4 I__5718 (
            .O(N__24556),
            .I(beamYZ0Z_0));
    InMux I__5717 (
            .O(N__24545),
            .I(N__24537));
    InMux I__5716 (
            .O(N__24544),
            .I(N__24532));
    InMux I__5715 (
            .O(N__24543),
            .I(N__24529));
    InMux I__5714 (
            .O(N__24542),
            .I(N__24526));
    InMux I__5713 (
            .O(N__24541),
            .I(N__24521));
    InMux I__5712 (
            .O(N__24540),
            .I(N__24518));
    LocalMux I__5711 (
            .O(N__24537),
            .I(N__24515));
    InMux I__5710 (
            .O(N__24536),
            .I(N__24499));
    InMux I__5709 (
            .O(N__24535),
            .I(N__24499));
    LocalMux I__5708 (
            .O(N__24532),
            .I(N__24496));
    LocalMux I__5707 (
            .O(N__24529),
            .I(N__24493));
    LocalMux I__5706 (
            .O(N__24526),
            .I(N__24490));
    InMux I__5705 (
            .O(N__24525),
            .I(N__24485));
    InMux I__5704 (
            .O(N__24524),
            .I(N__24485));
    LocalMux I__5703 (
            .O(N__24521),
            .I(N__24468));
    LocalMux I__5702 (
            .O(N__24518),
            .I(N__24463));
    Span4Mux_s3_h I__5701 (
            .O(N__24515),
            .I(N__24463));
    InMux I__5700 (
            .O(N__24514),
            .I(N__24458));
    InMux I__5699 (
            .O(N__24513),
            .I(N__24458));
    InMux I__5698 (
            .O(N__24512),
            .I(N__24451));
    InMux I__5697 (
            .O(N__24511),
            .I(N__24451));
    InMux I__5696 (
            .O(N__24510),
            .I(N__24451));
    InMux I__5695 (
            .O(N__24509),
            .I(N__24440));
    InMux I__5694 (
            .O(N__24508),
            .I(N__24440));
    InMux I__5693 (
            .O(N__24507),
            .I(N__24440));
    InMux I__5692 (
            .O(N__24506),
            .I(N__24440));
    InMux I__5691 (
            .O(N__24505),
            .I(N__24440));
    InMux I__5690 (
            .O(N__24504),
            .I(N__24437));
    LocalMux I__5689 (
            .O(N__24499),
            .I(N__24432));
    Span4Mux_s3_h I__5688 (
            .O(N__24496),
            .I(N__24432));
    Span4Mux_h I__5687 (
            .O(N__24493),
            .I(N__24425));
    Span4Mux_v I__5686 (
            .O(N__24490),
            .I(N__24425));
    LocalMux I__5685 (
            .O(N__24485),
            .I(N__24425));
    InMux I__5684 (
            .O(N__24484),
            .I(N__24420));
    InMux I__5683 (
            .O(N__24483),
            .I(N__24420));
    InMux I__5682 (
            .O(N__24482),
            .I(N__24413));
    InMux I__5681 (
            .O(N__24481),
            .I(N__24413));
    InMux I__5680 (
            .O(N__24480),
            .I(N__24413));
    InMux I__5679 (
            .O(N__24479),
            .I(N__24404));
    InMux I__5678 (
            .O(N__24478),
            .I(N__24404));
    InMux I__5677 (
            .O(N__24477),
            .I(N__24404));
    InMux I__5676 (
            .O(N__24476),
            .I(N__24404));
    InMux I__5675 (
            .O(N__24475),
            .I(N__24393));
    InMux I__5674 (
            .O(N__24474),
            .I(N__24393));
    InMux I__5673 (
            .O(N__24473),
            .I(N__24393));
    InMux I__5672 (
            .O(N__24472),
            .I(N__24393));
    InMux I__5671 (
            .O(N__24471),
            .I(N__24393));
    Odrv12 I__5670 (
            .O(N__24468),
            .I(currentchar_1_0));
    Odrv4 I__5669 (
            .O(N__24463),
            .I(currentchar_1_0));
    LocalMux I__5668 (
            .O(N__24458),
            .I(currentchar_1_0));
    LocalMux I__5667 (
            .O(N__24451),
            .I(currentchar_1_0));
    LocalMux I__5666 (
            .O(N__24440),
            .I(currentchar_1_0));
    LocalMux I__5665 (
            .O(N__24437),
            .I(currentchar_1_0));
    Odrv4 I__5664 (
            .O(N__24432),
            .I(currentchar_1_0));
    Odrv4 I__5663 (
            .O(N__24425),
            .I(currentchar_1_0));
    LocalMux I__5662 (
            .O(N__24420),
            .I(currentchar_1_0));
    LocalMux I__5661 (
            .O(N__24413),
            .I(currentchar_1_0));
    LocalMux I__5660 (
            .O(N__24404),
            .I(currentchar_1_0));
    LocalMux I__5659 (
            .O(N__24393),
            .I(currentchar_1_0));
    InMux I__5658 (
            .O(N__24368),
            .I(N__24365));
    LocalMux I__5657 (
            .O(N__24365),
            .I(un115_pixel_3_am_2));
    InMux I__5656 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__5655 (
            .O(N__24359),
            .I(N__24355));
    CascadeMux I__5654 (
            .O(N__24358),
            .I(N__24350));
    Span4Mux_s0_h I__5653 (
            .O(N__24355),
            .I(N__24344));
    InMux I__5652 (
            .O(N__24354),
            .I(N__24333));
    InMux I__5651 (
            .O(N__24353),
            .I(N__24333));
    InMux I__5650 (
            .O(N__24350),
            .I(N__24333));
    InMux I__5649 (
            .O(N__24349),
            .I(N__24333));
    InMux I__5648 (
            .O(N__24348),
            .I(N__24333));
    CascadeMux I__5647 (
            .O(N__24347),
            .I(N__24330));
    Span4Mux_h I__5646 (
            .O(N__24344),
            .I(N__24325));
    LocalMux I__5645 (
            .O(N__24333),
            .I(N__24325));
    InMux I__5644 (
            .O(N__24330),
            .I(N__24322));
    Sp12to4 I__5643 (
            .O(N__24325),
            .I(N__24317));
    LocalMux I__5642 (
            .O(N__24322),
            .I(N__24317));
    Odrv12 I__5641 (
            .O(N__24317),
            .I(charx_if_generate_plus_mult1_un75_sum));
    CascadeMux I__5640 (
            .O(N__24314),
            .I(N__24311));
    InMux I__5639 (
            .O(N__24311),
            .I(N__24308));
    LocalMux I__5638 (
            .O(N__24308),
            .I(column_1_if_generate_plus_mult1_un75_sum_iZ0));
    InMux I__5637 (
            .O(N__24305),
            .I(N__24302));
    LocalMux I__5636 (
            .O(N__24302),
            .I(G_673));
    CascadeMux I__5635 (
            .O(N__24299),
            .I(N__24296));
    InMux I__5634 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__5633 (
            .O(N__24293),
            .I(if_generate_plus_mult1_un75_sum_cry_2_s));
    CascadeMux I__5632 (
            .O(N__24290),
            .I(N__24287));
    InMux I__5631 (
            .O(N__24287),
            .I(N__24284));
    LocalMux I__5630 (
            .O(N__24284),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__5629 (
            .O(N__24281),
            .I(N__24278));
    LocalMux I__5628 (
            .O(N__24278),
            .I(G_674));
    InMux I__5627 (
            .O(N__24275),
            .I(N__24272));
    LocalMux I__5626 (
            .O(N__24272),
            .I(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__5625 (
            .O(N__24269),
            .I(column_1_if_generate_plus_mult1_un82_sum_cry_4));
    InMux I__5624 (
            .O(N__24266),
            .I(N__24263));
    LocalMux I__5623 (
            .O(N__24263),
            .I(N_1303_0));
    CascadeMux I__5622 (
            .O(N__24260),
            .I(g0_16_x0_cascade_));
    InMux I__5621 (
            .O(N__24257),
            .I(N__24254));
    LocalMux I__5620 (
            .O(N__24254),
            .I(g0_16_x1));
    InMux I__5619 (
            .O(N__24251),
            .I(N__24248));
    LocalMux I__5618 (
            .O(N__24248),
            .I(N__24245));
    Odrv4 I__5617 (
            .O(N__24245),
            .I(N_4560_0));
    InMux I__5616 (
            .O(N__24242),
            .I(N__24239));
    LocalMux I__5615 (
            .O(N__24239),
            .I(N__24236));
    Span4Mux_h I__5614 (
            .O(N__24236),
            .I(N__24233));
    Odrv4 I__5613 (
            .O(N__24233),
            .I(N_1309_0));
    InMux I__5612 (
            .O(N__24230),
            .I(N__24226));
    InMux I__5611 (
            .O(N__24229),
            .I(N__24223));
    LocalMux I__5610 (
            .O(N__24226),
            .I(N__24220));
    LocalMux I__5609 (
            .O(N__24223),
            .I(N__24217));
    Odrv4 I__5608 (
            .O(N__24220),
            .I(un113_pixel_4_0_15__N_2));
    Odrv4 I__5607 (
            .O(N__24217),
            .I(un113_pixel_4_0_15__N_2));
    InMux I__5606 (
            .O(N__24212),
            .I(N__24209));
    LocalMux I__5605 (
            .O(N__24209),
            .I(N__24206));
    Span4Mux_s3_h I__5604 (
            .O(N__24206),
            .I(N__24203));
    Odrv4 I__5603 (
            .O(N__24203),
            .I(un113_pixel_7_1_7__N_9));
    CascadeMux I__5602 (
            .O(N__24200),
            .I(beamY_RNIJIDRG11Z0Z_0_cascade_));
    InMux I__5601 (
            .O(N__24197),
            .I(N__24194));
    LocalMux I__5600 (
            .O(N__24194),
            .I(N__24191));
    Span4Mux_s2_h I__5599 (
            .O(N__24191),
            .I(N__24188));
    Odrv4 I__5598 (
            .O(N__24188),
            .I(beamY_RNIJIDRG11_0Z0Z_0));
    CascadeMux I__5597 (
            .O(N__24185),
            .I(beamY_RNIRG0LHO1Z0Z_0_cascade_));
    InMux I__5596 (
            .O(N__24182),
            .I(N__24176));
    InMux I__5595 (
            .O(N__24181),
            .I(N__24176));
    LocalMux I__5594 (
            .O(N__24176),
            .I(N__24173));
    Odrv4 I__5593 (
            .O(N__24173),
            .I(ScreenBuffer_0_7_RNIB3R6U63Z0Z_0));
    InMux I__5592 (
            .O(N__24170),
            .I(N__24163));
    InMux I__5591 (
            .O(N__24169),
            .I(N__24163));
    InMux I__5590 (
            .O(N__24168),
            .I(N__24155));
    LocalMux I__5589 (
            .O(N__24163),
            .I(N__24150));
    CascadeMux I__5588 (
            .O(N__24162),
            .I(N__24147));
    InMux I__5587 (
            .O(N__24161),
            .I(N__24139));
    InMux I__5586 (
            .O(N__24160),
            .I(N__24139));
    InMux I__5585 (
            .O(N__24159),
            .I(N__24139));
    CascadeMux I__5584 (
            .O(N__24158),
            .I(N__24132));
    LocalMux I__5583 (
            .O(N__24155),
            .I(N__24127));
    InMux I__5582 (
            .O(N__24154),
            .I(N__24124));
    InMux I__5581 (
            .O(N__24153),
            .I(N__24121));
    Span4Mux_s2_v I__5580 (
            .O(N__24150),
            .I(N__24118));
    InMux I__5579 (
            .O(N__24147),
            .I(N__24114));
    InMux I__5578 (
            .O(N__24146),
            .I(N__24111));
    LocalMux I__5577 (
            .O(N__24139),
            .I(N__24108));
    InMux I__5576 (
            .O(N__24138),
            .I(N__24105));
    InMux I__5575 (
            .O(N__24137),
            .I(N__24100));
    InMux I__5574 (
            .O(N__24136),
            .I(N__24100));
    InMux I__5573 (
            .O(N__24135),
            .I(N__24093));
    InMux I__5572 (
            .O(N__24132),
            .I(N__24093));
    InMux I__5571 (
            .O(N__24131),
            .I(N__24093));
    InMux I__5570 (
            .O(N__24130),
            .I(N__24090));
    Span4Mux_v I__5569 (
            .O(N__24127),
            .I(N__24081));
    LocalMux I__5568 (
            .O(N__24124),
            .I(N__24081));
    LocalMux I__5567 (
            .O(N__24121),
            .I(N__24081));
    Span4Mux_h I__5566 (
            .O(N__24118),
            .I(N__24081));
    InMux I__5565 (
            .O(N__24117),
            .I(N__24078));
    LocalMux I__5564 (
            .O(N__24114),
            .I(N__24071));
    LocalMux I__5563 (
            .O(N__24111),
            .I(N__24071));
    Span4Mux_s3_v I__5562 (
            .O(N__24108),
            .I(N__24071));
    LocalMux I__5561 (
            .O(N__24105),
            .I(N__24068));
    LocalMux I__5560 (
            .O(N__24100),
            .I(N__24063));
    LocalMux I__5559 (
            .O(N__24093),
            .I(N__24063));
    LocalMux I__5558 (
            .O(N__24090),
            .I(N__24060));
    Span4Mux_v I__5557 (
            .O(N__24081),
            .I(N__24057));
    LocalMux I__5556 (
            .O(N__24078),
            .I(N__24052));
    Span4Mux_v I__5555 (
            .O(N__24071),
            .I(N__24052));
    Span4Mux_v I__5554 (
            .O(N__24068),
            .I(N__24049));
    Span4Mux_v I__5553 (
            .O(N__24063),
            .I(N__24046));
    Odrv12 I__5552 (
            .O(N__24060),
            .I(font_un28_pixel_29));
    Odrv4 I__5551 (
            .O(N__24057),
            .I(font_un28_pixel_29));
    Odrv4 I__5550 (
            .O(N__24052),
            .I(font_un28_pixel_29));
    Odrv4 I__5549 (
            .O(N__24049),
            .I(font_un28_pixel_29));
    Odrv4 I__5548 (
            .O(N__24046),
            .I(font_un28_pixel_29));
    InMux I__5547 (
            .O(N__24035),
            .I(N__24032));
    LocalMux I__5546 (
            .O(N__24032),
            .I(beamY_RNIRG0LHO1Z0Z_0));
    InMux I__5545 (
            .O(N__24029),
            .I(N__24026));
    LocalMux I__5544 (
            .O(N__24026),
            .I(N__24023));
    Odrv12 I__5543 (
            .O(N__24023),
            .I(ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0));
    CascadeMux I__5542 (
            .O(N__24020),
            .I(g0_2_x1_cascade_));
    InMux I__5541 (
            .O(N__24017),
            .I(N__24014));
    LocalMux I__5540 (
            .O(N__24014),
            .I(g0_2_x0));
    InMux I__5539 (
            .O(N__24011),
            .I(N__24005));
    InMux I__5538 (
            .O(N__24010),
            .I(N__24005));
    LocalMux I__5537 (
            .O(N__24005),
            .I(N_1331_0));
    InMux I__5536 (
            .O(N__24002),
            .I(N__23995));
    InMux I__5535 (
            .O(N__24001),
            .I(N__23991));
    InMux I__5534 (
            .O(N__24000),
            .I(N__23988));
    InMux I__5533 (
            .O(N__23999),
            .I(N__23982));
    InMux I__5532 (
            .O(N__23998),
            .I(N__23982));
    LocalMux I__5531 (
            .O(N__23995),
            .I(N__23979));
    InMux I__5530 (
            .O(N__23994),
            .I(N__23976));
    LocalMux I__5529 (
            .O(N__23991),
            .I(N__23973));
    LocalMux I__5528 (
            .O(N__23988),
            .I(N__23963));
    InMux I__5527 (
            .O(N__23987),
            .I(N__23960));
    LocalMux I__5526 (
            .O(N__23982),
            .I(N__23951));
    Span4Mux_s2_v I__5525 (
            .O(N__23979),
            .I(N__23944));
    LocalMux I__5524 (
            .O(N__23976),
            .I(N__23944));
    Span4Mux_s3_h I__5523 (
            .O(N__23973),
            .I(N__23944));
    InMux I__5522 (
            .O(N__23972),
            .I(N__23941));
    InMux I__5521 (
            .O(N__23971),
            .I(N__23936));
    InMux I__5520 (
            .O(N__23970),
            .I(N__23936));
    InMux I__5519 (
            .O(N__23969),
            .I(N__23927));
    InMux I__5518 (
            .O(N__23968),
            .I(N__23927));
    InMux I__5517 (
            .O(N__23967),
            .I(N__23927));
    InMux I__5516 (
            .O(N__23966),
            .I(N__23927));
    Span12Mux_s4_h I__5515 (
            .O(N__23963),
            .I(N__23922));
    LocalMux I__5514 (
            .O(N__23960),
            .I(N__23922));
    InMux I__5513 (
            .O(N__23959),
            .I(N__23917));
    InMux I__5512 (
            .O(N__23958),
            .I(N__23917));
    InMux I__5511 (
            .O(N__23957),
            .I(N__23908));
    InMux I__5510 (
            .O(N__23956),
            .I(N__23908));
    InMux I__5509 (
            .O(N__23955),
            .I(N__23908));
    InMux I__5508 (
            .O(N__23954),
            .I(N__23908));
    Odrv4 I__5507 (
            .O(N__23951),
            .I(currentchar_1_2));
    Odrv4 I__5506 (
            .O(N__23944),
            .I(currentchar_1_2));
    LocalMux I__5505 (
            .O(N__23941),
            .I(currentchar_1_2));
    LocalMux I__5504 (
            .O(N__23936),
            .I(currentchar_1_2));
    LocalMux I__5503 (
            .O(N__23927),
            .I(currentchar_1_2));
    Odrv12 I__5502 (
            .O(N__23922),
            .I(currentchar_1_2));
    LocalMux I__5501 (
            .O(N__23917),
            .I(currentchar_1_2));
    LocalMux I__5500 (
            .O(N__23908),
            .I(currentchar_1_2));
    CascadeMux I__5499 (
            .O(N__23891),
            .I(N__23888));
    InMux I__5498 (
            .O(N__23888),
            .I(N__23874));
    InMux I__5497 (
            .O(N__23887),
            .I(N__23871));
    InMux I__5496 (
            .O(N__23886),
            .I(N__23867));
    CascadeMux I__5495 (
            .O(N__23885),
            .I(N__23861));
    CascadeMux I__5494 (
            .O(N__23884),
            .I(N__23856));
    CascadeMux I__5493 (
            .O(N__23883),
            .I(N__23853));
    CascadeMux I__5492 (
            .O(N__23882),
            .I(N__23849));
    CascadeMux I__5491 (
            .O(N__23881),
            .I(N__23846));
    InMux I__5490 (
            .O(N__23880),
            .I(N__23839));
    InMux I__5489 (
            .O(N__23879),
            .I(N__23839));
    InMux I__5488 (
            .O(N__23878),
            .I(N__23836));
    InMux I__5487 (
            .O(N__23877),
            .I(N__23833));
    LocalMux I__5486 (
            .O(N__23874),
            .I(N__23830));
    LocalMux I__5485 (
            .O(N__23871),
            .I(N__23827));
    InMux I__5484 (
            .O(N__23870),
            .I(N__23824));
    LocalMux I__5483 (
            .O(N__23867),
            .I(N__23821));
    CascadeMux I__5482 (
            .O(N__23866),
            .I(N__23818));
    CascadeMux I__5481 (
            .O(N__23865),
            .I(N__23815));
    InMux I__5480 (
            .O(N__23864),
            .I(N__23810));
    InMux I__5479 (
            .O(N__23861),
            .I(N__23810));
    InMux I__5478 (
            .O(N__23860),
            .I(N__23807));
    InMux I__5477 (
            .O(N__23859),
            .I(N__23802));
    InMux I__5476 (
            .O(N__23856),
            .I(N__23802));
    InMux I__5475 (
            .O(N__23853),
            .I(N__23799));
    InMux I__5474 (
            .O(N__23852),
            .I(N__23792));
    InMux I__5473 (
            .O(N__23849),
            .I(N__23792));
    InMux I__5472 (
            .O(N__23846),
            .I(N__23792));
    CascadeMux I__5471 (
            .O(N__23845),
            .I(N__23785));
    InMux I__5470 (
            .O(N__23844),
            .I(N__23782));
    LocalMux I__5469 (
            .O(N__23839),
            .I(N__23779));
    LocalMux I__5468 (
            .O(N__23836),
            .I(N__23774));
    LocalMux I__5467 (
            .O(N__23833),
            .I(N__23774));
    Span4Mux_s1_h I__5466 (
            .O(N__23830),
            .I(N__23765));
    Span4Mux_v I__5465 (
            .O(N__23827),
            .I(N__23765));
    LocalMux I__5464 (
            .O(N__23824),
            .I(N__23765));
    Span4Mux_v I__5463 (
            .O(N__23821),
            .I(N__23765));
    InMux I__5462 (
            .O(N__23818),
            .I(N__23760));
    InMux I__5461 (
            .O(N__23815),
            .I(N__23760));
    LocalMux I__5460 (
            .O(N__23810),
            .I(N__23753));
    LocalMux I__5459 (
            .O(N__23807),
            .I(N__23753));
    LocalMux I__5458 (
            .O(N__23802),
            .I(N__23753));
    LocalMux I__5457 (
            .O(N__23799),
            .I(N__23748));
    LocalMux I__5456 (
            .O(N__23792),
            .I(N__23748));
    InMux I__5455 (
            .O(N__23791),
            .I(N__23745));
    InMux I__5454 (
            .O(N__23790),
            .I(N__23736));
    InMux I__5453 (
            .O(N__23789),
            .I(N__23736));
    InMux I__5452 (
            .O(N__23788),
            .I(N__23736));
    InMux I__5451 (
            .O(N__23785),
            .I(N__23736));
    LocalMux I__5450 (
            .O(N__23782),
            .I(currentchar_m7_0));
    Odrv12 I__5449 (
            .O(N__23779),
            .I(currentchar_m7_0));
    Odrv4 I__5448 (
            .O(N__23774),
            .I(currentchar_m7_0));
    Odrv4 I__5447 (
            .O(N__23765),
            .I(currentchar_m7_0));
    LocalMux I__5446 (
            .O(N__23760),
            .I(currentchar_m7_0));
    Odrv4 I__5445 (
            .O(N__23753),
            .I(currentchar_m7_0));
    Odrv12 I__5444 (
            .O(N__23748),
            .I(currentchar_m7_0));
    LocalMux I__5443 (
            .O(N__23745),
            .I(currentchar_m7_0));
    LocalMux I__5442 (
            .O(N__23736),
            .I(currentchar_m7_0));
    InMux I__5441 (
            .O(N__23717),
            .I(N__23714));
    LocalMux I__5440 (
            .O(N__23714),
            .I(N__23711));
    Span4Mux_v I__5439 (
            .O(N__23711),
            .I(N__23708));
    Span4Mux_h I__5438 (
            .O(N__23708),
            .I(N__23704));
    InMux I__5437 (
            .O(N__23707),
            .I(N__23701));
    Span4Mux_h I__5436 (
            .O(N__23704),
            .I(N__23698));
    LocalMux I__5435 (
            .O(N__23701),
            .I(ScreenBuffer_0_10Z0Z_0));
    Odrv4 I__5434 (
            .O(N__23698),
            .I(ScreenBuffer_0_10Z0Z_0));
    InMux I__5433 (
            .O(N__23693),
            .I(N__23690));
    LocalMux I__5432 (
            .O(N__23690),
            .I(N__23687));
    Span4Mux_s1_h I__5431 (
            .O(N__23687),
            .I(N__23683));
    InMux I__5430 (
            .O(N__23686),
            .I(N__23680));
    Span4Mux_h I__5429 (
            .O(N__23683),
            .I(N__23677));
    LocalMux I__5428 (
            .O(N__23680),
            .I(ScreenBuffer_0_11Z0Z_0));
    Odrv4 I__5427 (
            .O(N__23677),
            .I(ScreenBuffer_0_11Z0Z_0));
    InMux I__5426 (
            .O(N__23672),
            .I(N__23669));
    LocalMux I__5425 (
            .O(N__23669),
            .I(N__23666));
    Span4Mux_v I__5424 (
            .O(N__23666),
            .I(N__23663));
    Odrv4 I__5423 (
            .O(N__23663),
            .I(ScreenBuffer_1_3Z0Z_0));
    CascadeMux I__5422 (
            .O(N__23660),
            .I(currentchar_1_5_ns_1_0_cascade_));
    InMux I__5421 (
            .O(N__23657),
            .I(N__23654));
    LocalMux I__5420 (
            .O(N__23654),
            .I(N__23651));
    Span4Mux_v I__5419 (
            .O(N__23651),
            .I(N__23648));
    Span4Mux_h I__5418 (
            .O(N__23648),
            .I(N__23644));
    InMux I__5417 (
            .O(N__23647),
            .I(N__23641));
    Span4Mux_h I__5416 (
            .O(N__23644),
            .I(N__23638));
    LocalMux I__5415 (
            .O(N__23641),
            .I(ScreenBuffer_0_3Z0Z_0));
    Odrv4 I__5414 (
            .O(N__23638),
            .I(ScreenBuffer_0_3Z0Z_0));
    InMux I__5413 (
            .O(N__23633),
            .I(N__23630));
    LocalMux I__5412 (
            .O(N__23630),
            .I(N__23627));
    Span4Mux_s2_h I__5411 (
            .O(N__23627),
            .I(N__23624));
    Odrv4 I__5410 (
            .O(N__23624),
            .I(beamY_RNIVDIFFI1Z0Z_0));
    InMux I__5409 (
            .O(N__23621),
            .I(N__23618));
    LocalMux I__5408 (
            .O(N__23618),
            .I(beamY_RNI2RNL4M2Z0Z_0));
    InMux I__5407 (
            .O(N__23615),
            .I(N__23609));
    InMux I__5406 (
            .O(N__23614),
            .I(N__23600));
    InMux I__5405 (
            .O(N__23613),
            .I(N__23595));
    InMux I__5404 (
            .O(N__23612),
            .I(N__23595));
    LocalMux I__5403 (
            .O(N__23609),
            .I(N__23592));
    CascadeMux I__5402 (
            .O(N__23608),
            .I(N__23589));
    CascadeMux I__5401 (
            .O(N__23607),
            .I(N__23586));
    CascadeMux I__5400 (
            .O(N__23606),
            .I(N__23582));
    CascadeMux I__5399 (
            .O(N__23605),
            .I(N__23579));
    CascadeMux I__5398 (
            .O(N__23604),
            .I(N__23576));
    CascadeMux I__5397 (
            .O(N__23603),
            .I(N__23573));
    LocalMux I__5396 (
            .O(N__23600),
            .I(N__23568));
    LocalMux I__5395 (
            .O(N__23595),
            .I(N__23568));
    Span4Mux_h I__5394 (
            .O(N__23592),
            .I(N__23565));
    InMux I__5393 (
            .O(N__23589),
            .I(N__23560));
    InMux I__5392 (
            .O(N__23586),
            .I(N__23560));
    InMux I__5391 (
            .O(N__23585),
            .I(N__23555));
    InMux I__5390 (
            .O(N__23582),
            .I(N__23555));
    InMux I__5389 (
            .O(N__23579),
            .I(N__23548));
    InMux I__5388 (
            .O(N__23576),
            .I(N__23548));
    InMux I__5387 (
            .O(N__23573),
            .I(N__23548));
    Span4Mux_v I__5386 (
            .O(N__23568),
            .I(N__23545));
    Odrv4 I__5385 (
            .O(N__23565),
            .I(un3_rowlto1));
    LocalMux I__5384 (
            .O(N__23560),
            .I(un3_rowlto1));
    LocalMux I__5383 (
            .O(N__23555),
            .I(un3_rowlto1));
    LocalMux I__5382 (
            .O(N__23548),
            .I(un3_rowlto1));
    Odrv4 I__5381 (
            .O(N__23545),
            .I(un3_rowlto1));
    CascadeMux I__5380 (
            .O(N__23534),
            .I(N__23531));
    InMux I__5379 (
            .O(N__23531),
            .I(N__23524));
    InMux I__5378 (
            .O(N__23530),
            .I(N__23519));
    InMux I__5377 (
            .O(N__23529),
            .I(N__23519));
    InMux I__5376 (
            .O(N__23528),
            .I(N__23514));
    InMux I__5375 (
            .O(N__23527),
            .I(N__23514));
    LocalMux I__5374 (
            .O(N__23524),
            .I(N__23505));
    LocalMux I__5373 (
            .O(N__23519),
            .I(N__23505));
    LocalMux I__5372 (
            .O(N__23514),
            .I(N__23499));
    InMux I__5371 (
            .O(N__23513),
            .I(N__23496));
    InMux I__5370 (
            .O(N__23512),
            .I(N__23489));
    InMux I__5369 (
            .O(N__23511),
            .I(N__23489));
    InMux I__5368 (
            .O(N__23510),
            .I(N__23489));
    Span4Mux_v I__5367 (
            .O(N__23505),
            .I(N__23486));
    InMux I__5366 (
            .O(N__23504),
            .I(N__23479));
    InMux I__5365 (
            .O(N__23503),
            .I(N__23479));
    InMux I__5364 (
            .O(N__23502),
            .I(N__23479));
    Span4Mux_v I__5363 (
            .O(N__23499),
            .I(N__23468));
    LocalMux I__5362 (
            .O(N__23496),
            .I(N__23468));
    LocalMux I__5361 (
            .O(N__23489),
            .I(N__23468));
    Span4Mux_h I__5360 (
            .O(N__23486),
            .I(N__23468));
    LocalMux I__5359 (
            .O(N__23479),
            .I(N__23468));
    Odrv4 I__5358 (
            .O(N__23468),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1));
    CascadeMux I__5357 (
            .O(N__23465),
            .I(N__23461));
    CascadeMux I__5356 (
            .O(N__23464),
            .I(N__23458));
    InMux I__5355 (
            .O(N__23461),
            .I(N__23453));
    InMux I__5354 (
            .O(N__23458),
            .I(N__23453));
    LocalMux I__5353 (
            .O(N__23453),
            .I(N__23450));
    Odrv4 I__5352 (
            .O(N__23450),
            .I(N_52));
    CascadeMux I__5351 (
            .O(N__23447),
            .I(N__23444));
    InMux I__5350 (
            .O(N__23444),
            .I(N__23440));
    InMux I__5349 (
            .O(N__23443),
            .I(N__23436));
    LocalMux I__5348 (
            .O(N__23440),
            .I(N__23430));
    CascadeMux I__5347 (
            .O(N__23439),
            .I(N__23426));
    LocalMux I__5346 (
            .O(N__23436),
            .I(N__23418));
    InMux I__5345 (
            .O(N__23435),
            .I(N__23413));
    InMux I__5344 (
            .O(N__23434),
            .I(N__23413));
    InMux I__5343 (
            .O(N__23433),
            .I(N__23410));
    Span4Mux_s3_h I__5342 (
            .O(N__23430),
            .I(N__23407));
    InMux I__5341 (
            .O(N__23429),
            .I(N__23404));
    InMux I__5340 (
            .O(N__23426),
            .I(N__23399));
    InMux I__5339 (
            .O(N__23425),
            .I(N__23399));
    InMux I__5338 (
            .O(N__23424),
            .I(N__23390));
    InMux I__5337 (
            .O(N__23423),
            .I(N__23390));
    InMux I__5336 (
            .O(N__23422),
            .I(N__23390));
    InMux I__5335 (
            .O(N__23421),
            .I(N__23390));
    Odrv4 I__5334 (
            .O(N__23418),
            .I(un112_pixel_2_8));
    LocalMux I__5333 (
            .O(N__23413),
            .I(un112_pixel_2_8));
    LocalMux I__5332 (
            .O(N__23410),
            .I(un112_pixel_2_8));
    Odrv4 I__5331 (
            .O(N__23407),
            .I(un112_pixel_2_8));
    LocalMux I__5330 (
            .O(N__23404),
            .I(un112_pixel_2_8));
    LocalMux I__5329 (
            .O(N__23399),
            .I(un112_pixel_2_8));
    LocalMux I__5328 (
            .O(N__23390),
            .I(un112_pixel_2_8));
    CascadeMux I__5327 (
            .O(N__23375),
            .I(N_4581_0_cascade_));
    CascadeMux I__5326 (
            .O(N__23372),
            .I(N_1296_0_cascade_));
    InMux I__5325 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__5324 (
            .O(N__23366),
            .I(N_1296_0));
    CascadeMux I__5323 (
            .O(N__23363),
            .I(N__23360));
    InMux I__5322 (
            .O(N__23360),
            .I(N__23354));
    InMux I__5321 (
            .O(N__23359),
            .I(N__23354));
    LocalMux I__5320 (
            .O(N__23354),
            .I(N__23350));
    InMux I__5319 (
            .O(N__23353),
            .I(N__23340));
    Span4Mux_v I__5318 (
            .O(N__23350),
            .I(N__23337));
    CascadeMux I__5317 (
            .O(N__23349),
            .I(N__23332));
    InMux I__5316 (
            .O(N__23348),
            .I(N__23329));
    InMux I__5315 (
            .O(N__23347),
            .I(N__23326));
    InMux I__5314 (
            .O(N__23346),
            .I(N__23323));
    CascadeMux I__5313 (
            .O(N__23345),
            .I(N__23319));
    InMux I__5312 (
            .O(N__23344),
            .I(N__23314));
    InMux I__5311 (
            .O(N__23343),
            .I(N__23314));
    LocalMux I__5310 (
            .O(N__23340),
            .I(N__23311));
    IoSpan4Mux I__5309 (
            .O(N__23337),
            .I(N__23308));
    InMux I__5308 (
            .O(N__23336),
            .I(N__23303));
    InMux I__5307 (
            .O(N__23335),
            .I(N__23303));
    InMux I__5306 (
            .O(N__23332),
            .I(N__23297));
    LocalMux I__5305 (
            .O(N__23329),
            .I(N__23294));
    LocalMux I__5304 (
            .O(N__23326),
            .I(N__23289));
    LocalMux I__5303 (
            .O(N__23323),
            .I(N__23289));
    InMux I__5302 (
            .O(N__23322),
            .I(N__23286));
    InMux I__5301 (
            .O(N__23319),
            .I(N__23281));
    LocalMux I__5300 (
            .O(N__23314),
            .I(N__23272));
    Span4Mux_v I__5299 (
            .O(N__23311),
            .I(N__23272));
    Span4Mux_s2_h I__5298 (
            .O(N__23308),
            .I(N__23272));
    LocalMux I__5297 (
            .O(N__23303),
            .I(N__23272));
    InMux I__5296 (
            .O(N__23302),
            .I(N__23269));
    InMux I__5295 (
            .O(N__23301),
            .I(N__23266));
    InMux I__5294 (
            .O(N__23300),
            .I(N__23261));
    LocalMux I__5293 (
            .O(N__23297),
            .I(N__23254));
    Span4Mux_h I__5292 (
            .O(N__23294),
            .I(N__23254));
    Span4Mux_s3_v I__5291 (
            .O(N__23289),
            .I(N__23254));
    LocalMux I__5290 (
            .O(N__23286),
            .I(N__23251));
    InMux I__5289 (
            .O(N__23285),
            .I(N__23248));
    InMux I__5288 (
            .O(N__23284),
            .I(N__23245));
    LocalMux I__5287 (
            .O(N__23281),
            .I(N__23236));
    Span4Mux_v I__5286 (
            .O(N__23272),
            .I(N__23236));
    LocalMux I__5285 (
            .O(N__23269),
            .I(N__23236));
    LocalMux I__5284 (
            .O(N__23266),
            .I(N__23233));
    InMux I__5283 (
            .O(N__23265),
            .I(N__23226));
    InMux I__5282 (
            .O(N__23264),
            .I(N__23226));
    LocalMux I__5281 (
            .O(N__23261),
            .I(N__23217));
    Span4Mux_v I__5280 (
            .O(N__23254),
            .I(N__23217));
    Span4Mux_v I__5279 (
            .O(N__23251),
            .I(N__23217));
    LocalMux I__5278 (
            .O(N__23248),
            .I(N__23217));
    LocalMux I__5277 (
            .O(N__23245),
            .I(N__23214));
    InMux I__5276 (
            .O(N__23244),
            .I(N__23209));
    InMux I__5275 (
            .O(N__23243),
            .I(N__23209));
    Span4Mux_h I__5274 (
            .O(N__23236),
            .I(N__23206));
    Span4Mux_h I__5273 (
            .O(N__23233),
            .I(N__23203));
    InMux I__5272 (
            .O(N__23232),
            .I(N__23200));
    InMux I__5271 (
            .O(N__23231),
            .I(N__23197));
    LocalMux I__5270 (
            .O(N__23226),
            .I(N__23192));
    Span4Mux_v I__5269 (
            .O(N__23217),
            .I(N__23192));
    Span4Mux_h I__5268 (
            .O(N__23214),
            .I(N__23185));
    LocalMux I__5267 (
            .O(N__23209),
            .I(N__23185));
    Span4Mux_v I__5266 (
            .O(N__23206),
            .I(N__23185));
    Odrv4 I__5265 (
            .O(N__23203),
            .I(beamYZ0Z_1));
    LocalMux I__5264 (
            .O(N__23200),
            .I(beamYZ0Z_1));
    LocalMux I__5263 (
            .O(N__23197),
            .I(beamYZ0Z_1));
    Odrv4 I__5262 (
            .O(N__23192),
            .I(beamYZ0Z_1));
    Odrv4 I__5261 (
            .O(N__23185),
            .I(beamYZ0Z_1));
    CascadeMux I__5260 (
            .O(N__23174),
            .I(N__23171));
    InMux I__5259 (
            .O(N__23171),
            .I(N__23168));
    LocalMux I__5258 (
            .O(N__23168),
            .I(N__23165));
    Span4Mux_v I__5257 (
            .O(N__23165),
            .I(N__23162));
    Odrv4 I__5256 (
            .O(N__23162),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    InMux I__5255 (
            .O(N__23159),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__5254 (
            .O(N__23156),
            .I(N__23153));
    LocalMux I__5253 (
            .O(N__23153),
            .I(if_generate_plus_mult1_un75_sum_axb_4_l_fx));
    CascadeMux I__5252 (
            .O(N__23150),
            .I(N__23147));
    InMux I__5251 (
            .O(N__23147),
            .I(N__23143));
    InMux I__5250 (
            .O(N__23146),
            .I(N__23140));
    LocalMux I__5249 (
            .O(N__23143),
            .I(N__23137));
    LocalMux I__5248 (
            .O(N__23140),
            .I(N__23134));
    Span4Mux_s3_h I__5247 (
            .O(N__23137),
            .I(N__23131));
    Odrv4 I__5246 (
            .O(N__23134),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    Odrv4 I__5245 (
            .O(N__23131),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    InMux I__5244 (
            .O(N__23126),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__5243 (
            .O(N__23123),
            .I(N__23120));
    LocalMux I__5242 (
            .O(N__23120),
            .I(N__23117));
    Span4Mux_s3_h I__5241 (
            .O(N__23117),
            .I(N__23114));
    Odrv4 I__5240 (
            .O(N__23114),
            .I(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__5239 (
            .O(N__23111),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__5238 (
            .O(N__23108),
            .I(N__23105));
    LocalMux I__5237 (
            .O(N__23105),
            .I(N__23102));
    Span4Mux_h I__5236 (
            .O(N__23102),
            .I(N__23099));
    Span4Mux_h I__5235 (
            .O(N__23099),
            .I(N__23096));
    Odrv4 I__5234 (
            .O(N__23096),
            .I(un6_rowlt7_0));
    InMux I__5233 (
            .O(N__23093),
            .I(N__23090));
    LocalMux I__5232 (
            .O(N__23090),
            .I(N__23085));
    InMux I__5231 (
            .O(N__23089),
            .I(N__23082));
    InMux I__5230 (
            .O(N__23088),
            .I(N__23077));
    Span4Mux_v I__5229 (
            .O(N__23085),
            .I(N__23074));
    LocalMux I__5228 (
            .O(N__23082),
            .I(N__23071));
    InMux I__5227 (
            .O(N__23081),
            .I(N__23068));
    InMux I__5226 (
            .O(N__23080),
            .I(N__23065));
    LocalMux I__5225 (
            .O(N__23077),
            .I(N__23062));
    Span4Mux_h I__5224 (
            .O(N__23074),
            .I(N__23059));
    Span4Mux_v I__5223 (
            .O(N__23071),
            .I(N__23054));
    LocalMux I__5222 (
            .O(N__23068),
            .I(N__23054));
    LocalMux I__5221 (
            .O(N__23065),
            .I(N__23051));
    Odrv12 I__5220 (
            .O(N__23062),
            .I(chessboardpixel_un151_pixel_24));
    Odrv4 I__5219 (
            .O(N__23059),
            .I(chessboardpixel_un151_pixel_24));
    Odrv4 I__5218 (
            .O(N__23054),
            .I(chessboardpixel_un151_pixel_24));
    Odrv12 I__5217 (
            .O(N__23051),
            .I(chessboardpixel_un151_pixel_24));
    CascadeMux I__5216 (
            .O(N__23042),
            .I(N__23039));
    InMux I__5215 (
            .O(N__23039),
            .I(N__23036));
    LocalMux I__5214 (
            .O(N__23036),
            .I(column_1_if_generate_plus_mult1_un68_sum_iZ0));
    CascadeMux I__5213 (
            .O(N__23033),
            .I(N__23027));
    InMux I__5212 (
            .O(N__23032),
            .I(N__23024));
    CascadeMux I__5211 (
            .O(N__23031),
            .I(N__23021));
    CascadeMux I__5210 (
            .O(N__23030),
            .I(N__23012));
    InMux I__5209 (
            .O(N__23027),
            .I(N__23009));
    LocalMux I__5208 (
            .O(N__23024),
            .I(N__23006));
    InMux I__5207 (
            .O(N__23021),
            .I(N__23003));
    InMux I__5206 (
            .O(N__23020),
            .I(N__22998));
    InMux I__5205 (
            .O(N__23019),
            .I(N__22998));
    CascadeMux I__5204 (
            .O(N__23018),
            .I(N__22995));
    InMux I__5203 (
            .O(N__23017),
            .I(N__22991));
    CascadeMux I__5202 (
            .O(N__23016),
            .I(N__22987));
    InMux I__5201 (
            .O(N__23015),
            .I(N__22979));
    InMux I__5200 (
            .O(N__23012),
            .I(N__22979));
    LocalMux I__5199 (
            .O(N__23009),
            .I(N__22970));
    Span4Mux_v I__5198 (
            .O(N__23006),
            .I(N__22970));
    LocalMux I__5197 (
            .O(N__23003),
            .I(N__22970));
    LocalMux I__5196 (
            .O(N__22998),
            .I(N__22970));
    InMux I__5195 (
            .O(N__22995),
            .I(N__22965));
    InMux I__5194 (
            .O(N__22994),
            .I(N__22965));
    LocalMux I__5193 (
            .O(N__22991),
            .I(N__22962));
    InMux I__5192 (
            .O(N__22990),
            .I(N__22957));
    InMux I__5191 (
            .O(N__22987),
            .I(N__22957));
    CascadeMux I__5190 (
            .O(N__22986),
            .I(N__22954));
    CascadeMux I__5189 (
            .O(N__22985),
            .I(N__22951));
    InMux I__5188 (
            .O(N__22984),
            .I(N__22948));
    LocalMux I__5187 (
            .O(N__22979),
            .I(N__22945));
    Span4Mux_h I__5186 (
            .O(N__22970),
            .I(N__22940));
    LocalMux I__5185 (
            .O(N__22965),
            .I(N__22940));
    Span4Mux_v I__5184 (
            .O(N__22962),
            .I(N__22935));
    LocalMux I__5183 (
            .O(N__22957),
            .I(N__22935));
    InMux I__5182 (
            .O(N__22954),
            .I(N__22930));
    InMux I__5181 (
            .O(N__22951),
            .I(N__22930));
    LocalMux I__5180 (
            .O(N__22948),
            .I(un3_rowlto0));
    Odrv12 I__5179 (
            .O(N__22945),
            .I(un3_rowlto0));
    Odrv4 I__5178 (
            .O(N__22940),
            .I(un3_rowlto0));
    Odrv4 I__5177 (
            .O(N__22935),
            .I(un3_rowlto0));
    LocalMux I__5176 (
            .O(N__22930),
            .I(un3_rowlto0));
    InMux I__5175 (
            .O(N__22919),
            .I(N__22916));
    LocalMux I__5174 (
            .O(N__22916),
            .I(N__22913));
    Span4Mux_h I__5173 (
            .O(N__22913),
            .I(N__22910));
    Odrv4 I__5172 (
            .O(N__22910),
            .I(un113_pixel_3_0_11__currentchar_m7_0Z0Z_1));
    CascadeMux I__5171 (
            .O(N__22907),
            .I(d_N_3_mux_cascade_));
    InMux I__5170 (
            .O(N__22904),
            .I(N__22901));
    LocalMux I__5169 (
            .O(N__22901),
            .I(N__22898));
    Span4Mux_v I__5168 (
            .O(N__22898),
            .I(N__22895));
    Span4Mux_h I__5167 (
            .O(N__22895),
            .I(N__22892));
    Odrv4 I__5166 (
            .O(N__22892),
            .I(ScreenBuffer_1_2Z0Z_2));
    InMux I__5165 (
            .O(N__22889),
            .I(N__22886));
    LocalMux I__5164 (
            .O(N__22886),
            .I(N__22883));
    Span4Mux_s2_h I__5163 (
            .O(N__22883),
            .I(N__22880));
    Span4Mux_h I__5162 (
            .O(N__22880),
            .I(N__22877));
    Odrv4 I__5161 (
            .O(N__22877),
            .I(ScreenBuffer_1_1Z0Z_2));
    InMux I__5160 (
            .O(N__22874),
            .I(N__22871));
    LocalMux I__5159 (
            .O(N__22871),
            .I(N__22868));
    Span4Mux_h I__5158 (
            .O(N__22868),
            .I(N__22865));
    Odrv4 I__5157 (
            .O(N__22865),
            .I(un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2));
    CascadeMux I__5156 (
            .O(N__22862),
            .I(N__22859));
    InMux I__5155 (
            .O(N__22859),
            .I(N__22856));
    LocalMux I__5154 (
            .O(N__22856),
            .I(N__22853));
    Odrv12 I__5153 (
            .O(N__22853),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0));
    CascadeMux I__5152 (
            .O(N__22850),
            .I(N__22847));
    InMux I__5151 (
            .O(N__22847),
            .I(N__22844));
    LocalMux I__5150 (
            .O(N__22844),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2));
    InMux I__5149 (
            .O(N__22841),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__5148 (
            .O(N__22838),
            .I(N__22835));
    LocalMux I__5147 (
            .O(N__22835),
            .I(charx_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__5146 (
            .O(N__22832),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__5145 (
            .O(N__22829),
            .I(N__22826));
    LocalMux I__5144 (
            .O(N__22826),
            .I(N__22823));
    Odrv12 I__5143 (
            .O(N__22823),
            .I(charx_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__5142 (
            .O(N__22820),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__5141 (
            .O(N__22817),
            .I(N__22814));
    LocalMux I__5140 (
            .O(N__22814),
            .I(N__22809));
    InMux I__5139 (
            .O(N__22813),
            .I(N__22806));
    InMux I__5138 (
            .O(N__22812),
            .I(N__22803));
    Span4Mux_h I__5137 (
            .O(N__22809),
            .I(N__22800));
    LocalMux I__5136 (
            .O(N__22806),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    LocalMux I__5135 (
            .O(N__22803),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    Odrv4 I__5134 (
            .O(N__22800),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    CascadeMux I__5133 (
            .O(N__22793),
            .I(N__22789));
    InMux I__5132 (
            .O(N__22792),
            .I(N__22784));
    InMux I__5131 (
            .O(N__22789),
            .I(N__22784));
    LocalMux I__5130 (
            .O(N__22784),
            .I(N__22781));
    Odrv12 I__5129 (
            .O(N__22781),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1));
    InMux I__5128 (
            .O(N__22778),
            .I(N__22773));
    InMux I__5127 (
            .O(N__22777),
            .I(N__22770));
    InMux I__5126 (
            .O(N__22776),
            .I(N__22766));
    LocalMux I__5125 (
            .O(N__22773),
            .I(N__22761));
    LocalMux I__5124 (
            .O(N__22770),
            .I(N__22761));
    InMux I__5123 (
            .O(N__22769),
            .I(N__22758));
    LocalMux I__5122 (
            .O(N__22766),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    Odrv12 I__5121 (
            .O(N__22761),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    LocalMux I__5120 (
            .O(N__22758),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    InMux I__5119 (
            .O(N__22751),
            .I(N__22748));
    LocalMux I__5118 (
            .O(N__22748),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73));
    CascadeMux I__5117 (
            .O(N__22745),
            .I(N__22740));
    InMux I__5116 (
            .O(N__22744),
            .I(N__22737));
    InMux I__5115 (
            .O(N__22743),
            .I(N__22733));
    InMux I__5114 (
            .O(N__22740),
            .I(N__22727));
    LocalMux I__5113 (
            .O(N__22737),
            .I(N__22724));
    InMux I__5112 (
            .O(N__22736),
            .I(N__22721));
    LocalMux I__5111 (
            .O(N__22733),
            .I(N__22717));
    InMux I__5110 (
            .O(N__22732),
            .I(N__22712));
    InMux I__5109 (
            .O(N__22731),
            .I(N__22712));
    InMux I__5108 (
            .O(N__22730),
            .I(N__22709));
    LocalMux I__5107 (
            .O(N__22727),
            .I(N__22704));
    Span4Mux_v I__5106 (
            .O(N__22724),
            .I(N__22704));
    LocalMux I__5105 (
            .O(N__22721),
            .I(N__22701));
    InMux I__5104 (
            .O(N__22720),
            .I(N__22698));
    Span4Mux_v I__5103 (
            .O(N__22717),
            .I(N__22695));
    LocalMux I__5102 (
            .O(N__22712),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__5101 (
            .O(N__22709),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__5100 (
            .O(N__22704),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv12 I__5099 (
            .O(N__22701),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__5098 (
            .O(N__22698),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__5097 (
            .O(N__22695),
            .I(charx_if_generate_plus_mult1_un40_sum));
    CascadeMux I__5096 (
            .O(N__22682),
            .I(N__22679));
    InMux I__5095 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__5094 (
            .O(N__22676),
            .I(charx_if_generate_plus_mult1_un40_sum_i));
    InMux I__5093 (
            .O(N__22673),
            .I(N__22669));
    InMux I__5092 (
            .O(N__22672),
            .I(N__22666));
    LocalMux I__5091 (
            .O(N__22669),
            .I(N__22659));
    LocalMux I__5090 (
            .O(N__22666),
            .I(N__22659));
    InMux I__5089 (
            .O(N__22665),
            .I(N__22656));
    InMux I__5088 (
            .O(N__22664),
            .I(N__22653));
    Span4Mux_v I__5087 (
            .O(N__22659),
            .I(N__22650));
    LocalMux I__5086 (
            .O(N__22656),
            .I(N__22645));
    LocalMux I__5085 (
            .O(N__22653),
            .I(N__22645));
    Span4Mux_h I__5084 (
            .O(N__22650),
            .I(N__22642));
    Span4Mux_v I__5083 (
            .O(N__22645),
            .I(N__22639));
    Odrv4 I__5082 (
            .O(N__22642),
            .I(charx_if_generate_plus_mult1_un68_sum));
    Odrv4 I__5081 (
            .O(N__22639),
            .I(charx_if_generate_plus_mult1_un68_sum));
    InMux I__5080 (
            .O(N__22634),
            .I(N__22631));
    LocalMux I__5079 (
            .O(N__22631),
            .I(N__22628));
    Odrv12 I__5078 (
            .O(N__22628),
            .I(column_1_i_i_2));
    InMux I__5077 (
            .O(N__22625),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_1));
    CascadeMux I__5076 (
            .O(N__22622),
            .I(N__22615));
    CascadeMux I__5075 (
            .O(N__22621),
            .I(N__22612));
    InMux I__5074 (
            .O(N__22620),
            .I(N__22608));
    InMux I__5073 (
            .O(N__22619),
            .I(N__22604));
    InMux I__5072 (
            .O(N__22618),
            .I(N__22601));
    InMux I__5071 (
            .O(N__22615),
            .I(N__22598));
    InMux I__5070 (
            .O(N__22612),
            .I(N__22593));
    InMux I__5069 (
            .O(N__22611),
            .I(N__22593));
    LocalMux I__5068 (
            .O(N__22608),
            .I(N__22590));
    InMux I__5067 (
            .O(N__22607),
            .I(N__22587));
    LocalMux I__5066 (
            .O(N__22604),
            .I(N__22582));
    LocalMux I__5065 (
            .O(N__22601),
            .I(N__22582));
    LocalMux I__5064 (
            .O(N__22598),
            .I(N__22577));
    LocalMux I__5063 (
            .O(N__22593),
            .I(N__22577));
    Span4Mux_s3_h I__5062 (
            .O(N__22590),
            .I(N__22574));
    LocalMux I__5061 (
            .O(N__22587),
            .I(N__22569));
    Span4Mux_v I__5060 (
            .O(N__22582),
            .I(N__22569));
    Odrv4 I__5059 (
            .O(N__22577),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__5058 (
            .O(N__22574),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__5057 (
            .O(N__22569),
            .I(charx_if_generate_plus_mult1_un54_sum));
    CascadeMux I__5056 (
            .O(N__22562),
            .I(N__22559));
    InMux I__5055 (
            .O(N__22559),
            .I(N__22556));
    LocalMux I__5054 (
            .O(N__22556),
            .I(N__22553));
    Span4Mux_h I__5053 (
            .O(N__22553),
            .I(N__22550));
    Odrv4 I__5052 (
            .O(N__22550),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3));
    InMux I__5051 (
            .O(N__22547),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1));
    CascadeMux I__5050 (
            .O(N__22544),
            .I(N__22541));
    InMux I__5049 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__5048 (
            .O(N__22538),
            .I(N__22535));
    Span4Mux_h I__5047 (
            .O(N__22535),
            .I(N__22532));
    Odrv4 I__5046 (
            .O(N__22532),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5));
    InMux I__5045 (
            .O(N__22529),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__5044 (
            .O(N__22526),
            .I(N__22520));
    InMux I__5043 (
            .O(N__22525),
            .I(N__22520));
    LocalMux I__5042 (
            .O(N__22520),
            .I(N__22517));
    Odrv4 I__5041 (
            .O(N__22517),
            .I(charx_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__5040 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__5039 (
            .O(N__22511),
            .I(N__22508));
    Span4Mux_h I__5038 (
            .O(N__22508),
            .I(N__22505));
    Odrv4 I__5037 (
            .O(N__22505),
            .I(charx_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__5036 (
            .O(N__22502),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__5035 (
            .O(N__22499),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__5034 (
            .O(N__22496),
            .I(N__22493));
    LocalMux I__5033 (
            .O(N__22493),
            .I(N__22488));
    InMux I__5032 (
            .O(N__22492),
            .I(N__22485));
    InMux I__5031 (
            .O(N__22491),
            .I(N__22482));
    Span4Mux_v I__5030 (
            .O(N__22488),
            .I(N__22477));
    LocalMux I__5029 (
            .O(N__22485),
            .I(N__22477));
    LocalMux I__5028 (
            .O(N__22482),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8));
    Odrv4 I__5027 (
            .O(N__22477),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8));
    CascadeMux I__5026 (
            .O(N__22472),
            .I(N__22469));
    InMux I__5025 (
            .O(N__22469),
            .I(N__22466));
    LocalMux I__5024 (
            .O(N__22466),
            .I(charx_if_generate_plus_mult1_un47_sum_i));
    InMux I__5023 (
            .O(N__22463),
            .I(N__22456));
    InMux I__5022 (
            .O(N__22462),
            .I(N__22453));
    InMux I__5021 (
            .O(N__22461),
            .I(N__22450));
    InMux I__5020 (
            .O(N__22460),
            .I(N__22446));
    InMux I__5019 (
            .O(N__22459),
            .I(N__22443));
    LocalMux I__5018 (
            .O(N__22456),
            .I(N__22440));
    LocalMux I__5017 (
            .O(N__22453),
            .I(N__22437));
    LocalMux I__5016 (
            .O(N__22450),
            .I(N__22434));
    InMux I__5015 (
            .O(N__22449),
            .I(N__22431));
    LocalMux I__5014 (
            .O(N__22446),
            .I(N__22428));
    LocalMux I__5013 (
            .O(N__22443),
            .I(N__22425));
    Span4Mux_h I__5012 (
            .O(N__22440),
            .I(N__22422));
    Span4Mux_h I__5011 (
            .O(N__22437),
            .I(N__22413));
    Span4Mux_v I__5010 (
            .O(N__22434),
            .I(N__22413));
    LocalMux I__5009 (
            .O(N__22431),
            .I(N__22413));
    Span4Mux_s3_h I__5008 (
            .O(N__22428),
            .I(N__22413));
    Odrv4 I__5007 (
            .O(N__22425),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__5006 (
            .O(N__22422),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__5005 (
            .O(N__22413),
            .I(charx_if_generate_plus_mult1_un47_sum));
    InMux I__5004 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__5003 (
            .O(N__22403),
            .I(N__22400));
    Odrv4 I__5002 (
            .O(N__22400),
            .I(charx_if_generate_plus_mult1_un40_sum_i_5));
    CascadeMux I__5001 (
            .O(N__22397),
            .I(N__22394));
    InMux I__5000 (
            .O(N__22394),
            .I(N__22391));
    LocalMux I__4999 (
            .O(N__22391),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1));
    InMux I__4998 (
            .O(N__22388),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1));
    InMux I__4997 (
            .O(N__22385),
            .I(N__22382));
    LocalMux I__4996 (
            .O(N__22382),
            .I(N__22379));
    Odrv12 I__4995 (
            .O(N__22379),
            .I(column_1_if_generate_plus_mult1_un47_sum1_2));
    InMux I__4994 (
            .O(N__22376),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_1));
    InMux I__4993 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__4992 (
            .O(N__22370),
            .I(N__22367));
    Span4Mux_h I__4991 (
            .O(N__22367),
            .I(N__22364));
    Odrv4 I__4990 (
            .O(N__22364),
            .I(column_1_if_generate_plus_mult1_un47_sum1_3));
    InMux I__4989 (
            .O(N__22361),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_2));
    InMux I__4988 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__4987 (
            .O(N__22355),
            .I(N__22352));
    Odrv4 I__4986 (
            .O(N__22352),
            .I(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx));
    CascadeMux I__4985 (
            .O(N__22349),
            .I(N__22346));
    InMux I__4984 (
            .O(N__22346),
            .I(N__22343));
    LocalMux I__4983 (
            .O(N__22343),
            .I(N__22340));
    Span4Mux_h I__4982 (
            .O(N__22340),
            .I(N__22337));
    Odrv4 I__4981 (
            .O(N__22337),
            .I(column_1_if_generate_plus_mult1_un47_sum1_4));
    InMux I__4980 (
            .O(N__22334),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_3));
    CascadeMux I__4979 (
            .O(N__22331),
            .I(N__22327));
    InMux I__4978 (
            .O(N__22330),
            .I(N__22324));
    InMux I__4977 (
            .O(N__22327),
            .I(N__22321));
    LocalMux I__4976 (
            .O(N__22324),
            .I(N__22314));
    LocalMux I__4975 (
            .O(N__22321),
            .I(N__22314));
    CascadeMux I__4974 (
            .O(N__22320),
            .I(N__22311));
    InMux I__4973 (
            .O(N__22319),
            .I(N__22306));
    Span4Mux_s3_v I__4972 (
            .O(N__22314),
            .I(N__22302));
    InMux I__4971 (
            .O(N__22311),
            .I(N__22299));
    InMux I__4970 (
            .O(N__22310),
            .I(N__22296));
    InMux I__4969 (
            .O(N__22309),
            .I(N__22293));
    LocalMux I__4968 (
            .O(N__22306),
            .I(N__22290));
    InMux I__4967 (
            .O(N__22305),
            .I(N__22287));
    Odrv4 I__4966 (
            .O(N__22302),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__4965 (
            .O(N__22299),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__4964 (
            .O(N__22296),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__4963 (
            .O(N__22293),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    Odrv4 I__4962 (
            .O(N__22290),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__4961 (
            .O(N__22287),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    InMux I__4960 (
            .O(N__22274),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_4));
    InMux I__4959 (
            .O(N__22271),
            .I(N__22265));
    InMux I__4958 (
            .O(N__22270),
            .I(N__22265));
    LocalMux I__4957 (
            .O(N__22265),
            .I(N__22262));
    Odrv4 I__4956 (
            .O(N__22262),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5));
    InMux I__4955 (
            .O(N__22259),
            .I(N__22246));
    InMux I__4954 (
            .O(N__22258),
            .I(N__22246));
    InMux I__4953 (
            .O(N__22257),
            .I(N__22243));
    InMux I__4952 (
            .O(N__22256),
            .I(N__22238));
    InMux I__4951 (
            .O(N__22255),
            .I(N__22238));
    InMux I__4950 (
            .O(N__22254),
            .I(N__22235));
    InMux I__4949 (
            .O(N__22253),
            .I(N__22232));
    InMux I__4948 (
            .O(N__22252),
            .I(N__22229));
    InMux I__4947 (
            .O(N__22251),
            .I(N__22226));
    LocalMux I__4946 (
            .O(N__22246),
            .I(N__22223));
    LocalMux I__4945 (
            .O(N__22243),
            .I(N__22220));
    LocalMux I__4944 (
            .O(N__22238),
            .I(N__22217));
    LocalMux I__4943 (
            .O(N__22235),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__4942 (
            .O(N__22232),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__4941 (
            .O(N__22229),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__4940 (
            .O(N__22226),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv12 I__4939 (
            .O(N__22223),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv4 I__4938 (
            .O(N__22220),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv4 I__4937 (
            .O(N__22217),
            .I(charx_if_generate_plus_mult1_un33_sum));
    InMux I__4936 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__4935 (
            .O(N__22199),
            .I(N__22196));
    Odrv4 I__4934 (
            .O(N__22196),
            .I(un5_visiblex_i_0_25));
    InMux I__4933 (
            .O(N__22193),
            .I(N__22189));
    InMux I__4932 (
            .O(N__22192),
            .I(N__22185));
    LocalMux I__4931 (
            .O(N__22189),
            .I(N__22182));
    InMux I__4930 (
            .O(N__22188),
            .I(N__22179));
    LocalMux I__4929 (
            .O(N__22185),
            .I(N__22176));
    Span4Mux_s3_h I__4928 (
            .O(N__22182),
            .I(N__22171));
    LocalMux I__4927 (
            .O(N__22179),
            .I(N__22171));
    Span4Mux_s2_h I__4926 (
            .O(N__22176),
            .I(N__22168));
    Odrv4 I__4925 (
            .O(N__22171),
            .I(N_56));
    Odrv4 I__4924 (
            .O(N__22168),
            .I(N_56));
    InMux I__4923 (
            .O(N__22163),
            .I(N__22159));
    InMux I__4922 (
            .O(N__22162),
            .I(N__22154));
    LocalMux I__4921 (
            .O(N__22159),
            .I(N__22151));
    InMux I__4920 (
            .O(N__22158),
            .I(N__22148));
    CascadeMux I__4919 (
            .O(N__22157),
            .I(N__22144));
    LocalMux I__4918 (
            .O(N__22154),
            .I(N__22137));
    Span4Mux_s2_v I__4917 (
            .O(N__22151),
            .I(N__22132));
    LocalMux I__4916 (
            .O(N__22148),
            .I(N__22132));
    InMux I__4915 (
            .O(N__22147),
            .I(N__22127));
    InMux I__4914 (
            .O(N__22144),
            .I(N__22127));
    InMux I__4913 (
            .O(N__22143),
            .I(N__22120));
    InMux I__4912 (
            .O(N__22142),
            .I(N__22120));
    InMux I__4911 (
            .O(N__22141),
            .I(N__22120));
    InMux I__4910 (
            .O(N__22140),
            .I(N__22117));
    Span4Mux_h I__4909 (
            .O(N__22137),
            .I(N__22112));
    Span4Mux_h I__4908 (
            .O(N__22132),
            .I(N__22112));
    LocalMux I__4907 (
            .O(N__22127),
            .I(N__22107));
    LocalMux I__4906 (
            .O(N__22120),
            .I(N__22107));
    LocalMux I__4905 (
            .O(N__22117),
            .I(N_32_i));
    Odrv4 I__4904 (
            .O(N__22112),
            .I(N_32_i));
    Odrv4 I__4903 (
            .O(N__22107),
            .I(N_32_i));
    InMux I__4902 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__4901 (
            .O(N__22097),
            .I(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx));
    CascadeMux I__4900 (
            .O(N__22094),
            .I(N__22089));
    CascadeMux I__4899 (
            .O(N__22093),
            .I(N__22081));
    CascadeMux I__4898 (
            .O(N__22092),
            .I(N__22078));
    InMux I__4897 (
            .O(N__22089),
            .I(N__22068));
    InMux I__4896 (
            .O(N__22088),
            .I(N__22060));
    InMux I__4895 (
            .O(N__22087),
            .I(N__22060));
    InMux I__4894 (
            .O(N__22086),
            .I(N__22060));
    InMux I__4893 (
            .O(N__22085),
            .I(N__22057));
    InMux I__4892 (
            .O(N__22084),
            .I(N__22048));
    InMux I__4891 (
            .O(N__22081),
            .I(N__22048));
    InMux I__4890 (
            .O(N__22078),
            .I(N__22048));
    InMux I__4889 (
            .O(N__22077),
            .I(N__22048));
    InMux I__4888 (
            .O(N__22076),
            .I(N__22045));
    InMux I__4887 (
            .O(N__22075),
            .I(N__22036));
    InMux I__4886 (
            .O(N__22074),
            .I(N__22036));
    InMux I__4885 (
            .O(N__22073),
            .I(N__22036));
    InMux I__4884 (
            .O(N__22072),
            .I(N__22036));
    InMux I__4883 (
            .O(N__22071),
            .I(N__22033));
    LocalMux I__4882 (
            .O(N__22068),
            .I(N__22029));
    InMux I__4881 (
            .O(N__22067),
            .I(N__22026));
    LocalMux I__4880 (
            .O(N__22060),
            .I(N__22013));
    LocalMux I__4879 (
            .O(N__22057),
            .I(N__22013));
    LocalMux I__4878 (
            .O(N__22048),
            .I(N__22013));
    LocalMux I__4877 (
            .O(N__22045),
            .I(N__22006));
    LocalMux I__4876 (
            .O(N__22036),
            .I(N__22006));
    LocalMux I__4875 (
            .O(N__22033),
            .I(N__22006));
    InMux I__4874 (
            .O(N__22032),
            .I(N__22000));
    Span4Mux_s0_v I__4873 (
            .O(N__22029),
            .I(N__21995));
    LocalMux I__4872 (
            .O(N__22026),
            .I(N__21995));
    InMux I__4871 (
            .O(N__22025),
            .I(N__21984));
    InMux I__4870 (
            .O(N__22024),
            .I(N__21984));
    InMux I__4869 (
            .O(N__22023),
            .I(N__21984));
    InMux I__4868 (
            .O(N__22022),
            .I(N__21984));
    InMux I__4867 (
            .O(N__22021),
            .I(N__21984));
    InMux I__4866 (
            .O(N__22020),
            .I(N__21981));
    Span4Mux_s3_v I__4865 (
            .O(N__22013),
            .I(N__21978));
    Span4Mux_h I__4864 (
            .O(N__22006),
            .I(N__21975));
    InMux I__4863 (
            .O(N__22005),
            .I(N__21968));
    InMux I__4862 (
            .O(N__22004),
            .I(N__21968));
    InMux I__4861 (
            .O(N__22003),
            .I(N__21968));
    LocalMux I__4860 (
            .O(N__22000),
            .I(CO3_0));
    Odrv4 I__4859 (
            .O(N__21995),
            .I(CO3_0));
    LocalMux I__4858 (
            .O(N__21984),
            .I(CO3_0));
    LocalMux I__4857 (
            .O(N__21981),
            .I(CO3_0));
    Odrv4 I__4856 (
            .O(N__21978),
            .I(CO3_0));
    Odrv4 I__4855 (
            .O(N__21975),
            .I(CO3_0));
    LocalMux I__4854 (
            .O(N__21968),
            .I(CO3_0));
    CascadeMux I__4853 (
            .O(N__21953),
            .I(N__21950));
    InMux I__4852 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__4851 (
            .O(N__21947),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3_i));
    InMux I__4850 (
            .O(N__21944),
            .I(N__21940));
    InMux I__4849 (
            .O(N__21943),
            .I(N__21937));
    LocalMux I__4848 (
            .O(N__21940),
            .I(un113_pixel_1_0_3__N_10_mux));
    LocalMux I__4847 (
            .O(N__21937),
            .I(un113_pixel_1_0_3__N_10_mux));
    InMux I__4846 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__4845 (
            .O(N__21929),
            .I(beamY_RNIMR86ES2Z0Z_0));
    InMux I__4844 (
            .O(N__21926),
            .I(N__21923));
    LocalMux I__4843 (
            .O(N__21923),
            .I(N__21920));
    Odrv4 I__4842 (
            .O(N__21920),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254));
    InMux I__4841 (
            .O(N__21917),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__4840 (
            .O(N__21914),
            .I(N__21909));
    CascadeMux I__4839 (
            .O(N__21913),
            .I(N__21905));
    InMux I__4838 (
            .O(N__21912),
            .I(N__21901));
    InMux I__4837 (
            .O(N__21909),
            .I(N__21893));
    InMux I__4836 (
            .O(N__21908),
            .I(N__21893));
    InMux I__4835 (
            .O(N__21905),
            .I(N__21893));
    CascadeMux I__4834 (
            .O(N__21904),
            .I(N__21889));
    LocalMux I__4833 (
            .O(N__21901),
            .I(N__21884));
    CascadeMux I__4832 (
            .O(N__21900),
            .I(N__21881));
    LocalMux I__4831 (
            .O(N__21893),
            .I(N__21878));
    IoInMux I__4830 (
            .O(N__21892),
            .I(N__21875));
    InMux I__4829 (
            .O(N__21889),
            .I(N__21872));
    CascadeMux I__4828 (
            .O(N__21888),
            .I(N__21867));
    CascadeMux I__4827 (
            .O(N__21887),
            .I(N__21863));
    Span4Mux_v I__4826 (
            .O(N__21884),
            .I(N__21860));
    InMux I__4825 (
            .O(N__21881),
            .I(N__21857));
    IoSpan4Mux I__4824 (
            .O(N__21878),
            .I(N__21852));
    LocalMux I__4823 (
            .O(N__21875),
            .I(N__21852));
    LocalMux I__4822 (
            .O(N__21872),
            .I(N__21848));
    InMux I__4821 (
            .O(N__21871),
            .I(N__21845));
    CascadeMux I__4820 (
            .O(N__21870),
            .I(N__21841));
    InMux I__4819 (
            .O(N__21867),
            .I(N__21838));
    InMux I__4818 (
            .O(N__21866),
            .I(N__21833));
    InMux I__4817 (
            .O(N__21863),
            .I(N__21833));
    Span4Mux_v I__4816 (
            .O(N__21860),
            .I(N__21828));
    LocalMux I__4815 (
            .O(N__21857),
            .I(N__21828));
    IoSpan4Mux I__4814 (
            .O(N__21852),
            .I(N__21825));
    CascadeMux I__4813 (
            .O(N__21851),
            .I(N__21822));
    Span4Mux_s2_v I__4812 (
            .O(N__21848),
            .I(N__21819));
    LocalMux I__4811 (
            .O(N__21845),
            .I(N__21816));
    InMux I__4810 (
            .O(N__21844),
            .I(N__21811));
    InMux I__4809 (
            .O(N__21841),
            .I(N__21811));
    LocalMux I__4808 (
            .O(N__21838),
            .I(N__21808));
    LocalMux I__4807 (
            .O(N__21833),
            .I(N__21805));
    Span4Mux_h I__4806 (
            .O(N__21828),
            .I(N__21802));
    Span4Mux_s1_v I__4805 (
            .O(N__21825),
            .I(N__21799));
    InMux I__4804 (
            .O(N__21822),
            .I(N__21796));
    Sp12to4 I__4803 (
            .O(N__21819),
            .I(N__21789));
    Span12Mux_v I__4802 (
            .O(N__21816),
            .I(N__21789));
    LocalMux I__4801 (
            .O(N__21811),
            .I(N__21789));
    Odrv12 I__4800 (
            .O(N__21808),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4799 (
            .O(N__21805),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4798 (
            .O(N__21802),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4797 (
            .O(N__21799),
            .I(CONSTANT_ONE_NET));
    LocalMux I__4796 (
            .O(N__21796),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4795 (
            .O(N__21789),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4794 (
            .O(N__21776),
            .I(N__21773));
    InMux I__4793 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__4792 (
            .O(N__21770),
            .I(N__21767));
    Odrv4 I__4791 (
            .O(N__21767),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464));
    InMux I__4790 (
            .O(N__21764),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__4789 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__4788 (
            .O(N__21758),
            .I(N__21755));
    Odrv4 I__4787 (
            .O(N__21755),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO));
    InMux I__4786 (
            .O(N__21752),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__4785 (
            .O(N__21749),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7));
    CascadeMux I__4784 (
            .O(N__21746),
            .I(N__21743));
    InMux I__4783 (
            .O(N__21743),
            .I(N__21737));
    InMux I__4782 (
            .O(N__21742),
            .I(N__21737));
    LocalMux I__4781 (
            .O(N__21737),
            .I(N__21734));
    Odrv4 I__4780 (
            .O(N__21734),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    InMux I__4779 (
            .O(N__21731),
            .I(N__21728));
    LocalMux I__4778 (
            .O(N__21728),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf));
    InMux I__4777 (
            .O(N__21725),
            .I(N__21722));
    LocalMux I__4776 (
            .O(N__21722),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_2));
    InMux I__4775 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__4774 (
            .O(N__21716),
            .I(m17));
    InMux I__4773 (
            .O(N__21713),
            .I(N__21710));
    LocalMux I__4772 (
            .O(N__21710),
            .I(m12));
    InMux I__4771 (
            .O(N__21707),
            .I(N__21704));
    LocalMux I__4770 (
            .O(N__21704),
            .I(un115_pixel_5_ns_x1_0));
    InMux I__4769 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__4768 (
            .O(N__21698),
            .I(un115_pixel_5_ns_x0_0));
    CascadeMux I__4767 (
            .O(N__21695),
            .I(N_1325_cascade_));
    InMux I__4766 (
            .O(N__21692),
            .I(N__21689));
    LocalMux I__4765 (
            .O(N__21689),
            .I(N__21686));
    Span4Mux_v I__4764 (
            .O(N__21686),
            .I(N__21683));
    Odrv4 I__4763 (
            .O(N__21683),
            .I(un115_pixel_7_bm_0));
    CascadeMux I__4762 (
            .O(N__21680),
            .I(N_1315_cascade_));
    InMux I__4761 (
            .O(N__21677),
            .I(N__21674));
    LocalMux I__4760 (
            .O(N__21674),
            .I(N_1322));
    InMux I__4759 (
            .O(N__21671),
            .I(N__21668));
    LocalMux I__4758 (
            .O(N__21668),
            .I(N_1329));
    CascadeMux I__4757 (
            .O(N__21665),
            .I(N_1294_cascade_));
    InMux I__4756 (
            .O(N__21662),
            .I(N__21659));
    LocalMux I__4755 (
            .O(N__21659),
            .I(beamY_RNICJUESD2_1Z0Z_0));
    InMux I__4754 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__4753 (
            .O(N__21653),
            .I(N_1308));
    InMux I__4752 (
            .O(N__21650),
            .I(N__21647));
    LocalMux I__4751 (
            .O(N__21647),
            .I(un115_pixel_5_d_2));
    InMux I__4750 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__4749 (
            .O(N__21641),
            .I(N_1286_0_0_0));
    InMux I__4748 (
            .O(N__21638),
            .I(N__21635));
    LocalMux I__4747 (
            .O(N__21635),
            .I(N_1289));
    InMux I__4746 (
            .O(N__21632),
            .I(N__21629));
    LocalMux I__4745 (
            .O(N__21629),
            .I(N__21626));
    Span4Mux_v I__4744 (
            .O(N__21626),
            .I(N__21620));
    InMux I__4743 (
            .O(N__21625),
            .I(N__21615));
    InMux I__4742 (
            .O(N__21624),
            .I(N__21615));
    InMux I__4741 (
            .O(N__21623),
            .I(N__21612));
    Odrv4 I__4740 (
            .O(N__21620),
            .I(font_un3_pixel_29));
    LocalMux I__4739 (
            .O(N__21615),
            .I(font_un3_pixel_29));
    LocalMux I__4738 (
            .O(N__21612),
            .I(font_un3_pixel_29));
    CascadeMux I__4737 (
            .O(N__21605),
            .I(N_4562_0_0_0_cascade_));
    InMux I__4736 (
            .O(N__21602),
            .I(N__21599));
    LocalMux I__4735 (
            .O(N__21599),
            .I(N__21596));
    Odrv12 I__4734 (
            .O(N__21596),
            .I(N_1340_0));
    InMux I__4733 (
            .O(N__21593),
            .I(N__21590));
    LocalMux I__4732 (
            .O(N__21590),
            .I(beamY_RNICJUESD2_0Z0Z_0));
    InMux I__4731 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__4730 (
            .O(N__21584),
            .I(N__21581));
    Span4Mux_v I__4729 (
            .O(N__21581),
            .I(N__21578));
    Odrv4 I__4728 (
            .O(N__21578),
            .I(beamY_RNI1H36941Z0Z_0));
    InMux I__4727 (
            .O(N__21575),
            .I(N__21572));
    LocalMux I__4726 (
            .O(N__21572),
            .I(font_un125_pixel_1_bm));
    CascadeMux I__4725 (
            .O(N__21569),
            .I(un113_pixel_6_1_5__N_11_cascade_));
    InMux I__4724 (
            .O(N__21566),
            .I(N__21563));
    LocalMux I__4723 (
            .O(N__21563),
            .I(un113_pixel_2_0_3__N_8));
    InMux I__4722 (
            .O(N__21560),
            .I(N__21557));
    LocalMux I__4721 (
            .O(N__21557),
            .I(beamY_RNICJUESD2_2Z0Z_0));
    InMux I__4720 (
            .O(N__21554),
            .I(N__21551));
    LocalMux I__4719 (
            .O(N__21551),
            .I(un115_pixel_5_s_7));
    CascadeMux I__4718 (
            .O(N__21548),
            .I(un115_pixel_5_am_7_cascade_));
    InMux I__4717 (
            .O(N__21545),
            .I(N__21542));
    LocalMux I__4716 (
            .O(N__21542),
            .I(un115_pixel_5_bm_7));
    InMux I__4715 (
            .O(N__21539),
            .I(N__21536));
    LocalMux I__4714 (
            .O(N__21536),
            .I(N_1288));
    InMux I__4713 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__4712 (
            .O(N__21530),
            .I(N__21520));
    InMux I__4711 (
            .O(N__21529),
            .I(N__21517));
    InMux I__4710 (
            .O(N__21528),
            .I(N__21510));
    InMux I__4709 (
            .O(N__21527),
            .I(N__21510));
    InMux I__4708 (
            .O(N__21526),
            .I(N__21510));
    InMux I__4707 (
            .O(N__21525),
            .I(N__21503));
    InMux I__4706 (
            .O(N__21524),
            .I(N__21503));
    InMux I__4705 (
            .O(N__21523),
            .I(N__21503));
    Odrv4 I__4704 (
            .O(N__21520),
            .I(un113_pixel_3_0_11__currentchar_1_4Z0Z_2));
    LocalMux I__4703 (
            .O(N__21517),
            .I(un113_pixel_3_0_11__currentchar_1_4Z0Z_2));
    LocalMux I__4702 (
            .O(N__21510),
            .I(un113_pixel_3_0_11__currentchar_1_4Z0Z_2));
    LocalMux I__4701 (
            .O(N__21503),
            .I(un113_pixel_3_0_11__currentchar_1_4Z0Z_2));
    InMux I__4700 (
            .O(N__21494),
            .I(N__21491));
    LocalMux I__4699 (
            .O(N__21491),
            .I(N__21488));
    Span4Mux_s3_h I__4698 (
            .O(N__21488),
            .I(N__21485));
    Odrv4 I__4697 (
            .O(N__21485),
            .I(un113_pixel_4_0_15__g1Z0Z_0));
    InMux I__4696 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__4695 (
            .O(N__21479),
            .I(N__21476));
    Span4Mux_s3_h I__4694 (
            .O(N__21476),
            .I(N__21473));
    Odrv4 I__4693 (
            .O(N__21473),
            .I(m9));
    CascadeMux I__4692 (
            .O(N__21470),
            .I(m9_cascade_));
    InMux I__4691 (
            .O(N__21467),
            .I(N__21464));
    LocalMux I__4690 (
            .O(N__21464),
            .I(m6));
    CascadeMux I__4689 (
            .O(N__21461),
            .I(m6_cascade_));
    InMux I__4688 (
            .O(N__21458),
            .I(N__21455));
    LocalMux I__4687 (
            .O(N__21455),
            .I(N__21452));
    Odrv12 I__4686 (
            .O(N__21452),
            .I(beamY_RNICJUESD2Z0Z_0));
    CascadeMux I__4685 (
            .O(N__21449),
            .I(un115_pixel_2_s_6_cascade_));
    CascadeMux I__4684 (
            .O(N__21446),
            .I(un115_pixel_2_d_0_6_cascade_));
    InMux I__4683 (
            .O(N__21443),
            .I(N__21440));
    LocalMux I__4682 (
            .O(N__21440),
            .I(un115_pixel_3_bm_6));
    InMux I__4681 (
            .O(N__21437),
            .I(N__21433));
    InMux I__4680 (
            .O(N__21436),
            .I(N__21430));
    LocalMux I__4679 (
            .O(N__21433),
            .I(N__21425));
    LocalMux I__4678 (
            .O(N__21430),
            .I(N__21425));
    Odrv4 I__4677 (
            .O(N__21425),
            .I(ScreenBuffer_1_2Z0Z_1));
    InMux I__4676 (
            .O(N__21422),
            .I(N__21418));
    InMux I__4675 (
            .O(N__21421),
            .I(N__21415));
    LocalMux I__4674 (
            .O(N__21418),
            .I(ScreenBuffer_1_0Z0Z_1));
    LocalMux I__4673 (
            .O(N__21415),
            .I(ScreenBuffer_1_0Z0Z_1));
    InMux I__4672 (
            .O(N__21410),
            .I(N__21407));
    LocalMux I__4671 (
            .O(N__21407),
            .I(N_1_7_0));
    InMux I__4670 (
            .O(N__21404),
            .I(N__21400));
    InMux I__4669 (
            .O(N__21403),
            .I(N__21397));
    LocalMux I__4668 (
            .O(N__21400),
            .I(N__21392));
    LocalMux I__4667 (
            .O(N__21397),
            .I(N__21392));
    Span4Mux_v I__4666 (
            .O(N__21392),
            .I(N__21389));
    Odrv4 I__4665 (
            .O(N__21389),
            .I(ScreenBuffer_1_3Z0Z_1));
    InMux I__4664 (
            .O(N__21386),
            .I(N__21382));
    InMux I__4663 (
            .O(N__21385),
            .I(N__21379));
    LocalMux I__4662 (
            .O(N__21382),
            .I(N__21374));
    LocalMux I__4661 (
            .O(N__21379),
            .I(N__21374));
    Span4Mux_v I__4660 (
            .O(N__21374),
            .I(N__21371));
    Span4Mux_h I__4659 (
            .O(N__21371),
            .I(N__21368));
    Odrv4 I__4658 (
            .O(N__21368),
            .I(ScreenBuffer_1_1Z0Z_1));
    InMux I__4657 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__4656 (
            .O(N__21362),
            .I(m8));
    InMux I__4655 (
            .O(N__21359),
            .I(N__21356));
    LocalMux I__4654 (
            .O(N__21356),
            .I(N__21352));
    InMux I__4653 (
            .O(N__21355),
            .I(N__21349));
    Span4Mux_h I__4652 (
            .O(N__21352),
            .I(N__21346));
    LocalMux I__4651 (
            .O(N__21349),
            .I(ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1));
    Odrv4 I__4650 (
            .O(N__21346),
            .I(ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1));
    InMux I__4649 (
            .O(N__21341),
            .I(N__21337));
    InMux I__4648 (
            .O(N__21340),
            .I(N__21334));
    LocalMux I__4647 (
            .O(N__21337),
            .I(N__21331));
    LocalMux I__4646 (
            .O(N__21334),
            .I(ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1));
    Odrv4 I__4645 (
            .O(N__21331),
            .I(ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1));
    InMux I__4644 (
            .O(N__21326),
            .I(N__21317));
    InMux I__4643 (
            .O(N__21325),
            .I(N__21317));
    InMux I__4642 (
            .O(N__21324),
            .I(N__21317));
    LocalMux I__4641 (
            .O(N__21317),
            .I(N__21313));
    InMux I__4640 (
            .O(N__21316),
            .I(N__21310));
    Odrv4 I__4639 (
            .O(N__21313),
            .I(ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1));
    LocalMux I__4638 (
            .O(N__21310),
            .I(ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1));
    CascadeMux I__4637 (
            .O(N__21305),
            .I(ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_));
    InMux I__4636 (
            .O(N__21302),
            .I(N__21299));
    LocalMux I__4635 (
            .O(N__21299),
            .I(un113_pixel_3_0_11__gZ0Z1));
    InMux I__4634 (
            .O(N__21296),
            .I(N__21293));
    LocalMux I__4633 (
            .O(N__21293),
            .I(N__21290));
    Span4Mux_v I__4632 (
            .O(N__21290),
            .I(N__21286));
    InMux I__4631 (
            .O(N__21289),
            .I(N__21283));
    Odrv4 I__4630 (
            .O(N__21286),
            .I(font_un3_pixel_28));
    LocalMux I__4629 (
            .O(N__21283),
            .I(font_un3_pixel_28));
    CascadeMux I__4628 (
            .O(N__21278),
            .I(N__21275));
    InMux I__4627 (
            .O(N__21275),
            .I(N__21272));
    LocalMux I__4626 (
            .O(N__21272),
            .I(N_1342));
    InMux I__4625 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__4624 (
            .O(N__21266),
            .I(N__21263));
    Odrv12 I__4623 (
            .O(N__21263),
            .I(un113_pixel_4_0_15__g0_5Z0Z_1));
    InMux I__4622 (
            .O(N__21260),
            .I(N__21255));
    InMux I__4621 (
            .O(N__21259),
            .I(N__21250));
    InMux I__4620 (
            .O(N__21258),
            .I(N__21250));
    LocalMux I__4619 (
            .O(N__21255),
            .I(font_un71_pixellt7_0_1));
    LocalMux I__4618 (
            .O(N__21250),
            .I(font_un71_pixellt7_0_1));
    CascadeMux I__4617 (
            .O(N__21245),
            .I(N__21242));
    InMux I__4616 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__4615 (
            .O(N__21239),
            .I(font_un64_pixel_ac0_5_0));
    InMux I__4614 (
            .O(N__21236),
            .I(N__21232));
    InMux I__4613 (
            .O(N__21235),
            .I(N__21229));
    LocalMux I__4612 (
            .O(N__21232),
            .I(N__21226));
    LocalMux I__4611 (
            .O(N__21229),
            .I(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3));
    Odrv4 I__4610 (
            .O(N__21226),
            .I(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3));
    InMux I__4609 (
            .O(N__21221),
            .I(N__21218));
    LocalMux I__4608 (
            .O(N__21218),
            .I(N__21215));
    Span4Mux_h I__4607 (
            .O(N__21215),
            .I(N__21212));
    Odrv4 I__4606 (
            .O(N__21212),
            .I(font_un3_pixel_0_29));
    CascadeMux I__4605 (
            .O(N__21209),
            .I(un113_pixel_4_0_15__g0_5Z0Z_4_cascade_));
    InMux I__4604 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__4603 (
            .O(N__21203),
            .I(N_9));
    CascadeMux I__4602 (
            .O(N__21200),
            .I(un113_pixel_4_0_15__g2Z0Z_0_cascade_));
    InMux I__4601 (
            .O(N__21197),
            .I(N__21194));
    LocalMux I__4600 (
            .O(N__21194),
            .I(N__21191));
    Span4Mux_h I__4599 (
            .O(N__21191),
            .I(N__21188));
    Odrv4 I__4598 (
            .O(N__21188),
            .I(N_4566_0));
    InMux I__4597 (
            .O(N__21185),
            .I(N__21182));
    LocalMux I__4596 (
            .O(N__21182),
            .I(un115_pixel_4));
    InMux I__4595 (
            .O(N__21179),
            .I(N__21176));
    LocalMux I__4594 (
            .O(N__21176),
            .I(N_4564_0));
    InMux I__4593 (
            .O(N__21173),
            .I(N__21170));
    LocalMux I__4592 (
            .O(N__21170),
            .I(N_5_0));
    InMux I__4591 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__4590 (
            .O(N__21164),
            .I(N__21160));
    CascadeMux I__4589 (
            .O(N__21163),
            .I(N__21154));
    Span4Mux_h I__4588 (
            .O(N__21160),
            .I(N__21151));
    InMux I__4587 (
            .O(N__21159),
            .I(N__21148));
    InMux I__4586 (
            .O(N__21158),
            .I(N__21141));
    InMux I__4585 (
            .O(N__21157),
            .I(N__21141));
    InMux I__4584 (
            .O(N__21154),
            .I(N__21141));
    Odrv4 I__4583 (
            .O(N__21151),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1));
    LocalMux I__4582 (
            .O(N__21148),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1));
    LocalMux I__4581 (
            .O(N__21141),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1));
    InMux I__4580 (
            .O(N__21134),
            .I(N__21131));
    LocalMux I__4579 (
            .O(N__21131),
            .I(N__21128));
    Span4Mux_s3_h I__4578 (
            .O(N__21128),
            .I(N__21125));
    Odrv4 I__4577 (
            .O(N__21125),
            .I(N_4561_0));
    CascadeMux I__4576 (
            .O(N__21122),
            .I(N__21119));
    InMux I__4575 (
            .O(N__21119),
            .I(N__21116));
    LocalMux I__4574 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_v I__4573 (
            .O(N__21113),
            .I(N__21110));
    Span4Mux_s3_h I__4572 (
            .O(N__21110),
            .I(N__21107));
    Odrv4 I__4571 (
            .O(N__21107),
            .I(g1_0));
    CascadeMux I__4570 (
            .O(N__21104),
            .I(N__21101));
    InMux I__4569 (
            .O(N__21101),
            .I(N__21098));
    LocalMux I__4568 (
            .O(N__21098),
            .I(N_2075));
    InMux I__4567 (
            .O(N__21095),
            .I(N__21092));
    LocalMux I__4566 (
            .O(N__21092),
            .I(N__21089));
    Span4Mux_v I__4565 (
            .O(N__21089),
            .I(N__21086));
    Odrv4 I__4564 (
            .O(N__21086),
            .I(N_11));
    InMux I__4563 (
            .O(N__21083),
            .I(N__21080));
    LocalMux I__4562 (
            .O(N__21080),
            .I(un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0));
    InMux I__4561 (
            .O(N__21077),
            .I(N__21074));
    LocalMux I__4560 (
            .O(N__21074),
            .I(un113_pixel_4_0_15__g0_i_a3_2));
    IoInMux I__4559 (
            .O(N__21071),
            .I(N__21068));
    LocalMux I__4558 (
            .O(N__21068),
            .I(N__21065));
    Odrv12 I__4557 (
            .O(N__21065),
            .I(Pixel_c));
    ClkMux I__4556 (
            .O(N__21062),
            .I(N__21029));
    ClkMux I__4555 (
            .O(N__21061),
            .I(N__21029));
    ClkMux I__4554 (
            .O(N__21060),
            .I(N__21029));
    ClkMux I__4553 (
            .O(N__21059),
            .I(N__21029));
    ClkMux I__4552 (
            .O(N__21058),
            .I(N__21029));
    ClkMux I__4551 (
            .O(N__21057),
            .I(N__21029));
    ClkMux I__4550 (
            .O(N__21056),
            .I(N__21029));
    ClkMux I__4549 (
            .O(N__21055),
            .I(N__21029));
    ClkMux I__4548 (
            .O(N__21054),
            .I(N__21029));
    ClkMux I__4547 (
            .O(N__21053),
            .I(N__21029));
    ClkMux I__4546 (
            .O(N__21052),
            .I(N__21029));
    GlobalMux I__4545 (
            .O(N__21029),
            .I(N__21026));
    gio2CtrlBuf I__4544 (
            .O(N__21026),
            .I(PixelClock_g));
    InMux I__4543 (
            .O(N__21023),
            .I(N__21020));
    LocalMux I__4542 (
            .O(N__21020),
            .I(N__21017));
    Odrv12 I__4541 (
            .O(N__21017),
            .I(un113_pixel_7_1_7__g0_6Z0Z_0));
    CascadeMux I__4540 (
            .O(N__21014),
            .I(N__21011));
    InMux I__4539 (
            .O(N__21011),
            .I(N__21008));
    LocalMux I__4538 (
            .O(N__21008),
            .I(N__21005));
    Sp12to4 I__4537 (
            .O(N__21005),
            .I(N__21002));
    Odrv12 I__4536 (
            .O(N__21002),
            .I(N_3078_0));
    CascadeMux I__4535 (
            .O(N__20999),
            .I(N_1297_0_cascade_));
    InMux I__4534 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__4533 (
            .O(N__20993),
            .I(N__20990));
    Span4Mux_v I__4532 (
            .O(N__20990),
            .I(N__20987));
    Odrv4 I__4531 (
            .O(N__20987),
            .I(font_un67_pixel_ac0_5_0));
    InMux I__4530 (
            .O(N__20984),
            .I(N__20978));
    InMux I__4529 (
            .O(N__20983),
            .I(N__20975));
    InMux I__4528 (
            .O(N__20982),
            .I(N__20970));
    InMux I__4527 (
            .O(N__20981),
            .I(N__20970));
    LocalMux I__4526 (
            .O(N__20978),
            .I(N__20967));
    LocalMux I__4525 (
            .O(N__20975),
            .I(N__20963));
    LocalMux I__4524 (
            .O(N__20970),
            .I(N__20960));
    Span4Mux_h I__4523 (
            .O(N__20967),
            .I(N__20957));
    InMux I__4522 (
            .O(N__20966),
            .I(N__20954));
    Span4Mux_h I__4521 (
            .O(N__20963),
            .I(N__20951));
    Span4Mux_h I__4520 (
            .O(N__20960),
            .I(N__20948));
    Odrv4 I__4519 (
            .O(N__20957),
            .I(chary_if_generate_plus_mult1_un68_sum_c5));
    LocalMux I__4518 (
            .O(N__20954),
            .I(chary_if_generate_plus_mult1_un68_sum_c5));
    Odrv4 I__4517 (
            .O(N__20951),
            .I(chary_if_generate_plus_mult1_un68_sum_c5));
    Odrv4 I__4516 (
            .O(N__20948),
            .I(chary_if_generate_plus_mult1_un68_sum_c5));
    InMux I__4515 (
            .O(N__20939),
            .I(N__20936));
    LocalMux I__4514 (
            .O(N__20936),
            .I(N__20930));
    InMux I__4513 (
            .O(N__20935),
            .I(N__20925));
    InMux I__4512 (
            .O(N__20934),
            .I(N__20925));
    InMux I__4511 (
            .O(N__20933),
            .I(N__20921));
    Span4Mux_s3_h I__4510 (
            .O(N__20930),
            .I(N__20916));
    LocalMux I__4509 (
            .O(N__20925),
            .I(N__20916));
    InMux I__4508 (
            .O(N__20924),
            .I(N__20913));
    LocalMux I__4507 (
            .O(N__20921),
            .I(N__20910));
    Span4Mux_h I__4506 (
            .O(N__20916),
            .I(N__20907));
    LocalMux I__4505 (
            .O(N__20913),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_2));
    Odrv12 I__4504 (
            .O(N__20910),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_2));
    Odrv4 I__4503 (
            .O(N__20907),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_2));
    InMux I__4502 (
            .O(N__20900),
            .I(N__20897));
    LocalMux I__4501 (
            .O(N__20897),
            .I(un113_pixel_4_0_15__g0_4_0Z0Z_0));
    CascadeMux I__4500 (
            .O(N__20894),
            .I(N__20889));
    CascadeMux I__4499 (
            .O(N__20893),
            .I(N__20879));
    InMux I__4498 (
            .O(N__20892),
            .I(N__20876));
    InMux I__4497 (
            .O(N__20889),
            .I(N__20873));
    InMux I__4496 (
            .O(N__20888),
            .I(N__20866));
    InMux I__4495 (
            .O(N__20887),
            .I(N__20866));
    InMux I__4494 (
            .O(N__20886),
            .I(N__20866));
    CascadeMux I__4493 (
            .O(N__20885),
            .I(N__20862));
    CascadeMux I__4492 (
            .O(N__20884),
            .I(N__20859));
    InMux I__4491 (
            .O(N__20883),
            .I(N__20855));
    InMux I__4490 (
            .O(N__20882),
            .I(N__20850));
    InMux I__4489 (
            .O(N__20879),
            .I(N__20850));
    LocalMux I__4488 (
            .O(N__20876),
            .I(N__20847));
    LocalMux I__4487 (
            .O(N__20873),
            .I(N__20842));
    LocalMux I__4486 (
            .O(N__20866),
            .I(N__20842));
    InMux I__4485 (
            .O(N__20865),
            .I(N__20833));
    InMux I__4484 (
            .O(N__20862),
            .I(N__20833));
    InMux I__4483 (
            .O(N__20859),
            .I(N__20833));
    CascadeMux I__4482 (
            .O(N__20858),
            .I(N__20828));
    LocalMux I__4481 (
            .O(N__20855),
            .I(N__20822));
    LocalMux I__4480 (
            .O(N__20850),
            .I(N__20819));
    Span4Mux_v I__4479 (
            .O(N__20847),
            .I(N__20816));
    Span4Mux_h I__4478 (
            .O(N__20842),
            .I(N__20813));
    InMux I__4477 (
            .O(N__20841),
            .I(N__20810));
    InMux I__4476 (
            .O(N__20840),
            .I(N__20807));
    LocalMux I__4475 (
            .O(N__20833),
            .I(N__20804));
    InMux I__4474 (
            .O(N__20832),
            .I(N__20801));
    InMux I__4473 (
            .O(N__20831),
            .I(N__20798));
    InMux I__4472 (
            .O(N__20828),
            .I(N__20791));
    InMux I__4471 (
            .O(N__20827),
            .I(N__20791));
    InMux I__4470 (
            .O(N__20826),
            .I(N__20791));
    InMux I__4469 (
            .O(N__20825),
            .I(N__20786));
    Span4Mux_v I__4468 (
            .O(N__20822),
            .I(N__20783));
    Span4Mux_v I__4467 (
            .O(N__20819),
            .I(N__20780));
    Span4Mux_h I__4466 (
            .O(N__20816),
            .I(N__20773));
    Span4Mux_v I__4465 (
            .O(N__20813),
            .I(N__20773));
    LocalMux I__4464 (
            .O(N__20810),
            .I(N__20773));
    LocalMux I__4463 (
            .O(N__20807),
            .I(N__20770));
    Span4Mux_v I__4462 (
            .O(N__20804),
            .I(N__20767));
    LocalMux I__4461 (
            .O(N__20801),
            .I(N__20764));
    LocalMux I__4460 (
            .O(N__20798),
            .I(N__20759));
    LocalMux I__4459 (
            .O(N__20791),
            .I(N__20759));
    InMux I__4458 (
            .O(N__20790),
            .I(N__20756));
    InMux I__4457 (
            .O(N__20789),
            .I(N__20748));
    LocalMux I__4456 (
            .O(N__20786),
            .I(N__20745));
    Span4Mux_h I__4455 (
            .O(N__20783),
            .I(N__20742));
    Span4Mux_h I__4454 (
            .O(N__20780),
            .I(N__20739));
    Span4Mux_h I__4453 (
            .O(N__20773),
            .I(N__20736));
    Span4Mux_v I__4452 (
            .O(N__20770),
            .I(N__20725));
    Span4Mux_h I__4451 (
            .O(N__20767),
            .I(N__20725));
    Span4Mux_v I__4450 (
            .O(N__20764),
            .I(N__20725));
    Span4Mux_v I__4449 (
            .O(N__20759),
            .I(N__20725));
    LocalMux I__4448 (
            .O(N__20756),
            .I(N__20725));
    InMux I__4447 (
            .O(N__20755),
            .I(N__20720));
    InMux I__4446 (
            .O(N__20754),
            .I(N__20720));
    InMux I__4445 (
            .O(N__20753),
            .I(N__20717));
    InMux I__4444 (
            .O(N__20752),
            .I(N__20712));
    InMux I__4443 (
            .O(N__20751),
            .I(N__20712));
    LocalMux I__4442 (
            .O(N__20748),
            .I(beamYZ0Z_2));
    Odrv4 I__4441 (
            .O(N__20745),
            .I(beamYZ0Z_2));
    Odrv4 I__4440 (
            .O(N__20742),
            .I(beamYZ0Z_2));
    Odrv4 I__4439 (
            .O(N__20739),
            .I(beamYZ0Z_2));
    Odrv4 I__4438 (
            .O(N__20736),
            .I(beamYZ0Z_2));
    Odrv4 I__4437 (
            .O(N__20725),
            .I(beamYZ0Z_2));
    LocalMux I__4436 (
            .O(N__20720),
            .I(beamYZ0Z_2));
    LocalMux I__4435 (
            .O(N__20717),
            .I(beamYZ0Z_2));
    LocalMux I__4434 (
            .O(N__20712),
            .I(beamYZ0Z_2));
    InMux I__4433 (
            .O(N__20693),
            .I(N__20682));
    InMux I__4432 (
            .O(N__20692),
            .I(N__20682));
    InMux I__4431 (
            .O(N__20691),
            .I(N__20682));
    CascadeMux I__4430 (
            .O(N__20690),
            .I(N__20679));
    InMux I__4429 (
            .O(N__20689),
            .I(N__20673));
    LocalMux I__4428 (
            .O(N__20682),
            .I(N__20669));
    InMux I__4427 (
            .O(N__20679),
            .I(N__20664));
    InMux I__4426 (
            .O(N__20678),
            .I(N__20664));
    InMux I__4425 (
            .O(N__20677),
            .I(N__20659));
    InMux I__4424 (
            .O(N__20676),
            .I(N__20659));
    LocalMux I__4423 (
            .O(N__20673),
            .I(N__20656));
    InMux I__4422 (
            .O(N__20672),
            .I(N__20653));
    Span4Mux_s3_h I__4421 (
            .O(N__20669),
            .I(N__20648));
    LocalMux I__4420 (
            .O(N__20664),
            .I(N__20648));
    LocalMux I__4419 (
            .O(N__20659),
            .I(N__20641));
    Span4Mux_v I__4418 (
            .O(N__20656),
            .I(N__20641));
    LocalMux I__4417 (
            .O(N__20653),
            .I(N__20641));
    Span4Mux_h I__4416 (
            .O(N__20648),
            .I(N__20638));
    Odrv4 I__4415 (
            .O(N__20641),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i));
    Odrv4 I__4414 (
            .O(N__20638),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i));
    CascadeMux I__4413 (
            .O(N__20633),
            .I(un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_));
    CascadeMux I__4412 (
            .O(N__20630),
            .I(N__20627));
    InMux I__4411 (
            .O(N__20627),
            .I(N__20624));
    LocalMux I__4410 (
            .O(N__20624),
            .I(charx_if_generate_plus_mult1_un61_sum_i));
    InMux I__4409 (
            .O(N__20621),
            .I(N__20616));
    InMux I__4408 (
            .O(N__20620),
            .I(N__20613));
    InMux I__4407 (
            .O(N__20619),
            .I(N__20610));
    LocalMux I__4406 (
            .O(N__20616),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0));
    LocalMux I__4405 (
            .O(N__20613),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0));
    LocalMux I__4404 (
            .O(N__20610),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0));
    InMux I__4403 (
            .O(N__20603),
            .I(N__20597));
    InMux I__4402 (
            .O(N__20602),
            .I(N__20597));
    LocalMux I__4401 (
            .O(N__20597),
            .I(charx_if_generate_plus_mult1_un61_sum_i_5));
    InMux I__4400 (
            .O(N__20594),
            .I(N__20591));
    LocalMux I__4399 (
            .O(N__20591),
            .I(N_2096_i));
    CascadeMux I__4398 (
            .O(N__20588),
            .I(N__20585));
    InMux I__4397 (
            .O(N__20585),
            .I(N__20582));
    LocalMux I__4396 (
            .O(N__20582),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__4395 (
            .O(N__20579),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__4394 (
            .O(N__20576),
            .I(N__20573));
    LocalMux I__4393 (
            .O(N__20573),
            .I(N__20569));
    InMux I__4392 (
            .O(N__20572),
            .I(N__20566));
    Span4Mux_v I__4391 (
            .O(N__20569),
            .I(N__20562));
    LocalMux I__4390 (
            .O(N__20566),
            .I(N__20559));
    InMux I__4389 (
            .O(N__20565),
            .I(N__20556));
    Odrv4 I__4388 (
            .O(N__20562),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    Odrv4 I__4387 (
            .O(N__20559),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__4386 (
            .O(N__20556),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    CascadeMux I__4385 (
            .O(N__20549),
            .I(N__20546));
    InMux I__4384 (
            .O(N__20546),
            .I(N__20543));
    LocalMux I__4383 (
            .O(N__20543),
            .I(N__20540));
    Odrv12 I__4382 (
            .O(N__20540),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    CascadeMux I__4381 (
            .O(N__20537),
            .I(N__20534));
    InMux I__4380 (
            .O(N__20534),
            .I(N__20531));
    LocalMux I__4379 (
            .O(N__20531),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__4378 (
            .O(N__20528),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__4377 (
            .O(N__20525),
            .I(N__20521));
    InMux I__4376 (
            .O(N__20524),
            .I(N__20518));
    InMux I__4375 (
            .O(N__20521),
            .I(N__20515));
    LocalMux I__4374 (
            .O(N__20518),
            .I(N__20510));
    LocalMux I__4373 (
            .O(N__20515),
            .I(N__20510));
    Odrv4 I__4372 (
            .O(N__20510),
            .I(column_1_if_generate_plus_mult1_un54_sum_i_5));
    CascadeMux I__4371 (
            .O(N__20507),
            .I(N__20504));
    InMux I__4370 (
            .O(N__20504),
            .I(N__20501));
    LocalMux I__4369 (
            .O(N__20501),
            .I(N__20498));
    Odrv4 I__4368 (
            .O(N__20498),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__4367 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__4366 (
            .O(N__20492),
            .I(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__4365 (
            .O(N__20489),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__4364 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__4363 (
            .O(N__20483),
            .I(N__20480));
    Odrv4 I__4362 (
            .O(N__20480),
            .I(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__4361 (
            .O(N__20477),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__4360 (
            .O(N__20474),
            .I(N__20468));
    InMux I__4359 (
            .O(N__20473),
            .I(N__20468));
    LocalMux I__4358 (
            .O(N__20468),
            .I(column_1_i_i_3));
    InMux I__4357 (
            .O(N__20465),
            .I(N__20459));
    InMux I__4356 (
            .O(N__20464),
            .I(N__20459));
    LocalMux I__4355 (
            .O(N__20459),
            .I(charx_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__4354 (
            .O(N__20456),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__4353 (
            .O(N__20453),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__4352 (
            .O(N__20450),
            .I(N__20447));
    InMux I__4351 (
            .O(N__20447),
            .I(N__20444));
    LocalMux I__4350 (
            .O(N__20444),
            .I(charx_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__4349 (
            .O(N__20441),
            .I(N__20438));
    InMux I__4348 (
            .O(N__20438),
            .I(N__20435));
    LocalMux I__4347 (
            .O(N__20435),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0));
    InMux I__4346 (
            .O(N__20432),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__4345 (
            .O(N__20429),
            .I(N__20426));
    InMux I__4344 (
            .O(N__20426),
            .I(N__20423));
    LocalMux I__4343 (
            .O(N__20423),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8));
    CascadeMux I__4342 (
            .O(N__20420),
            .I(N__20417));
    InMux I__4341 (
            .O(N__20417),
            .I(N__20414));
    LocalMux I__4340 (
            .O(N__20414),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0));
    InMux I__4339 (
            .O(N__20411),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2));
    CascadeMux I__4338 (
            .O(N__20408),
            .I(N__20405));
    InMux I__4337 (
            .O(N__20405),
            .I(N__20402));
    LocalMux I__4336 (
            .O(N__20402),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0));
    InMux I__4335 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__4334 (
            .O(N__20396),
            .I(charx_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__4333 (
            .O(N__20393),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__4332 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__4331 (
            .O(N__20387),
            .I(charx_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__4330 (
            .O(N__20384),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__4329 (
            .O(N__20381),
            .I(N__20376));
    InMux I__4328 (
            .O(N__20380),
            .I(N__20373));
    InMux I__4327 (
            .O(N__20379),
            .I(N__20370));
    LocalMux I__4326 (
            .O(N__20376),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0));
    LocalMux I__4325 (
            .O(N__20373),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0));
    LocalMux I__4324 (
            .O(N__20370),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0));
    InMux I__4323 (
            .O(N__20363),
            .I(N__20360));
    LocalMux I__4322 (
            .O(N__20360),
            .I(N__20357));
    Odrv4 I__4321 (
            .O(N__20357),
            .I(if_generate_plus_mult1_un54_sum_axb_2_l_fx));
    InMux I__4320 (
            .O(N__20354),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__4319 (
            .O(N__20351),
            .I(N__20345));
    CascadeMux I__4318 (
            .O(N__20350),
            .I(N__20341));
    CascadeMux I__4317 (
            .O(N__20349),
            .I(N__20338));
    InMux I__4316 (
            .O(N__20348),
            .I(N__20334));
    LocalMux I__4315 (
            .O(N__20345),
            .I(N__20331));
    InMux I__4314 (
            .O(N__20344),
            .I(N__20328));
    InMux I__4313 (
            .O(N__20341),
            .I(N__20321));
    InMux I__4312 (
            .O(N__20338),
            .I(N__20321));
    InMux I__4311 (
            .O(N__20337),
            .I(N__20321));
    LocalMux I__4310 (
            .O(N__20334),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    Odrv4 I__4309 (
            .O(N__20331),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    LocalMux I__4308 (
            .O(N__20328),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    LocalMux I__4307 (
            .O(N__20321),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    CascadeMux I__4306 (
            .O(N__20312),
            .I(N__20309));
    InMux I__4305 (
            .O(N__20309),
            .I(N__20306));
    LocalMux I__4304 (
            .O(N__20306),
            .I(N__20303));
    Odrv4 I__4303 (
            .O(N__20303),
            .I(if_generate_plus_mult1_un54_sum_axb_3_l_fx));
    InMux I__4302 (
            .O(N__20300),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__4301 (
            .O(N__20297),
            .I(N__20294));
    LocalMux I__4300 (
            .O(N__20294),
            .I(if_generate_plus_mult1_un54_sum_axb_4_l_fx));
    CascadeMux I__4299 (
            .O(N__20291),
            .I(N__20287));
    CascadeMux I__4298 (
            .O(N__20290),
            .I(N__20284));
    InMux I__4297 (
            .O(N__20287),
            .I(N__20279));
    InMux I__4296 (
            .O(N__20284),
            .I(N__20279));
    LocalMux I__4295 (
            .O(N__20279),
            .I(N__20275));
    InMux I__4294 (
            .O(N__20278),
            .I(N__20272));
    Odrv4 I__4293 (
            .O(N__20275),
            .I(N_2110_i));
    LocalMux I__4292 (
            .O(N__20272),
            .I(N_2110_i));
    InMux I__4291 (
            .O(N__20267),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__4290 (
            .O(N__20264),
            .I(N__20261));
    LocalMux I__4289 (
            .O(N__20261),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__4288 (
            .O(N__20258),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__4287 (
            .O(N__20255),
            .I(if_generate_plus_mult1_un54_sum_s_5_cascade_));
    InMux I__4286 (
            .O(N__20252),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__4285 (
            .O(N__20249),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__4284 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__4283 (
            .O(N__20243),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2));
    InMux I__4282 (
            .O(N__20240),
            .I(N__20237));
    LocalMux I__4281 (
            .O(N__20237),
            .I(column_1_if_generate_plus_mult1_un47_sum0_3));
    CascadeMux I__4280 (
            .O(N__20234),
            .I(N__20231));
    InMux I__4279 (
            .O(N__20231),
            .I(N__20228));
    LocalMux I__4278 (
            .O(N__20228),
            .I(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx));
    InMux I__4277 (
            .O(N__20225),
            .I(N__20222));
    LocalMux I__4276 (
            .O(N__20222),
            .I(column_1_if_generate_plus_mult1_un47_sum0_2));
    InMux I__4275 (
            .O(N__20219),
            .I(N__20211));
    InMux I__4274 (
            .O(N__20218),
            .I(N__20211));
    InMux I__4273 (
            .O(N__20217),
            .I(N__20200));
    InMux I__4272 (
            .O(N__20216),
            .I(N__20196));
    LocalMux I__4271 (
            .O(N__20211),
            .I(N__20190));
    InMux I__4270 (
            .O(N__20210),
            .I(N__20187));
    InMux I__4269 (
            .O(N__20209),
            .I(N__20178));
    InMux I__4268 (
            .O(N__20208),
            .I(N__20178));
    InMux I__4267 (
            .O(N__20207),
            .I(N__20178));
    InMux I__4266 (
            .O(N__20206),
            .I(N__20178));
    InMux I__4265 (
            .O(N__20205),
            .I(N__20175));
    InMux I__4264 (
            .O(N__20204),
            .I(N__20170));
    InMux I__4263 (
            .O(N__20203),
            .I(N__20170));
    LocalMux I__4262 (
            .O(N__20200),
            .I(N__20167));
    InMux I__4261 (
            .O(N__20199),
            .I(N__20164));
    LocalMux I__4260 (
            .O(N__20196),
            .I(N__20158));
    InMux I__4259 (
            .O(N__20195),
            .I(N__20155));
    InMux I__4258 (
            .O(N__20194),
            .I(N__20150));
    InMux I__4257 (
            .O(N__20193),
            .I(N__20150));
    Span4Mux_h I__4256 (
            .O(N__20190),
            .I(N__20145));
    LocalMux I__4255 (
            .O(N__20187),
            .I(N__20145));
    LocalMux I__4254 (
            .O(N__20178),
            .I(N__20142));
    LocalMux I__4253 (
            .O(N__20175),
            .I(N__20137));
    LocalMux I__4252 (
            .O(N__20170),
            .I(N__20137));
    Span4Mux_s1_h I__4251 (
            .O(N__20167),
            .I(N__20132));
    LocalMux I__4250 (
            .O(N__20164),
            .I(N__20132));
    InMux I__4249 (
            .O(N__20163),
            .I(N__20125));
    InMux I__4248 (
            .O(N__20162),
            .I(N__20125));
    InMux I__4247 (
            .O(N__20161),
            .I(N__20125));
    Sp12to4 I__4246 (
            .O(N__20158),
            .I(N__20122));
    LocalMux I__4245 (
            .O(N__20155),
            .I(N__20117));
    LocalMux I__4244 (
            .O(N__20150),
            .I(N__20117));
    Span4Mux_v I__4243 (
            .O(N__20145),
            .I(N__20114));
    Span4Mux_v I__4242 (
            .O(N__20142),
            .I(N__20111));
    Span4Mux_v I__4241 (
            .O(N__20137),
            .I(N__20104));
    Span4Mux_h I__4240 (
            .O(N__20132),
            .I(N__20104));
    LocalMux I__4239 (
            .O(N__20125),
            .I(N__20104));
    Span12Mux_v I__4238 (
            .O(N__20122),
            .I(N__20099));
    Span12Mux_s9_h I__4237 (
            .O(N__20117),
            .I(N__20099));
    IoSpan4Mux I__4236 (
            .O(N__20114),
            .I(N__20096));
    Span4Mux_h I__4235 (
            .O(N__20111),
            .I(N__20091));
    Span4Mux_h I__4234 (
            .O(N__20104),
            .I(N__20091));
    Odrv12 I__4233 (
            .O(N__20099),
            .I(SDATA1_c));
    Odrv4 I__4232 (
            .O(N__20096),
            .I(SDATA1_c));
    Odrv4 I__4231 (
            .O(N__20091),
            .I(SDATA1_c));
    InMux I__4230 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__4229 (
            .O(N__20081),
            .I(N__20078));
    Span4Mux_v I__4228 (
            .O(N__20078),
            .I(N__20075));
    Span4Mux_v I__4227 (
            .O(N__20075),
            .I(N__20071));
    InMux I__4226 (
            .O(N__20074),
            .I(N__20068));
    Span4Mux_v I__4225 (
            .O(N__20071),
            .I(N__20063));
    LocalMux I__4224 (
            .O(N__20068),
            .I(N__20063));
    Span4Mux_h I__4223 (
            .O(N__20063),
            .I(N__20058));
    InMux I__4222 (
            .O(N__20062),
            .I(N__20052));
    InMux I__4221 (
            .O(N__20061),
            .I(N__20052));
    Span4Mux_h I__4220 (
            .O(N__20058),
            .I(N__20049));
    InMux I__4219 (
            .O(N__20057),
            .I(N__20046));
    LocalMux I__4218 (
            .O(N__20052),
            .I(un1_sclk17_9_0_3));
    Odrv4 I__4217 (
            .O(N__20049),
            .I(un1_sclk17_9_0_3));
    LocalMux I__4216 (
            .O(N__20046),
            .I(un1_sclk17_9_0_3));
    CascadeMux I__4215 (
            .O(N__20039),
            .I(N__20036));
    InMux I__4214 (
            .O(N__20036),
            .I(N__20033));
    LocalMux I__4213 (
            .O(N__20033),
            .I(N__20030));
    Span4Mux_v I__4212 (
            .O(N__20030),
            .I(N__20027));
    Span4Mux_v I__4211 (
            .O(N__20027),
            .I(N__20024));
    Span4Mux_h I__4210 (
            .O(N__20024),
            .I(N__20021));
    Odrv4 I__4209 (
            .O(N__20021),
            .I(un1_sclk17_5_1_0));
    InMux I__4208 (
            .O(N__20018),
            .I(N__20015));
    LocalMux I__4207 (
            .O(N__20015),
            .I(N__20012));
    Span4Mux_h I__4206 (
            .O(N__20012),
            .I(N__20008));
    InMux I__4205 (
            .O(N__20011),
            .I(N__20005));
    Span4Mux_v I__4204 (
            .O(N__20008),
            .I(N__20002));
    LocalMux I__4203 (
            .O(N__20005),
            .I(ScreenBuffer_0_9Z0Z_0));
    Odrv4 I__4202 (
            .O(N__20002),
            .I(ScreenBuffer_0_9Z0Z_0));
    CascadeMux I__4201 (
            .O(N__19997),
            .I(N__19994));
    InMux I__4200 (
            .O(N__19994),
            .I(N__19990));
    InMux I__4199 (
            .O(N__19993),
            .I(N__19987));
    LocalMux I__4198 (
            .O(N__19990),
            .I(N__19984));
    LocalMux I__4197 (
            .O(N__19987),
            .I(N__19957));
    Glb2LocalMux I__4196 (
            .O(N__19984),
            .I(N__19892));
    ClkMux I__4195 (
            .O(N__19983),
            .I(N__19892));
    ClkMux I__4194 (
            .O(N__19982),
            .I(N__19892));
    ClkMux I__4193 (
            .O(N__19981),
            .I(N__19892));
    ClkMux I__4192 (
            .O(N__19980),
            .I(N__19892));
    ClkMux I__4191 (
            .O(N__19979),
            .I(N__19892));
    ClkMux I__4190 (
            .O(N__19978),
            .I(N__19892));
    ClkMux I__4189 (
            .O(N__19977),
            .I(N__19892));
    ClkMux I__4188 (
            .O(N__19976),
            .I(N__19892));
    ClkMux I__4187 (
            .O(N__19975),
            .I(N__19892));
    ClkMux I__4186 (
            .O(N__19974),
            .I(N__19892));
    ClkMux I__4185 (
            .O(N__19973),
            .I(N__19892));
    ClkMux I__4184 (
            .O(N__19972),
            .I(N__19892));
    ClkMux I__4183 (
            .O(N__19971),
            .I(N__19892));
    ClkMux I__4182 (
            .O(N__19970),
            .I(N__19892));
    ClkMux I__4181 (
            .O(N__19969),
            .I(N__19892));
    ClkMux I__4180 (
            .O(N__19968),
            .I(N__19892));
    ClkMux I__4179 (
            .O(N__19967),
            .I(N__19892));
    ClkMux I__4178 (
            .O(N__19966),
            .I(N__19892));
    ClkMux I__4177 (
            .O(N__19965),
            .I(N__19892));
    ClkMux I__4176 (
            .O(N__19964),
            .I(N__19892));
    ClkMux I__4175 (
            .O(N__19963),
            .I(N__19892));
    ClkMux I__4174 (
            .O(N__19962),
            .I(N__19892));
    ClkMux I__4173 (
            .O(N__19961),
            .I(N__19892));
    ClkMux I__4172 (
            .O(N__19960),
            .I(N__19892));
    Glb2LocalMux I__4171 (
            .O(N__19957),
            .I(N__19892));
    ClkMux I__4170 (
            .O(N__19956),
            .I(N__19892));
    ClkMux I__4169 (
            .O(N__19955),
            .I(N__19892));
    ClkMux I__4168 (
            .O(N__19954),
            .I(N__19892));
    ClkMux I__4167 (
            .O(N__19953),
            .I(N__19892));
    GlobalMux I__4166 (
            .O(N__19892),
            .I(N__19889));
    gio2CtrlBuf I__4165 (
            .O(N__19889),
            .I(Clock12MHz_c_g));
    InMux I__4164 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__4163 (
            .O(N__19883),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4));
    InMux I__4162 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__4161 (
            .O(N__19877),
            .I(N__19874));
    Odrv4 I__4160 (
            .O(N__19874),
            .I(column_1_if_generate_plus_mult1_un47_sum0_4));
    InMux I__4159 (
            .O(N__19871),
            .I(N__19868));
    LocalMux I__4158 (
            .O(N__19868),
            .I(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx));
    InMux I__4157 (
            .O(N__19865),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_1));
    InMux I__4156 (
            .O(N__19862),
            .I(N__19859));
    LocalMux I__4155 (
            .O(N__19859),
            .I(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx));
    CascadeMux I__4154 (
            .O(N__19856),
            .I(N__19853));
    InMux I__4153 (
            .O(N__19853),
            .I(N__19850));
    LocalMux I__4152 (
            .O(N__19850),
            .I(if_generate_plus_mult1_un47_sum_0_cry_3_ma));
    InMux I__4151 (
            .O(N__19847),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_2));
    InMux I__4150 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__4149 (
            .O(N__19841),
            .I(N_1184_0_i));
    InMux I__4148 (
            .O(N__19838),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_3));
    InMux I__4147 (
            .O(N__19835),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_4));
    CascadeMux I__4146 (
            .O(N__19832),
            .I(N__19829));
    InMux I__4145 (
            .O(N__19829),
            .I(N__19826));
    LocalMux I__4144 (
            .O(N__19826),
            .I(un5_visiblex_i_25));
    CascadeMux I__4143 (
            .O(N__19823),
            .I(N_2110_i_cascade_));
    InMux I__4142 (
            .O(N__19820),
            .I(N__19814));
    InMux I__4141 (
            .O(N__19819),
            .I(N__19814));
    LocalMux I__4140 (
            .O(N__19814),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    CascadeMux I__4139 (
            .O(N__19811),
            .I(un115_pixel_6_bm_2_cascade_));
    InMux I__4138 (
            .O(N__19808),
            .I(N__19805));
    LocalMux I__4137 (
            .O(N__19805),
            .I(N__19802));
    Odrv12 I__4136 (
            .O(N__19802),
            .I(N_1330));
    InMux I__4135 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__4134 (
            .O(N__19796),
            .I(un115_pixel_6_am_2));
    InMux I__4133 (
            .O(N__19793),
            .I(N__19789));
    CascadeMux I__4132 (
            .O(N__19792),
            .I(N__19786));
    LocalMux I__4131 (
            .O(N__19789),
            .I(N__19783));
    InMux I__4130 (
            .O(N__19786),
            .I(N__19780));
    Odrv4 I__4129 (
            .O(N__19783),
            .I(un5_visiblex_i_24));
    LocalMux I__4128 (
            .O(N__19780),
            .I(un5_visiblex_i_24));
    CascadeMux I__4127 (
            .O(N__19775),
            .I(N__19772));
    InMux I__4126 (
            .O(N__19772),
            .I(N__19769));
    LocalMux I__4125 (
            .O(N__19769),
            .I(N__19766));
    Span4Mux_h I__4124 (
            .O(N__19766),
            .I(N__19763));
    Odrv4 I__4123 (
            .O(N__19763),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0));
    InMux I__4122 (
            .O(N__19760),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__4121 (
            .O(N__19757),
            .I(N__19753));
    InMux I__4120 (
            .O(N__19756),
            .I(N__19748));
    InMux I__4119 (
            .O(N__19753),
            .I(N__19748));
    LocalMux I__4118 (
            .O(N__19748),
            .I(N__19745));
    Span4Mux_h I__4117 (
            .O(N__19745),
            .I(N__19742));
    Odrv4 I__4116 (
            .O(N__19742),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0));
    InMux I__4115 (
            .O(N__19739),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__4114 (
            .O(N__19736),
            .I(N__19733));
    LocalMux I__4113 (
            .O(N__19733),
            .I(N__19730));
    Span4Mux_h I__4112 (
            .O(N__19730),
            .I(N__19727));
    Odrv4 I__4111 (
            .O(N__19727),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__4110 (
            .O(N__19724),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__4109 (
            .O(N__19721),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__4108 (
            .O(N__19718),
            .I(N__19712));
    InMux I__4107 (
            .O(N__19717),
            .I(N__19709));
    InMux I__4106 (
            .O(N__19716),
            .I(N__19706));
    InMux I__4105 (
            .O(N__19715),
            .I(N__19703));
    LocalMux I__4104 (
            .O(N__19712),
            .I(N__19698));
    LocalMux I__4103 (
            .O(N__19709),
            .I(N__19698));
    LocalMux I__4102 (
            .O(N__19706),
            .I(N__19691));
    LocalMux I__4101 (
            .O(N__19703),
            .I(N__19691));
    Span4Mux_v I__4100 (
            .O(N__19698),
            .I(N__19691));
    Odrv4 I__4099 (
            .O(N__19691),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0));
    InMux I__4098 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__4097 (
            .O(N__19685),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__4096 (
            .O(N__19682),
            .I(N__19678));
    InMux I__4095 (
            .O(N__19681),
            .I(N__19670));
    InMux I__4094 (
            .O(N__19678),
            .I(N__19670));
    InMux I__4093 (
            .O(N__19677),
            .I(N__19670));
    LocalMux I__4092 (
            .O(N__19670),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12));
    CascadeMux I__4091 (
            .O(N__19667),
            .I(m14_cascade_));
    InMux I__4090 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__4089 (
            .O(N__19661),
            .I(beamY_RNI7RM4IFZ0Z_0));
    InMux I__4088 (
            .O(N__19658),
            .I(N__19655));
    LocalMux I__4087 (
            .O(N__19655),
            .I(un113_pixel_3_0_11__g1_1_0));
    InMux I__4086 (
            .O(N__19652),
            .I(N__19649));
    LocalMux I__4085 (
            .O(N__19649),
            .I(beamY_RNIPQEDM42Z0Z_0));
    InMux I__4084 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__4083 (
            .O(N__19643),
            .I(N_1293));
    CascadeMux I__4082 (
            .O(N__19640),
            .I(N_1306_cascade_));
    InMux I__4081 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__4080 (
            .O(N__19634),
            .I(N_1327_0));
    CascadeMux I__4079 (
            .O(N__19631),
            .I(m11_cascade_));
    InMux I__4078 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__4077 (
            .O(N__19625),
            .I(un113_pixel_4_0_15__N_17));
    InMux I__4076 (
            .O(N__19622),
            .I(N__19619));
    LocalMux I__4075 (
            .O(N__19619),
            .I(un115_pixel_4_am_7));
    CascadeMux I__4074 (
            .O(N__19616),
            .I(N_1287_cascade_));
    CascadeMux I__4073 (
            .O(N__19613),
            .I(currentchar_1_0_cascade_));
    InMux I__4072 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__4071 (
            .O(N__19607),
            .I(un115_pixel_4_bm_7));
    InMux I__4070 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__4069 (
            .O(N__19601),
            .I(N__19595));
    InMux I__4068 (
            .O(N__19600),
            .I(N__19590));
    InMux I__4067 (
            .O(N__19599),
            .I(N__19590));
    InMux I__4066 (
            .O(N__19598),
            .I(N__19587));
    Odrv4 I__4065 (
            .O(N__19595),
            .I(ScreenBuffer_0_7_RNII0GVLQZ0Z_0));
    LocalMux I__4064 (
            .O(N__19590),
            .I(ScreenBuffer_0_7_RNII0GVLQZ0Z_0));
    LocalMux I__4063 (
            .O(N__19587),
            .I(ScreenBuffer_0_7_RNII0GVLQZ0Z_0));
    CascadeMux I__4062 (
            .O(N__19580),
            .I(un113_pixel_1_0_3__N_10_mux_cascade_));
    CascadeMux I__4061 (
            .O(N__19577),
            .I(N_1285_0_0_0_cascade_));
    InMux I__4060 (
            .O(N__19574),
            .I(N__19571));
    LocalMux I__4059 (
            .O(N__19571),
            .I(N__19568));
    Span4Mux_v I__4058 (
            .O(N__19568),
            .I(N__19565));
    Span4Mux_h I__4057 (
            .O(N__19565),
            .I(N__19562));
    Odrv4 I__4056 (
            .O(N__19562),
            .I(un113_pixel_3_0_11__g1_0_0_0));
    InMux I__4055 (
            .O(N__19559),
            .I(N__19556));
    LocalMux I__4054 (
            .O(N__19556),
            .I(m14));
    CascadeMux I__4053 (
            .O(N__19553),
            .I(ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_));
    CascadeMux I__4052 (
            .O(N__19550),
            .I(currentchar_m7_0_cascade_));
    CascadeMux I__4051 (
            .O(N__19547),
            .I(N__19543));
    InMux I__4050 (
            .O(N__19546),
            .I(N__19540));
    InMux I__4049 (
            .O(N__19543),
            .I(N__19537));
    LocalMux I__4048 (
            .O(N__19540),
            .I(N__19534));
    LocalMux I__4047 (
            .O(N__19537),
            .I(N__19529));
    Span4Mux_v I__4046 (
            .O(N__19534),
            .I(N__19529));
    Odrv4 I__4045 (
            .O(N__19529),
            .I(ScreenBuffer_0_7Z0Z_0));
    InMux I__4044 (
            .O(N__19526),
            .I(N__19522));
    InMux I__4043 (
            .O(N__19525),
            .I(N__19519));
    LocalMux I__4042 (
            .O(N__19522),
            .I(N__19516));
    LocalMux I__4041 (
            .O(N__19519),
            .I(ScreenBuffer_0_5Z0Z_0));
    Odrv4 I__4040 (
            .O(N__19516),
            .I(ScreenBuffer_0_5Z0Z_0));
    InMux I__4039 (
            .O(N__19511),
            .I(N__19507));
    InMux I__4038 (
            .O(N__19510),
            .I(N__19504));
    LocalMux I__4037 (
            .O(N__19507),
            .I(N__19500));
    LocalMux I__4036 (
            .O(N__19504),
            .I(N__19497));
    InMux I__4035 (
            .O(N__19503),
            .I(N__19494));
    Odrv4 I__4034 (
            .O(N__19500),
            .I(un113_pixel_3_0_11__currentchar_N_13));
    Odrv4 I__4033 (
            .O(N__19497),
            .I(un113_pixel_3_0_11__currentchar_N_13));
    LocalMux I__4032 (
            .O(N__19494),
            .I(un113_pixel_3_0_11__currentchar_N_13));
    InMux I__4031 (
            .O(N__19487),
            .I(N__19484));
    LocalMux I__4030 (
            .O(N__19484),
            .I(un112_pixel_1_2_x1));
    CascadeMux I__4029 (
            .O(N__19481),
            .I(un112_pixel_2_8_cascade_));
    InMux I__4028 (
            .O(N__19478),
            .I(N__19475));
    LocalMux I__4027 (
            .O(N__19475),
            .I(N__19472));
    Odrv4 I__4026 (
            .O(N__19472),
            .I(ScreenBuffer_1_2Z0Z_3));
    CascadeMux I__4025 (
            .O(N__19469),
            .I(un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_));
    CascadeMux I__4024 (
            .O(N__19466),
            .I(un113_pixel_3_0_11__currentchar_N_13_cascade_));
    InMux I__4023 (
            .O(N__19463),
            .I(N__19459));
    InMux I__4022 (
            .O(N__19462),
            .I(N__19456));
    LocalMux I__4021 (
            .O(N__19459),
            .I(N__19451));
    LocalMux I__4020 (
            .O(N__19456),
            .I(N__19451));
    Span12Mux_s11_v I__4019 (
            .O(N__19451),
            .I(N__19446));
    InMux I__4018 (
            .O(N__19450),
            .I(N__19443));
    InMux I__4017 (
            .O(N__19449),
            .I(N__19440));
    Odrv12 I__4016 (
            .O(N__19446),
            .I(voltage_3Z0Z_3));
    LocalMux I__4015 (
            .O(N__19443),
            .I(voltage_3Z0Z_3));
    LocalMux I__4014 (
            .O(N__19440),
            .I(voltage_3Z0Z_3));
    InMux I__4013 (
            .O(N__19433),
            .I(N__19429));
    InMux I__4012 (
            .O(N__19432),
            .I(N__19426));
    LocalMux I__4011 (
            .O(N__19429),
            .I(N__19423));
    LocalMux I__4010 (
            .O(N__19426),
            .I(N__19420));
    Span4Mux_v I__4009 (
            .O(N__19423),
            .I(N__19413));
    Span4Mux_v I__4008 (
            .O(N__19420),
            .I(N__19413));
    InMux I__4007 (
            .O(N__19419),
            .I(N__19407));
    InMux I__4006 (
            .O(N__19418),
            .I(N__19407));
    Span4Mux_h I__4005 (
            .O(N__19413),
            .I(N__19404));
    InMux I__4004 (
            .O(N__19412),
            .I(N__19401));
    LocalMux I__4003 (
            .O(N__19407),
            .I(N__19398));
    Odrv4 I__4002 (
            .O(N__19404),
            .I(voltage_0Z0Z_3));
    LocalMux I__4001 (
            .O(N__19401),
            .I(voltage_0Z0Z_3));
    Odrv4 I__4000 (
            .O(N__19398),
            .I(voltage_0Z0Z_3));
    InMux I__3999 (
            .O(N__19391),
            .I(N__19388));
    LocalMux I__3998 (
            .O(N__19388),
            .I(ScreenBuffer_1_0Z0Z_3));
    InMux I__3997 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__3996 (
            .O(N__19382),
            .I(un113_pixel_4_0_15__g0_1Z0Z_0));
    InMux I__3995 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__3994 (
            .O(N__19376),
            .I(un113_pixel_4_0_15__g0_3_0));
    InMux I__3993 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__3992 (
            .O(N__19370),
            .I(N__19365));
    InMux I__3991 (
            .O(N__19369),
            .I(N__19362));
    InMux I__3990 (
            .O(N__19368),
            .I(N__19359));
    Span4Mux_v I__3989 (
            .O(N__19365),
            .I(N__19356));
    LocalMux I__3988 (
            .O(N__19362),
            .I(N__19353));
    LocalMux I__3987 (
            .O(N__19359),
            .I(N__19349));
    Span4Mux_h I__3986 (
            .O(N__19356),
            .I(N__19344));
    Span4Mux_s3_h I__3985 (
            .O(N__19353),
            .I(N__19344));
    InMux I__3984 (
            .O(N__19352),
            .I(N__19341));
    Odrv12 I__3983 (
            .O(N__19349),
            .I(voltage_3Z0Z_1));
    Odrv4 I__3982 (
            .O(N__19344),
            .I(voltage_3Z0Z_1));
    LocalMux I__3981 (
            .O(N__19341),
            .I(voltage_3Z0Z_1));
    InMux I__3980 (
            .O(N__19334),
            .I(N__19323));
    InMux I__3979 (
            .O(N__19333),
            .I(N__19315));
    InMux I__3978 (
            .O(N__19332),
            .I(N__19310));
    InMux I__3977 (
            .O(N__19331),
            .I(N__19310));
    InMux I__3976 (
            .O(N__19330),
            .I(N__19296));
    InMux I__3975 (
            .O(N__19329),
            .I(N__19293));
    CascadeMux I__3974 (
            .O(N__19328),
            .I(N__19285));
    CascadeMux I__3973 (
            .O(N__19327),
            .I(N__19281));
    InMux I__3972 (
            .O(N__19326),
            .I(N__19277));
    LocalMux I__3971 (
            .O(N__19323),
            .I(N__19274));
    InMux I__3970 (
            .O(N__19322),
            .I(N__19265));
    InMux I__3969 (
            .O(N__19321),
            .I(N__19265));
    InMux I__3968 (
            .O(N__19320),
            .I(N__19265));
    InMux I__3967 (
            .O(N__19319),
            .I(N__19265));
    InMux I__3966 (
            .O(N__19318),
            .I(N__19262));
    LocalMux I__3965 (
            .O(N__19315),
            .I(N__19257));
    LocalMux I__3964 (
            .O(N__19310),
            .I(N__19257));
    InMux I__3963 (
            .O(N__19309),
            .I(N__19252));
    InMux I__3962 (
            .O(N__19308),
            .I(N__19252));
    InMux I__3961 (
            .O(N__19307),
            .I(N__19243));
    InMux I__3960 (
            .O(N__19306),
            .I(N__19243));
    InMux I__3959 (
            .O(N__19305),
            .I(N__19234));
    InMux I__3958 (
            .O(N__19304),
            .I(N__19234));
    InMux I__3957 (
            .O(N__19303),
            .I(N__19234));
    InMux I__3956 (
            .O(N__19302),
            .I(N__19234));
    InMux I__3955 (
            .O(N__19301),
            .I(N__19229));
    InMux I__3954 (
            .O(N__19300),
            .I(N__19229));
    InMux I__3953 (
            .O(N__19299),
            .I(N__19226));
    LocalMux I__3952 (
            .O(N__19296),
            .I(N__19221));
    LocalMux I__3951 (
            .O(N__19293),
            .I(N__19221));
    InMux I__3950 (
            .O(N__19292),
            .I(N__19218));
    InMux I__3949 (
            .O(N__19291),
            .I(N__19213));
    InMux I__3948 (
            .O(N__19290),
            .I(N__19213));
    InMux I__3947 (
            .O(N__19289),
            .I(N__19210));
    InMux I__3946 (
            .O(N__19288),
            .I(N__19203));
    InMux I__3945 (
            .O(N__19285),
            .I(N__19203));
    InMux I__3944 (
            .O(N__19284),
            .I(N__19203));
    InMux I__3943 (
            .O(N__19281),
            .I(N__19198));
    InMux I__3942 (
            .O(N__19280),
            .I(N__19198));
    LocalMux I__3941 (
            .O(N__19277),
            .I(N__19187));
    Span4Mux_h I__3940 (
            .O(N__19274),
            .I(N__19187));
    LocalMux I__3939 (
            .O(N__19265),
            .I(N__19187));
    LocalMux I__3938 (
            .O(N__19262),
            .I(N__19187));
    Span4Mux_s3_v I__3937 (
            .O(N__19257),
            .I(N__19187));
    LocalMux I__3936 (
            .O(N__19252),
            .I(N__19184));
    InMux I__3935 (
            .O(N__19251),
            .I(N__19167));
    InMux I__3934 (
            .O(N__19250),
            .I(N__19167));
    InMux I__3933 (
            .O(N__19249),
            .I(N__19167));
    InMux I__3932 (
            .O(N__19248),
            .I(N__19167));
    LocalMux I__3931 (
            .O(N__19243),
            .I(N__19146));
    LocalMux I__3930 (
            .O(N__19234),
            .I(N__19146));
    LocalMux I__3929 (
            .O(N__19229),
            .I(N__19146));
    LocalMux I__3928 (
            .O(N__19226),
            .I(N__19146));
    Span4Mux_v I__3927 (
            .O(N__19221),
            .I(N__19146));
    LocalMux I__3926 (
            .O(N__19218),
            .I(N__19146));
    LocalMux I__3925 (
            .O(N__19213),
            .I(N__19146));
    LocalMux I__3924 (
            .O(N__19210),
            .I(N__19146));
    LocalMux I__3923 (
            .O(N__19203),
            .I(N__19146));
    LocalMux I__3922 (
            .O(N__19198),
            .I(N__19146));
    Span4Mux_v I__3921 (
            .O(N__19187),
            .I(N__19143));
    Span4Mux_v I__3920 (
            .O(N__19184),
            .I(N__19140));
    InMux I__3919 (
            .O(N__19183),
            .I(N__19135));
    InMux I__3918 (
            .O(N__19182),
            .I(N__19135));
    InMux I__3917 (
            .O(N__19181),
            .I(N__19132));
    InMux I__3916 (
            .O(N__19180),
            .I(N__19127));
    InMux I__3915 (
            .O(N__19179),
            .I(N__19127));
    InMux I__3914 (
            .O(N__19178),
            .I(N__19124));
    InMux I__3913 (
            .O(N__19177),
            .I(N__19121));
    InMux I__3912 (
            .O(N__19176),
            .I(N__19118));
    LocalMux I__3911 (
            .O(N__19167),
            .I(N__19115));
    Span4Mux_v I__3910 (
            .O(N__19146),
            .I(N__19107));
    Span4Mux_v I__3909 (
            .O(N__19143),
            .I(N__19102));
    Span4Mux_v I__3908 (
            .O(N__19140),
            .I(N__19102));
    LocalMux I__3907 (
            .O(N__19135),
            .I(N__19093));
    LocalMux I__3906 (
            .O(N__19132),
            .I(N__19093));
    LocalMux I__3905 (
            .O(N__19127),
            .I(N__19093));
    LocalMux I__3904 (
            .O(N__19124),
            .I(N__19093));
    LocalMux I__3903 (
            .O(N__19121),
            .I(N__19086));
    LocalMux I__3902 (
            .O(N__19118),
            .I(N__19086));
    Span4Mux_h I__3901 (
            .O(N__19115),
            .I(N__19086));
    InMux I__3900 (
            .O(N__19114),
            .I(N__19081));
    InMux I__3899 (
            .O(N__19113),
            .I(N__19081));
    InMux I__3898 (
            .O(N__19112),
            .I(N__19074));
    InMux I__3897 (
            .O(N__19111),
            .I(N__19074));
    InMux I__3896 (
            .O(N__19110),
            .I(N__19074));
    Span4Mux_h I__3895 (
            .O(N__19107),
            .I(N__19071));
    Sp12to4 I__3894 (
            .O(N__19102),
            .I(N__19066));
    Span12Mux_s11_v I__3893 (
            .O(N__19093),
            .I(N__19066));
    Span4Mux_v I__3892 (
            .O(N__19086),
            .I(N__19063));
    LocalMux I__3891 (
            .O(N__19081),
            .I(slaveselectZ0));
    LocalMux I__3890 (
            .O(N__19074),
            .I(slaveselectZ0));
    Odrv4 I__3889 (
            .O(N__19071),
            .I(slaveselectZ0));
    Odrv12 I__3888 (
            .O(N__19066),
            .I(slaveselectZ0));
    Odrv4 I__3887 (
            .O(N__19063),
            .I(slaveselectZ0));
    InMux I__3886 (
            .O(N__19052),
            .I(N__19048));
    InMux I__3885 (
            .O(N__19051),
            .I(N__19043));
    LocalMux I__3884 (
            .O(N__19048),
            .I(N__19040));
    InMux I__3883 (
            .O(N__19047),
            .I(N__19037));
    InMux I__3882 (
            .O(N__19046),
            .I(N__19034));
    LocalMux I__3881 (
            .O(N__19043),
            .I(N__19031));
    Span4Mux_v I__3880 (
            .O(N__19040),
            .I(N__19027));
    LocalMux I__3879 (
            .O(N__19037),
            .I(N__19024));
    LocalMux I__3878 (
            .O(N__19034),
            .I(N__19021));
    Span4Mux_v I__3877 (
            .O(N__19031),
            .I(N__19018));
    InMux I__3876 (
            .O(N__19030),
            .I(N__19015));
    Span4Mux_h I__3875 (
            .O(N__19027),
            .I(N__19010));
    Span4Mux_v I__3874 (
            .O(N__19024),
            .I(N__19010));
    Span4Mux_v I__3873 (
            .O(N__19021),
            .I(N__19005));
    Span4Mux_h I__3872 (
            .O(N__19018),
            .I(N__19005));
    LocalMux I__3871 (
            .O(N__19015),
            .I(voltage_0Z0Z_1));
    Odrv4 I__3870 (
            .O(N__19010),
            .I(voltage_0Z0Z_1));
    Odrv4 I__3869 (
            .O(N__19005),
            .I(voltage_0Z0Z_1));
    CEMux I__3868 (
            .O(N__18998),
            .I(N__18994));
    CEMux I__3867 (
            .O(N__18997),
            .I(N__18991));
    LocalMux I__3866 (
            .O(N__18994),
            .I(N__18988));
    LocalMux I__3865 (
            .O(N__18991),
            .I(N__18985));
    Span4Mux_v I__3864 (
            .O(N__18988),
            .I(N__18982));
    Span4Mux_h I__3863 (
            .O(N__18985),
            .I(N__18979));
    Odrv4 I__3862 (
            .O(N__18982),
            .I(un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0));
    Odrv4 I__3861 (
            .O(N__18979),
            .I(un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0));
    InMux I__3860 (
            .O(N__18974),
            .I(N__18970));
    InMux I__3859 (
            .O(N__18973),
            .I(N__18967));
    LocalMux I__3858 (
            .O(N__18970),
            .I(N__18964));
    LocalMux I__3857 (
            .O(N__18967),
            .I(ScreenBuffer_0_12Z0Z_0));
    Odrv4 I__3856 (
            .O(N__18964),
            .I(ScreenBuffer_0_12Z0Z_0));
    InMux I__3855 (
            .O(N__18959),
            .I(N__18955));
    InMux I__3854 (
            .O(N__18958),
            .I(N__18952));
    LocalMux I__3853 (
            .O(N__18955),
            .I(N__18949));
    LocalMux I__3852 (
            .O(N__18952),
            .I(ScreenBuffer_0_4Z0Z_0));
    Odrv12 I__3851 (
            .O(N__18949),
            .I(ScreenBuffer_0_4Z0Z_0));
    CascadeMux I__3850 (
            .O(N__18944),
            .I(ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_));
    InMux I__3849 (
            .O(N__18941),
            .I(N__18937));
    CascadeMux I__3848 (
            .O(N__18940),
            .I(N__18934));
    LocalMux I__3847 (
            .O(N__18937),
            .I(N__18931));
    InMux I__3846 (
            .O(N__18934),
            .I(N__18928));
    Span4Mux_h I__3845 (
            .O(N__18931),
            .I(N__18925));
    LocalMux I__3844 (
            .O(N__18928),
            .I(ScreenBuffer_0_6Z0Z_0));
    Odrv4 I__3843 (
            .O(N__18925),
            .I(ScreenBuffer_0_6Z0Z_0));
    CascadeMux I__3842 (
            .O(N__18920),
            .I(beamY_RNIOEPPEK1Z0Z_0_cascade_));
    InMux I__3841 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__3840 (
            .O(N__18914),
            .I(un112_pixel_1_2));
    CascadeMux I__3839 (
            .O(N__18911),
            .I(N_3461_0_cascade_));
    CascadeMux I__3838 (
            .O(N__18908),
            .I(N_4568_0_cascade_));
    InMux I__3837 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__3836 (
            .O(N__18902),
            .I(N_1305_0));
    InMux I__3835 (
            .O(N__18899),
            .I(N__18896));
    LocalMux I__3834 (
            .O(N__18896),
            .I(un113_pixel_4_0_15__g0_0Z0Z_2));
    InMux I__3833 (
            .O(N__18893),
            .I(N__18890));
    LocalMux I__3832 (
            .O(N__18890),
            .I(N__18887));
    Span4Mux_v I__3831 (
            .O(N__18887),
            .I(N__18884));
    Odrv4 I__3830 (
            .O(N__18884),
            .I(Pixel_3_sqmuxa_0));
    InMux I__3829 (
            .O(N__18881),
            .I(N__18878));
    LocalMux I__3828 (
            .O(N__18878),
            .I(g0_1_1));
    CascadeMux I__3827 (
            .O(N__18875),
            .I(N_1_0_cascade_));
    InMux I__3826 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__3825 (
            .O(N__18869),
            .I(N__18866));
    Odrv12 I__3824 (
            .O(N__18866),
            .I(ScreenBuffer_1_3Z0Z_3));
    InMux I__3823 (
            .O(N__18863),
            .I(N__18860));
    LocalMux I__3822 (
            .O(N__18860),
            .I(N__18857));
    Span4Mux_v I__3821 (
            .O(N__18857),
            .I(N__18854));
    Odrv4 I__3820 (
            .O(N__18854),
            .I(ScreenBuffer_1_1Z0Z_3));
    CascadeMux I__3819 (
            .O(N__18851),
            .I(N__18848));
    InMux I__3818 (
            .O(N__18848),
            .I(N__18845));
    LocalMux I__3817 (
            .O(N__18845),
            .I(column_1_if_generate_plus_mult1_un61_sum_iZ0));
    CascadeMux I__3816 (
            .O(N__18842),
            .I(N__18839));
    InMux I__3815 (
            .O(N__18839),
            .I(N__18835));
    InMux I__3814 (
            .O(N__18838),
            .I(N__18832));
    LocalMux I__3813 (
            .O(N__18835),
            .I(chary_24));
    LocalMux I__3812 (
            .O(N__18832),
            .I(chary_24));
    CascadeMux I__3811 (
            .O(N__18827),
            .I(N__18824));
    InMux I__3810 (
            .O(N__18824),
            .I(N__18821));
    LocalMux I__3809 (
            .O(N__18821),
            .I(N__18818));
    Odrv4 I__3808 (
            .O(N__18818),
            .I(un113_pixel_4_0_15__gZ0Z2));
    InMux I__3807 (
            .O(N__18815),
            .I(N__18811));
    InMux I__3806 (
            .O(N__18814),
            .I(N__18808));
    LocalMux I__3805 (
            .O(N__18811),
            .I(font_un3_pixel_30));
    LocalMux I__3804 (
            .O(N__18808),
            .I(font_un3_pixel_30));
    InMux I__3803 (
            .O(N__18803),
            .I(N__18800));
    LocalMux I__3802 (
            .O(N__18800),
            .I(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1));
    CascadeMux I__3801 (
            .O(N__18797),
            .I(font_un57_pixel_cascade_));
    InMux I__3800 (
            .O(N__18794),
            .I(N__18791));
    LocalMux I__3799 (
            .O(N__18791),
            .I(currentchar_1_5));
    InMux I__3798 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__3797 (
            .O(N__18785),
            .I(N__18782));
    Odrv4 I__3796 (
            .O(N__18782),
            .I(font_un67_pixel_ac0_5));
    InMux I__3795 (
            .O(N__18779),
            .I(N__18776));
    LocalMux I__3794 (
            .O(N__18776),
            .I(font_un64_pixel_ac0_5));
    CascadeMux I__3793 (
            .O(N__18773),
            .I(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_));
    InMux I__3792 (
            .O(N__18770),
            .I(N__18767));
    LocalMux I__3791 (
            .O(N__18767),
            .I(N__18764));
    Span4Mux_h I__3790 (
            .O(N__18764),
            .I(N__18761));
    Odrv4 I__3789 (
            .O(N__18761),
            .I(N_12));
    CascadeMux I__3788 (
            .O(N__18758),
            .I(N__18755));
    InMux I__3787 (
            .O(N__18755),
            .I(N__18752));
    LocalMux I__3786 (
            .O(N__18752),
            .I(N__18749));
    Odrv4 I__3785 (
            .O(N__18749),
            .I(un113_pixel_4_0_15__g0_iZ0Z_2));
    CascadeMux I__3784 (
            .O(N__18746),
            .I(un113_pixel_4_0_15__g0_iZ0Z_5_cascade_));
    CascadeMux I__3783 (
            .O(N__18743),
            .I(N__18737));
    CascadeMux I__3782 (
            .O(N__18742),
            .I(N__18733));
    InMux I__3781 (
            .O(N__18741),
            .I(N__18726));
    InMux I__3780 (
            .O(N__18740),
            .I(N__18726));
    InMux I__3779 (
            .O(N__18737),
            .I(N__18726));
    CascadeMux I__3778 (
            .O(N__18736),
            .I(N__18721));
    InMux I__3777 (
            .O(N__18733),
            .I(N__18717));
    LocalMux I__3776 (
            .O(N__18726),
            .I(N__18714));
    InMux I__3775 (
            .O(N__18725),
            .I(N__18711));
    InMux I__3774 (
            .O(N__18724),
            .I(N__18708));
    InMux I__3773 (
            .O(N__18721),
            .I(N__18705));
    CascadeMux I__3772 (
            .O(N__18720),
            .I(N__18701));
    LocalMux I__3771 (
            .O(N__18717),
            .I(N__18695));
    Span4Mux_h I__3770 (
            .O(N__18714),
            .I(N__18692));
    LocalMux I__3769 (
            .O(N__18711),
            .I(N__18687));
    LocalMux I__3768 (
            .O(N__18708),
            .I(N__18687));
    LocalMux I__3767 (
            .O(N__18705),
            .I(N__18684));
    InMux I__3766 (
            .O(N__18704),
            .I(N__18679));
    InMux I__3765 (
            .O(N__18701),
            .I(N__18679));
    InMux I__3764 (
            .O(N__18700),
            .I(N__18676));
    InMux I__3763 (
            .O(N__18699),
            .I(N__18673));
    InMux I__3762 (
            .O(N__18698),
            .I(N__18670));
    Span4Mux_s2_v I__3761 (
            .O(N__18695),
            .I(N__18667));
    Span4Mux_v I__3760 (
            .O(N__18692),
            .I(N__18664));
    Span4Mux_v I__3759 (
            .O(N__18687),
            .I(N__18661));
    Span4Mux_v I__3758 (
            .O(N__18684),
            .I(N__18656));
    LocalMux I__3757 (
            .O(N__18679),
            .I(N__18656));
    LocalMux I__3756 (
            .O(N__18676),
            .I(N__18653));
    LocalMux I__3755 (
            .O(N__18673),
            .I(beamXZ0Z_0));
    LocalMux I__3754 (
            .O(N__18670),
            .I(beamXZ0Z_0));
    Odrv4 I__3753 (
            .O(N__18667),
            .I(beamXZ0Z_0));
    Odrv4 I__3752 (
            .O(N__18664),
            .I(beamXZ0Z_0));
    Odrv4 I__3751 (
            .O(N__18661),
            .I(beamXZ0Z_0));
    Odrv4 I__3750 (
            .O(N__18656),
            .I(beamXZ0Z_0));
    Odrv4 I__3749 (
            .O(N__18653),
            .I(beamXZ0Z_0));
    InMux I__3748 (
            .O(N__18638),
            .I(N__18632));
    InMux I__3747 (
            .O(N__18637),
            .I(N__18632));
    LocalMux I__3746 (
            .O(N__18632),
            .I(un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6));
    InMux I__3745 (
            .O(N__18629),
            .I(N__18623));
    InMux I__3744 (
            .O(N__18628),
            .I(N__18623));
    LocalMux I__3743 (
            .O(N__18623),
            .I(charx_if_generate_plus_mult1_un68_sum_i_5));
    InMux I__3742 (
            .O(N__18620),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__3741 (
            .O(N__18617),
            .I(N__18602));
    InMux I__3740 (
            .O(N__18616),
            .I(N__18602));
    InMux I__3739 (
            .O(N__18615),
            .I(N__18602));
    InMux I__3738 (
            .O(N__18614),
            .I(N__18602));
    InMux I__3737 (
            .O(N__18613),
            .I(N__18602));
    LocalMux I__3736 (
            .O(N__18602),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1));
    CascadeMux I__3735 (
            .O(N__18599),
            .I(N__18596));
    InMux I__3734 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__3733 (
            .O(N__18593),
            .I(charx_if_generate_plus_mult1_un68_sum_i));
    InMux I__3732 (
            .O(N__18590),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__3731 (
            .O(N__18587),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__3730 (
            .O(N__18584),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__3729 (
            .O(N__18581),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__3728 (
            .O(N__18578),
            .I(N__18572));
    InMux I__3727 (
            .O(N__18577),
            .I(N__18572));
    LocalMux I__3726 (
            .O(N__18572),
            .I(N__18569));
    Span4Mux_v I__3725 (
            .O(N__18569),
            .I(N__18565));
    InMux I__3724 (
            .O(N__18568),
            .I(N__18562));
    Span4Mux_h I__3723 (
            .O(N__18565),
            .I(N__18559));
    LocalMux I__3722 (
            .O(N__18562),
            .I(N__18556));
    Span4Mux_v I__3721 (
            .O(N__18559),
            .I(N__18551));
    Span4Mux_h I__3720 (
            .O(N__18556),
            .I(N__18551));
    Odrv4 I__3719 (
            .O(N__18551),
            .I(un1_counter_1_0));
    SRMux I__3718 (
            .O(N__18548),
            .I(N__18524));
    SRMux I__3717 (
            .O(N__18547),
            .I(N__18524));
    SRMux I__3716 (
            .O(N__18546),
            .I(N__18524));
    SRMux I__3715 (
            .O(N__18545),
            .I(N__18524));
    SRMux I__3714 (
            .O(N__18544),
            .I(N__18524));
    SRMux I__3713 (
            .O(N__18543),
            .I(N__18524));
    SRMux I__3712 (
            .O(N__18542),
            .I(N__18524));
    SRMux I__3711 (
            .O(N__18541),
            .I(N__18524));
    GlobalMux I__3710 (
            .O(N__18524),
            .I(N__18521));
    gio2CtrlBuf I__3709 (
            .O(N__18521),
            .I(voltage_0_0_sqmuxa_1_g));
    InMux I__3708 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__3707 (
            .O(N__18515),
            .I(N__18512));
    Span4Mux_v I__3706 (
            .O(N__18512),
            .I(N__18509));
    Span4Mux_h I__3705 (
            .O(N__18509),
            .I(N__18506));
    Span4Mux_h I__3704 (
            .O(N__18506),
            .I(N__18500));
    InMux I__3703 (
            .O(N__18505),
            .I(N__18497));
    InMux I__3702 (
            .O(N__18504),
            .I(N__18494));
    InMux I__3701 (
            .O(N__18503),
            .I(N__18491));
    Odrv4 I__3700 (
            .O(N__18500),
            .I(voltage_3Z0Z_0));
    LocalMux I__3699 (
            .O(N__18497),
            .I(voltage_3Z0Z_0));
    LocalMux I__3698 (
            .O(N__18494),
            .I(voltage_3Z0Z_0));
    LocalMux I__3697 (
            .O(N__18491),
            .I(voltage_3Z0Z_0));
    InMux I__3696 (
            .O(N__18482),
            .I(N__18469));
    InMux I__3695 (
            .O(N__18481),
            .I(N__18469));
    InMux I__3694 (
            .O(N__18480),
            .I(N__18469));
    InMux I__3693 (
            .O(N__18479),
            .I(N__18469));
    InMux I__3692 (
            .O(N__18478),
            .I(N__18466));
    LocalMux I__3691 (
            .O(N__18469),
            .I(N__18463));
    LocalMux I__3690 (
            .O(N__18466),
            .I(N__18460));
    Span4Mux_s3_h I__3689 (
            .O(N__18463),
            .I(N__18457));
    Span4Mux_v I__3688 (
            .O(N__18460),
            .I(N__18453));
    Span4Mux_h I__3687 (
            .O(N__18457),
            .I(N__18450));
    InMux I__3686 (
            .O(N__18456),
            .I(N__18447));
    Span4Mux_h I__3685 (
            .O(N__18453),
            .I(N__18444));
    Span4Mux_v I__3684 (
            .O(N__18450),
            .I(N__18441));
    LocalMux I__3683 (
            .O(N__18447),
            .I(voltage_0Z0Z_0));
    Odrv4 I__3682 (
            .O(N__18444),
            .I(voltage_0Z0Z_0));
    Odrv4 I__3681 (
            .O(N__18441),
            .I(voltage_0Z0Z_0));
    CEMux I__3680 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__3679 (
            .O(N__18431),
            .I(N__18427));
    CEMux I__3678 (
            .O(N__18430),
            .I(N__18424));
    Span4Mux_h I__3677 (
            .O(N__18427),
            .I(N__18421));
    LocalMux I__3676 (
            .O(N__18424),
            .I(N__18418));
    Span4Mux_v I__3675 (
            .O(N__18421),
            .I(N__18415));
    Span4Mux_v I__3674 (
            .O(N__18418),
            .I(N__18412));
    Odrv4 I__3673 (
            .O(N__18415),
            .I(un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0));
    Odrv4 I__3672 (
            .O(N__18412),
            .I(un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0));
    CascadeMux I__3671 (
            .O(N__18407),
            .I(N__18403));
    CascadeMux I__3670 (
            .O(N__18406),
            .I(N__18399));
    InMux I__3669 (
            .O(N__18403),
            .I(N__18389));
    InMux I__3668 (
            .O(N__18402),
            .I(N__18389));
    InMux I__3667 (
            .O(N__18399),
            .I(N__18389));
    InMux I__3666 (
            .O(N__18398),
            .I(N__18389));
    LocalMux I__3665 (
            .O(N__18389),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    InMux I__3664 (
            .O(N__18386),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__3663 (
            .O(N__18383),
            .I(N__18374));
    InMux I__3662 (
            .O(N__18382),
            .I(N__18374));
    InMux I__3661 (
            .O(N__18381),
            .I(N__18374));
    LocalMux I__3660 (
            .O(N__18374),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1));
    InMux I__3659 (
            .O(N__18371),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__3658 (
            .O(N__18368),
            .I(N__18364));
    InMux I__3657 (
            .O(N__18367),
            .I(N__18361));
    LocalMux I__3656 (
            .O(N__18364),
            .I(N__18354));
    LocalMux I__3655 (
            .O(N__18361),
            .I(N__18354));
    InMux I__3654 (
            .O(N__18360),
            .I(N__18351));
    InMux I__3653 (
            .O(N__18359),
            .I(N__18348));
    Span4Mux_v I__3652 (
            .O(N__18354),
            .I(N__18343));
    LocalMux I__3651 (
            .O(N__18351),
            .I(N__18343));
    LocalMux I__3650 (
            .O(N__18348),
            .I(beamXZ0Z_8));
    Odrv4 I__3649 (
            .O(N__18343),
            .I(beamXZ0Z_8));
    InMux I__3648 (
            .O(N__18338),
            .I(bfn_8_4_0_));
    InMux I__3647 (
            .O(N__18335),
            .I(N__18331));
    InMux I__3646 (
            .O(N__18334),
            .I(N__18328));
    LocalMux I__3645 (
            .O(N__18331),
            .I(N__18321));
    LocalMux I__3644 (
            .O(N__18328),
            .I(N__18321));
    InMux I__3643 (
            .O(N__18327),
            .I(N__18318));
    InMux I__3642 (
            .O(N__18326),
            .I(N__18315));
    Span4Mux_v I__3641 (
            .O(N__18321),
            .I(N__18310));
    LocalMux I__3640 (
            .O(N__18318),
            .I(N__18310));
    LocalMux I__3639 (
            .O(N__18315),
            .I(beamXZ0Z_9));
    Odrv4 I__3638 (
            .O(N__18310),
            .I(beamXZ0Z_9));
    InMux I__3637 (
            .O(N__18305),
            .I(un5_visiblex_cry_8));
    CascadeMux I__3636 (
            .O(N__18302),
            .I(CO3_0_cascade_));
    InMux I__3635 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__3634 (
            .O(N__18296),
            .I(charx_if_generate_plus_mult1_un26_sum_s_2_sf));
    InMux I__3633 (
            .O(N__18293),
            .I(N__18288));
    InMux I__3632 (
            .O(N__18292),
            .I(N__18280));
    InMux I__3631 (
            .O(N__18291),
            .I(N__18277));
    LocalMux I__3630 (
            .O(N__18288),
            .I(N__18274));
    InMux I__3629 (
            .O(N__18287),
            .I(N__18271));
    InMux I__3628 (
            .O(N__18286),
            .I(N__18266));
    InMux I__3627 (
            .O(N__18285),
            .I(N__18266));
    InMux I__3626 (
            .O(N__18284),
            .I(N__18263));
    CascadeMux I__3625 (
            .O(N__18283),
            .I(N__18257));
    LocalMux I__3624 (
            .O(N__18280),
            .I(N__18250));
    LocalMux I__3623 (
            .O(N__18277),
            .I(N__18247));
    Span4Mux_v I__3622 (
            .O(N__18274),
            .I(N__18242));
    LocalMux I__3621 (
            .O(N__18271),
            .I(N__18242));
    LocalMux I__3620 (
            .O(N__18266),
            .I(N__18237));
    LocalMux I__3619 (
            .O(N__18263),
            .I(N__18237));
    InMux I__3618 (
            .O(N__18262),
            .I(N__18230));
    InMux I__3617 (
            .O(N__18261),
            .I(N__18230));
    InMux I__3616 (
            .O(N__18260),
            .I(N__18230));
    InMux I__3615 (
            .O(N__18257),
            .I(N__18227));
    InMux I__3614 (
            .O(N__18256),
            .I(N__18213));
    InMux I__3613 (
            .O(N__18255),
            .I(N__18213));
    InMux I__3612 (
            .O(N__18254),
            .I(N__18213));
    InMux I__3611 (
            .O(N__18253),
            .I(N__18213));
    Span4Mux_h I__3610 (
            .O(N__18250),
            .I(N__18202));
    Span4Mux_v I__3609 (
            .O(N__18247),
            .I(N__18202));
    Span4Mux_h I__3608 (
            .O(N__18242),
            .I(N__18202));
    Span4Mux_v I__3607 (
            .O(N__18237),
            .I(N__18202));
    LocalMux I__3606 (
            .O(N__18230),
            .I(N__18202));
    LocalMux I__3605 (
            .O(N__18227),
            .I(N__18199));
    InMux I__3604 (
            .O(N__18226),
            .I(N__18196));
    InMux I__3603 (
            .O(N__18225),
            .I(N__18193));
    InMux I__3602 (
            .O(N__18224),
            .I(N__18186));
    InMux I__3601 (
            .O(N__18223),
            .I(N__18186));
    InMux I__3600 (
            .O(N__18222),
            .I(N__18186));
    LocalMux I__3599 (
            .O(N__18213),
            .I(N__18183));
    Odrv4 I__3598 (
            .O(N__18202),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__3597 (
            .O(N__18199),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__3596 (
            .O(N__18196),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__3595 (
            .O(N__18193),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__3594 (
            .O(N__18186),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__3593 (
            .O(N__18183),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    InMux I__3592 (
            .O(N__18170),
            .I(N__18165));
    CascadeMux I__3591 (
            .O(N__18169),
            .I(N__18159));
    InMux I__3590 (
            .O(N__18168),
            .I(N__18154));
    LocalMux I__3589 (
            .O(N__18165),
            .I(N__18151));
    InMux I__3588 (
            .O(N__18164),
            .I(N__18146));
    InMux I__3587 (
            .O(N__18163),
            .I(N__18146));
    InMux I__3586 (
            .O(N__18162),
            .I(N__18143));
    InMux I__3585 (
            .O(N__18159),
            .I(N__18132));
    InMux I__3584 (
            .O(N__18158),
            .I(N__18129));
    InMux I__3583 (
            .O(N__18157),
            .I(N__18126));
    LocalMux I__3582 (
            .O(N__18154),
            .I(N__18121));
    Span4Mux_v I__3581 (
            .O(N__18151),
            .I(N__18121));
    LocalMux I__3580 (
            .O(N__18146),
            .I(N__18116));
    LocalMux I__3579 (
            .O(N__18143),
            .I(N__18116));
    InMux I__3578 (
            .O(N__18142),
            .I(N__18109));
    InMux I__3577 (
            .O(N__18141),
            .I(N__18109));
    InMux I__3576 (
            .O(N__18140),
            .I(N__18109));
    CascadeMux I__3575 (
            .O(N__18139),
            .I(N__18103));
    InMux I__3574 (
            .O(N__18138),
            .I(N__18093));
    InMux I__3573 (
            .O(N__18137),
            .I(N__18093));
    InMux I__3572 (
            .O(N__18136),
            .I(N__18093));
    InMux I__3571 (
            .O(N__18135),
            .I(N__18093));
    LocalMux I__3570 (
            .O(N__18132),
            .I(N__18088));
    LocalMux I__3569 (
            .O(N__18129),
            .I(N__18088));
    LocalMux I__3568 (
            .O(N__18126),
            .I(N__18085));
    Span4Mux_h I__3567 (
            .O(N__18121),
            .I(N__18078));
    Span4Mux_v I__3566 (
            .O(N__18116),
            .I(N__18078));
    LocalMux I__3565 (
            .O(N__18109),
            .I(N__18078));
    InMux I__3564 (
            .O(N__18108),
            .I(N__18073));
    InMux I__3563 (
            .O(N__18107),
            .I(N__18073));
    InMux I__3562 (
            .O(N__18106),
            .I(N__18066));
    InMux I__3561 (
            .O(N__18103),
            .I(N__18066));
    InMux I__3560 (
            .O(N__18102),
            .I(N__18066));
    LocalMux I__3559 (
            .O(N__18093),
            .I(N__18063));
    Odrv12 I__3558 (
            .O(N__18088),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__3557 (
            .O(N__18085),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__3556 (
            .O(N__18078),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    LocalMux I__3555 (
            .O(N__18073),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    LocalMux I__3554 (
            .O(N__18066),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__3553 (
            .O(N__18063),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    CascadeMux I__3552 (
            .O(N__18050),
            .I(N__18047));
    InMux I__3551 (
            .O(N__18047),
            .I(N__18044));
    LocalMux I__3550 (
            .O(N__18044),
            .I(N_13));
    CascadeMux I__3549 (
            .O(N__18041),
            .I(N__18038));
    InMux I__3548 (
            .O(N__18038),
            .I(N__18035));
    LocalMux I__3547 (
            .O(N__18035),
            .I(N__18032));
    Span4Mux_h I__3546 (
            .O(N__18032),
            .I(N__18029));
    Odrv4 I__3545 (
            .O(N__18029),
            .I(un113_pixel_4_0_15__un4_rowZ0Z_1));
    InMux I__3544 (
            .O(N__18026),
            .I(N__18023));
    LocalMux I__3543 (
            .O(N__18023),
            .I(N__18020));
    Span4Mux_h I__3542 (
            .O(N__18020),
            .I(N__18017));
    Span4Mux_h I__3541 (
            .O(N__18017),
            .I(N__18014));
    Span4Mux_v I__3540 (
            .O(N__18014),
            .I(N__18011));
    Odrv4 I__3539 (
            .O(N__18011),
            .I(un1_voltage_0_axb_0));
    InMux I__3538 (
            .O(N__18008),
            .I(N__18005));
    LocalMux I__3537 (
            .O(N__18005),
            .I(N__18002));
    Span4Mux_h I__3536 (
            .O(N__18002),
            .I(N__17999));
    Span4Mux_v I__3535 (
            .O(N__17999),
            .I(N__17996));
    Span4Mux_h I__3534 (
            .O(N__17996),
            .I(N__17993));
    Odrv4 I__3533 (
            .O(N__17993),
            .I(voltage_0_10_iv_0_0));
    InMux I__3532 (
            .O(N__17990),
            .I(N__17984));
    InMux I__3531 (
            .O(N__17989),
            .I(N__17984));
    LocalMux I__3530 (
            .O(N__17984),
            .I(N__17980));
    CascadeMux I__3529 (
            .O(N__17983),
            .I(N__17977));
    Span4Mux_h I__3528 (
            .O(N__17980),
            .I(N__17973));
    InMux I__3527 (
            .O(N__17977),
            .I(N__17970));
    InMux I__3526 (
            .O(N__17976),
            .I(N__17967));
    Span4Mux_h I__3525 (
            .O(N__17973),
            .I(N__17964));
    LocalMux I__3524 (
            .O(N__17970),
            .I(un1_voltage_012_2_0));
    LocalMux I__3523 (
            .O(N__17967),
            .I(un1_voltage_012_2_0));
    Odrv4 I__3522 (
            .O(N__17964),
            .I(un1_voltage_012_2_0));
    InMux I__3521 (
            .O(N__17957),
            .I(N__17954));
    LocalMux I__3520 (
            .O(N__17954),
            .I(N__17951));
    Span12Mux_s10_h I__3519 (
            .O(N__17951),
            .I(N__17948));
    Odrv12 I__3518 (
            .O(N__17948),
            .I(voltage_0_10_iv_0_1));
    InMux I__3517 (
            .O(N__17945),
            .I(N__17942));
    LocalMux I__3516 (
            .O(N__17942),
            .I(N__17939));
    Span12Mux_s8_v I__3515 (
            .O(N__17939),
            .I(N__17936));
    Odrv12 I__3514 (
            .O(N__17936),
            .I(voltage_0_RNO_0Z0Z_1));
    IoInMux I__3513 (
            .O(N__17933),
            .I(N__17929));
    IoInMux I__3512 (
            .O(N__17932),
            .I(N__17926));
    LocalMux I__3511 (
            .O(N__17929),
            .I(N__17921));
    LocalMux I__3510 (
            .O(N__17926),
            .I(N__17921));
    Span4Mux_s3_v I__3509 (
            .O(N__17921),
            .I(N__17918));
    Span4Mux_v I__3508 (
            .O(N__17918),
            .I(N__17915));
    Span4Mux_v I__3507 (
            .O(N__17915),
            .I(N__17911));
    InMux I__3506 (
            .O(N__17914),
            .I(N__17908));
    Odrv4 I__3505 (
            .O(N__17911),
            .I(nCS1_c));
    LocalMux I__3504 (
            .O(N__17908),
            .I(nCS1_c));
    InMux I__3503 (
            .O(N__17903),
            .I(N__17897));
    InMux I__3502 (
            .O(N__17902),
            .I(N__17892));
    InMux I__3501 (
            .O(N__17901),
            .I(N__17892));
    InMux I__3500 (
            .O(N__17900),
            .I(N__17888));
    LocalMux I__3499 (
            .O(N__17897),
            .I(N__17885));
    LocalMux I__3498 (
            .O(N__17892),
            .I(N__17882));
    InMux I__3497 (
            .O(N__17891),
            .I(N__17879));
    LocalMux I__3496 (
            .O(N__17888),
            .I(beamXZ0Z_1));
    Odrv4 I__3495 (
            .O(N__17885),
            .I(beamXZ0Z_1));
    Odrv4 I__3494 (
            .O(N__17882),
            .I(beamXZ0Z_1));
    LocalMux I__3493 (
            .O(N__17879),
            .I(beamXZ0Z_1));
    InMux I__3492 (
            .O(N__17870),
            .I(un5_visiblex_cry_0));
    InMux I__3491 (
            .O(N__17867),
            .I(N__17861));
    InMux I__3490 (
            .O(N__17866),
            .I(N__17861));
    LocalMux I__3489 (
            .O(N__17861),
            .I(N__17856));
    InMux I__3488 (
            .O(N__17860),
            .I(N__17853));
    InMux I__3487 (
            .O(N__17859),
            .I(N__17850));
    Span4Mux_v I__3486 (
            .O(N__17856),
            .I(N__17847));
    LocalMux I__3485 (
            .O(N__17853),
            .I(N__17844));
    LocalMux I__3484 (
            .O(N__17850),
            .I(beamXZ0Z_2));
    Odrv4 I__3483 (
            .O(N__17847),
            .I(beamXZ0Z_2));
    Odrv4 I__3482 (
            .O(N__17844),
            .I(beamXZ0Z_2));
    InMux I__3481 (
            .O(N__17837),
            .I(un5_visiblex_cry_1));
    InMux I__3480 (
            .O(N__17834),
            .I(N__17831));
    LocalMux I__3479 (
            .O(N__17831),
            .I(N__17825));
    InMux I__3478 (
            .O(N__17830),
            .I(N__17820));
    InMux I__3477 (
            .O(N__17829),
            .I(N__17820));
    InMux I__3476 (
            .O(N__17828),
            .I(N__17816));
    Span4Mux_v I__3475 (
            .O(N__17825),
            .I(N__17811));
    LocalMux I__3474 (
            .O(N__17820),
            .I(N__17811));
    InMux I__3473 (
            .O(N__17819),
            .I(N__17808));
    LocalMux I__3472 (
            .O(N__17816),
            .I(N__17803));
    Span4Mux_v I__3471 (
            .O(N__17811),
            .I(N__17803));
    LocalMux I__3470 (
            .O(N__17808),
            .I(N__17800));
    Odrv4 I__3469 (
            .O(N__17803),
            .I(beamXZ0Z_3));
    Odrv4 I__3468 (
            .O(N__17800),
            .I(beamXZ0Z_3));
    InMux I__3467 (
            .O(N__17795),
            .I(un5_visiblex_cry_2));
    CascadeMux I__3466 (
            .O(N__17792),
            .I(N__17787));
    CascadeMux I__3465 (
            .O(N__17791),
            .I(N__17784));
    CascadeMux I__3464 (
            .O(N__17790),
            .I(N__17780));
    InMux I__3463 (
            .O(N__17787),
            .I(N__17777));
    InMux I__3462 (
            .O(N__17784),
            .I(N__17772));
    InMux I__3461 (
            .O(N__17783),
            .I(N__17772));
    InMux I__3460 (
            .O(N__17780),
            .I(N__17769));
    LocalMux I__3459 (
            .O(N__17777),
            .I(N__17764));
    LocalMux I__3458 (
            .O(N__17772),
            .I(N__17764));
    LocalMux I__3457 (
            .O(N__17769),
            .I(N__17759));
    Span4Mux_h I__3456 (
            .O(N__17764),
            .I(N__17756));
    InMux I__3455 (
            .O(N__17763),
            .I(N__17753));
    InMux I__3454 (
            .O(N__17762),
            .I(N__17750));
    Span4Mux_v I__3453 (
            .O(N__17759),
            .I(N__17747));
    Span4Mux_v I__3452 (
            .O(N__17756),
            .I(N__17744));
    LocalMux I__3451 (
            .O(N__17753),
            .I(N__17741));
    LocalMux I__3450 (
            .O(N__17750),
            .I(beamXZ0Z_4));
    Odrv4 I__3449 (
            .O(N__17747),
            .I(beamXZ0Z_4));
    Odrv4 I__3448 (
            .O(N__17744),
            .I(beamXZ0Z_4));
    Odrv4 I__3447 (
            .O(N__17741),
            .I(beamXZ0Z_4));
    InMux I__3446 (
            .O(N__17732),
            .I(un5_visiblex_cry_3));
    InMux I__3445 (
            .O(N__17729),
            .I(N__17717));
    InMux I__3444 (
            .O(N__17728),
            .I(N__17717));
    InMux I__3443 (
            .O(N__17727),
            .I(N__17717));
    InMux I__3442 (
            .O(N__17726),
            .I(N__17717));
    LocalMux I__3441 (
            .O(N__17717),
            .I(N__17714));
    Span4Mux_v I__3440 (
            .O(N__17714),
            .I(N__17709));
    InMux I__3439 (
            .O(N__17713),
            .I(N__17706));
    InMux I__3438 (
            .O(N__17712),
            .I(N__17703));
    Span4Mux_v I__3437 (
            .O(N__17709),
            .I(N__17700));
    LocalMux I__3436 (
            .O(N__17706),
            .I(N__17697));
    LocalMux I__3435 (
            .O(N__17703),
            .I(beamXZ0Z_5));
    Odrv4 I__3434 (
            .O(N__17700),
            .I(beamXZ0Z_5));
    Odrv4 I__3433 (
            .O(N__17697),
            .I(beamXZ0Z_5));
    InMux I__3432 (
            .O(N__17690),
            .I(un5_visiblex_cry_4));
    CascadeMux I__3431 (
            .O(N__17687),
            .I(N__17681));
    InMux I__3430 (
            .O(N__17686),
            .I(N__17676));
    InMux I__3429 (
            .O(N__17685),
            .I(N__17673));
    InMux I__3428 (
            .O(N__17684),
            .I(N__17668));
    InMux I__3427 (
            .O(N__17681),
            .I(N__17668));
    InMux I__3426 (
            .O(N__17680),
            .I(N__17665));
    CascadeMux I__3425 (
            .O(N__17679),
            .I(N__17662));
    LocalMux I__3424 (
            .O(N__17676),
            .I(N__17658));
    LocalMux I__3423 (
            .O(N__17673),
            .I(N__17653));
    LocalMux I__3422 (
            .O(N__17668),
            .I(N__17653));
    LocalMux I__3421 (
            .O(N__17665),
            .I(N__17650));
    InMux I__3420 (
            .O(N__17662),
            .I(N__17647));
    InMux I__3419 (
            .O(N__17661),
            .I(N__17644));
    Span4Mux_v I__3418 (
            .O(N__17658),
            .I(N__17641));
    Span12Mux_s7_h I__3417 (
            .O(N__17653),
            .I(N__17638));
    Span4Mux_v I__3416 (
            .O(N__17650),
            .I(N__17633));
    LocalMux I__3415 (
            .O(N__17647),
            .I(N__17633));
    LocalMux I__3414 (
            .O(N__17644),
            .I(beamXZ0Z_6));
    Odrv4 I__3413 (
            .O(N__17641),
            .I(beamXZ0Z_6));
    Odrv12 I__3412 (
            .O(N__17638),
            .I(beamXZ0Z_6));
    Odrv4 I__3411 (
            .O(N__17633),
            .I(beamXZ0Z_6));
    InMux I__3410 (
            .O(N__17624),
            .I(un5_visiblex_cry_5));
    CascadeMux I__3409 (
            .O(N__17621),
            .I(N__17616));
    CascadeMux I__3408 (
            .O(N__17620),
            .I(N__17611));
    InMux I__3407 (
            .O(N__17619),
            .I(N__17608));
    InMux I__3406 (
            .O(N__17616),
            .I(N__17601));
    InMux I__3405 (
            .O(N__17615),
            .I(N__17601));
    InMux I__3404 (
            .O(N__17614),
            .I(N__17601));
    InMux I__3403 (
            .O(N__17611),
            .I(N__17598));
    LocalMux I__3402 (
            .O(N__17608),
            .I(N__17591));
    LocalMux I__3401 (
            .O(N__17601),
            .I(N__17591));
    LocalMux I__3400 (
            .O(N__17598),
            .I(N__17588));
    InMux I__3399 (
            .O(N__17597),
            .I(N__17585));
    InMux I__3398 (
            .O(N__17596),
            .I(N__17582));
    Span12Mux_v I__3397 (
            .O(N__17591),
            .I(N__17579));
    Span4Mux_v I__3396 (
            .O(N__17588),
            .I(N__17576));
    LocalMux I__3395 (
            .O(N__17585),
            .I(N__17573));
    LocalMux I__3394 (
            .O(N__17582),
            .I(beamXZ0Z_7));
    Odrv12 I__3393 (
            .O(N__17579),
            .I(beamXZ0Z_7));
    Odrv4 I__3392 (
            .O(N__17576),
            .I(beamXZ0Z_7));
    Odrv4 I__3391 (
            .O(N__17573),
            .I(beamXZ0Z_7));
    InMux I__3390 (
            .O(N__17564),
            .I(un5_visiblex_cry_6));
    InMux I__3389 (
            .O(N__17561),
            .I(un8_beamx_cry_4));
    InMux I__3388 (
            .O(N__17558),
            .I(un8_beamx_cry_5));
    InMux I__3387 (
            .O(N__17555),
            .I(un8_beamx_cry_6));
    InMux I__3386 (
            .O(N__17552),
            .I(un8_beamx_cry_7));
    InMux I__3385 (
            .O(N__17549),
            .I(bfn_8_2_0_));
    CEMux I__3384 (
            .O(N__17546),
            .I(N__17542));
    InMux I__3383 (
            .O(N__17545),
            .I(N__17537));
    LocalMux I__3382 (
            .O(N__17542),
            .I(N__17534));
    CEMux I__3381 (
            .O(N__17541),
            .I(N__17530));
    InMux I__3380 (
            .O(N__17540),
            .I(N__17526));
    LocalMux I__3379 (
            .O(N__17537),
            .I(N__17523));
    Span4Mux_v I__3378 (
            .O(N__17534),
            .I(N__17520));
    InMux I__3377 (
            .O(N__17533),
            .I(N__17516));
    LocalMux I__3376 (
            .O(N__17530),
            .I(N__17513));
    InMux I__3375 (
            .O(N__17529),
            .I(N__17510));
    LocalMux I__3374 (
            .O(N__17526),
            .I(N__17507));
    Span4Mux_h I__3373 (
            .O(N__17523),
            .I(N__17504));
    Span4Mux_s1_h I__3372 (
            .O(N__17520),
            .I(N__17501));
    InMux I__3371 (
            .O(N__17519),
            .I(N__17498));
    LocalMux I__3370 (
            .O(N__17516),
            .I(N__17495));
    Span4Mux_s2_h I__3369 (
            .O(N__17513),
            .I(N__17492));
    LocalMux I__3368 (
            .O(N__17510),
            .I(N__17487));
    Span4Mux_h I__3367 (
            .O(N__17507),
            .I(N__17487));
    Span4Mux_v I__3366 (
            .O(N__17504),
            .I(N__17482));
    Span4Mux_h I__3365 (
            .O(N__17501),
            .I(N__17482));
    LocalMux I__3364 (
            .O(N__17498),
            .I(un3_beamx_0));
    Odrv4 I__3363 (
            .O(N__17495),
            .I(un3_beamx_0));
    Odrv4 I__3362 (
            .O(N__17492),
            .I(un3_beamx_0));
    Odrv4 I__3361 (
            .O(N__17487),
            .I(un3_beamx_0));
    Odrv4 I__3360 (
            .O(N__17482),
            .I(un3_beamx_0));
    InMux I__3359 (
            .O(N__17471),
            .I(un8_beamx_cry_9));
    InMux I__3358 (
            .O(N__17468),
            .I(N__17463));
    InMux I__3357 (
            .O(N__17467),
            .I(N__17459));
    InMux I__3356 (
            .O(N__17466),
            .I(N__17456));
    LocalMux I__3355 (
            .O(N__17463),
            .I(N__17453));
    InMux I__3354 (
            .O(N__17462),
            .I(N__17450));
    LocalMux I__3353 (
            .O(N__17459),
            .I(N__17445));
    LocalMux I__3352 (
            .O(N__17456),
            .I(N__17445));
    Span4Mux_h I__3351 (
            .O(N__17453),
            .I(N__17442));
    LocalMux I__3350 (
            .O(N__17450),
            .I(N__17437));
    Span4Mux_v I__3349 (
            .O(N__17445),
            .I(N__17437));
    Span4Mux_v I__3348 (
            .O(N__17442),
            .I(N__17434));
    Odrv4 I__3347 (
            .O(N__17437),
            .I(beamXZ0Z_10));
    Odrv4 I__3346 (
            .O(N__17434),
            .I(beamXZ0Z_10));
    InMux I__3345 (
            .O(N__17429),
            .I(N__17426));
    LocalMux I__3344 (
            .O(N__17426),
            .I(ScreenBuffer_0_7_RNIHMH43T2Z0Z_0));
    CascadeMux I__3343 (
            .O(N__17423),
            .I(beamY_RNIDQUNU91Z0Z_0_cascade_));
    CascadeMux I__3342 (
            .O(N__17420),
            .I(un115_pixel_2_sn_5_cascade_));
    CascadeMux I__3341 (
            .O(N__17417),
            .I(un112_pixel_7_cascade_));
    InMux I__3340 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__3339 (
            .O(N__17411),
            .I(beamY_RNIINK7J73Z0Z_0));
    InMux I__3338 (
            .O(N__17408),
            .I(un8_beamx_cry_1));
    InMux I__3337 (
            .O(N__17405),
            .I(un8_beamx_cry_2));
    InMux I__3336 (
            .O(N__17402),
            .I(un8_beamx_cry_3));
    InMux I__3335 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__3334 (
            .O(N__17396),
            .I(N__17393));
    Odrv12 I__3333 (
            .O(N__17393),
            .I(slaveselect_RNILOQC2Z0Z_0));
    InMux I__3332 (
            .O(N__17390),
            .I(N__17386));
    InMux I__3331 (
            .O(N__17389),
            .I(N__17383));
    LocalMux I__3330 (
            .O(N__17386),
            .I(N__17380));
    LocalMux I__3329 (
            .O(N__17383),
            .I(ScreenBuffer_1_2Z0Z_4));
    Odrv4 I__3328 (
            .O(N__17380),
            .I(ScreenBuffer_1_2Z0Z_4));
    InMux I__3327 (
            .O(N__17375),
            .I(N__17372));
    LocalMux I__3326 (
            .O(N__17372),
            .I(ScreenBuffer_1_3Z0Z_2));
    InMux I__3325 (
            .O(N__17369),
            .I(N__17366));
    LocalMux I__3324 (
            .O(N__17366),
            .I(N__17363));
    Span4Mux_v I__3323 (
            .O(N__17363),
            .I(N__17360));
    Span4Mux_h I__3322 (
            .O(N__17360),
            .I(N__17357));
    Odrv4 I__3321 (
            .O(N__17357),
            .I(ScreenBuffer_1_0Z0Z_2));
    CascadeMux I__3320 (
            .O(N__17354),
            .I(un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_));
    CascadeMux I__3319 (
            .O(N__17351),
            .I(un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_));
    InMux I__3318 (
            .O(N__17348),
            .I(N__17345));
    LocalMux I__3317 (
            .O(N__17345),
            .I(m10_0_x1));
    CascadeMux I__3316 (
            .O(N__17342),
            .I(un112_pixel_2_2_cascade_));
    InMux I__3315 (
            .O(N__17339),
            .I(N__17336));
    LocalMux I__3314 (
            .O(N__17336),
            .I(un113_pixel_3_0_11__g0_0Z0Z_0));
    InMux I__3313 (
            .O(N__17333),
            .I(N__17329));
    InMux I__3312 (
            .O(N__17332),
            .I(N__17326));
    LocalMux I__3311 (
            .O(N__17329),
            .I(N__17323));
    LocalMux I__3310 (
            .O(N__17326),
            .I(N__17318));
    Span4Mux_v I__3309 (
            .O(N__17323),
            .I(N__17318));
    Odrv4 I__3308 (
            .O(N__17318),
            .I(ScreenBuffer_1_3Z0Z_4));
    InMux I__3307 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__3306 (
            .O(N__17312),
            .I(ScreenBuffer_1_3_RNIVS9G2FZ0Z_4));
    CascadeMux I__3305 (
            .O(N__17309),
            .I(g1Z0Z_1_cascade_));
    CascadeMux I__3304 (
            .O(N__17306),
            .I(N_1428_0_cascade_));
    CascadeMux I__3303 (
            .O(N__17303),
            .I(un113_pixel_4_0_15__g1_1_cascade_));
    InMux I__3302 (
            .O(N__17300),
            .I(N__17297));
    LocalMux I__3301 (
            .O(N__17297),
            .I(N_1300_0));
    CascadeMux I__3300 (
            .O(N__17294),
            .I(un112_pixel_0_2_cascade_));
    InMux I__3299 (
            .O(N__17291),
            .I(N__17288));
    LocalMux I__3298 (
            .O(N__17288),
            .I(N_1293_0));
    CascadeMux I__3297 (
            .O(N__17285),
            .I(ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_));
    CascadeMux I__3296 (
            .O(N__17282),
            .I(ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_));
    InMux I__3295 (
            .O(N__17279),
            .I(N__17273));
    InMux I__3294 (
            .O(N__17278),
            .I(N__17273));
    LocalMux I__3293 (
            .O(N__17273),
            .I(N__17270));
    Span12Mux_s7_h I__3292 (
            .O(N__17270),
            .I(N__17267));
    Odrv12 I__3291 (
            .O(N__17267),
            .I(row_1_if_generate_plus_mult1_un75_sum_c5));
    CascadeMux I__3290 (
            .O(N__17264),
            .I(N__17261));
    InMux I__3289 (
            .O(N__17261),
            .I(N__17255));
    InMux I__3288 (
            .O(N__17260),
            .I(N__17255));
    LocalMux I__3287 (
            .O(N__17255),
            .I(N__17252));
    Span4Mux_v I__3286 (
            .O(N__17252),
            .I(N__17248));
    InMux I__3285 (
            .O(N__17251),
            .I(N__17245));
    Sp12to4 I__3284 (
            .O(N__17248),
            .I(N__17240));
    LocalMux I__3283 (
            .O(N__17245),
            .I(N__17240));
    Odrv12 I__3282 (
            .O(N__17240),
            .I(row_1_if_generate_plus_mult1_un68_sum_cZ0Z4));
    InMux I__3281 (
            .O(N__17237),
            .I(N__17231));
    InMux I__3280 (
            .O(N__17236),
            .I(N__17231));
    LocalMux I__3279 (
            .O(N__17231),
            .I(N__17228));
    Span4Mux_h I__3278 (
            .O(N__17228),
            .I(N__17225));
    Span4Mux_h I__3277 (
            .O(N__17225),
            .I(N__17222));
    Odrv4 I__3276 (
            .O(N__17222),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_0));
    InMux I__3275 (
            .O(N__17219),
            .I(N__17216));
    LocalMux I__3274 (
            .O(N__17216),
            .I(ScreenBuffer_1_2Z0Z_0));
    CascadeMux I__3273 (
            .O(N__17213),
            .I(un3_rowlto1_cascade_));
    CascadeMux I__3272 (
            .O(N__17210),
            .I(N__17207));
    InMux I__3271 (
            .O(N__17207),
            .I(N__17203));
    InMux I__3270 (
            .O(N__17206),
            .I(N__17200));
    LocalMux I__3269 (
            .O(N__17203),
            .I(N__17197));
    LocalMux I__3268 (
            .O(N__17200),
            .I(N__17194));
    Odrv4 I__3267 (
            .O(N__17197),
            .I(ScreenBuffer_0_2Z0Z_0));
    Odrv4 I__3266 (
            .O(N__17194),
            .I(ScreenBuffer_0_2Z0Z_0));
    InMux I__3265 (
            .O(N__17189),
            .I(N__17186));
    LocalMux I__3264 (
            .O(N__17186),
            .I(N__17182));
    InMux I__3263 (
            .O(N__17185),
            .I(N__17179));
    Span4Mux_h I__3262 (
            .O(N__17182),
            .I(N__17176));
    LocalMux I__3261 (
            .O(N__17179),
            .I(N__17173));
    Odrv4 I__3260 (
            .O(N__17176),
            .I(ScreenBuffer_1_1_1_sqmuxa));
    Odrv4 I__3259 (
            .O(N__17173),
            .I(ScreenBuffer_1_1_1_sqmuxa));
    CascadeMux I__3258 (
            .O(N__17168),
            .I(N__17165));
    InMux I__3257 (
            .O(N__17165),
            .I(N__17161));
    InMux I__3256 (
            .O(N__17164),
            .I(N__17158));
    LocalMux I__3255 (
            .O(N__17161),
            .I(ScreenBuffer_0_0Z0Z_0));
    LocalMux I__3254 (
            .O(N__17158),
            .I(ScreenBuffer_0_0Z0Z_0));
    InMux I__3253 (
            .O(N__17153),
            .I(N__17150));
    LocalMux I__3252 (
            .O(N__17150),
            .I(N__17146));
    InMux I__3251 (
            .O(N__17149),
            .I(N__17143));
    Span4Mux_h I__3250 (
            .O(N__17146),
            .I(N__17140));
    LocalMux I__3249 (
            .O(N__17143),
            .I(ScreenBuffer_1_1Z0Z_4));
    Odrv4 I__3248 (
            .O(N__17140),
            .I(ScreenBuffer_1_1Z0Z_4));
    CascadeMux I__3247 (
            .O(N__17135),
            .I(ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_));
    InMux I__3246 (
            .O(N__17132),
            .I(N__17129));
    LocalMux I__3245 (
            .O(N__17129),
            .I(currentchar_1_11_ns_1_4));
    InMux I__3244 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__3243 (
            .O(N__17123),
            .I(ScreenBuffer_1_2_RNIUP6F2FZ0Z_4));
    InMux I__3242 (
            .O(N__17120),
            .I(N__17110));
    InMux I__3241 (
            .O(N__17119),
            .I(N__17107));
    InMux I__3240 (
            .O(N__17118),
            .I(N__17104));
    InMux I__3239 (
            .O(N__17117),
            .I(N__17101));
    InMux I__3238 (
            .O(N__17116),
            .I(N__17092));
    InMux I__3237 (
            .O(N__17115),
            .I(N__17092));
    InMux I__3236 (
            .O(N__17114),
            .I(N__17092));
    InMux I__3235 (
            .O(N__17113),
            .I(N__17092));
    LocalMux I__3234 (
            .O(N__17110),
            .I(N__17087));
    LocalMux I__3233 (
            .O(N__17107),
            .I(N__17087));
    LocalMux I__3232 (
            .O(N__17104),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3));
    LocalMux I__3231 (
            .O(N__17101),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3));
    LocalMux I__3230 (
            .O(N__17092),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3));
    Odrv4 I__3229 (
            .O(N__17087),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3));
    InMux I__3228 (
            .O(N__17078),
            .I(N__17074));
    CascadeMux I__3227 (
            .O(N__17077),
            .I(N__17070));
    LocalMux I__3226 (
            .O(N__17074),
            .I(N__17062));
    InMux I__3225 (
            .O(N__17073),
            .I(N__17057));
    InMux I__3224 (
            .O(N__17070),
            .I(N__17057));
    InMux I__3223 (
            .O(N__17069),
            .I(N__17054));
    InMux I__3222 (
            .O(N__17068),
            .I(N__17045));
    InMux I__3221 (
            .O(N__17067),
            .I(N__17045));
    InMux I__3220 (
            .O(N__17066),
            .I(N__17045));
    InMux I__3219 (
            .O(N__17065),
            .I(N__17045));
    Span4Mux_v I__3218 (
            .O(N__17062),
            .I(N__17040));
    LocalMux I__3217 (
            .O(N__17057),
            .I(N__17040));
    LocalMux I__3216 (
            .O(N__17054),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__3215 (
            .O(N__17045),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    Odrv4 I__3214 (
            .O(N__17040),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    CascadeMux I__3213 (
            .O(N__17033),
            .I(N_9_i_cascade_));
    InMux I__3212 (
            .O(N__17030),
            .I(N__17027));
    LocalMux I__3211 (
            .O(N__17027),
            .I(N_13_0));
    InMux I__3210 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__3209 (
            .O(N__17021),
            .I(N__17017));
    InMux I__3208 (
            .O(N__17020),
            .I(N__17014));
    Span4Mux_v I__3207 (
            .O(N__17017),
            .I(N__17011));
    LocalMux I__3206 (
            .O(N__17014),
            .I(ScreenBuffer_0_8Z0Z_0));
    Odrv4 I__3205 (
            .O(N__17011),
            .I(ScreenBuffer_0_8Z0Z_0));
    InMux I__3204 (
            .O(N__17006),
            .I(N__17003));
    LocalMux I__3203 (
            .O(N__17003),
            .I(N__17000));
    Odrv12 I__3202 (
            .O(N__17000),
            .I(ScreenBuffer_1_0Z0Z_0));
    CascadeMux I__3201 (
            .O(N__16997),
            .I(currentchar_1_9_ns_1_0_cascade_));
    InMux I__3200 (
            .O(N__16994),
            .I(N__16991));
    LocalMux I__3199 (
            .O(N__16991),
            .I(N__16988));
    Span4Mux_h I__3198 (
            .O(N__16988),
            .I(N__16985));
    Odrv4 I__3197 (
            .O(N__16985),
            .I(ScreenBuffer_1_1Z0Z_0));
    CascadeMux I__3196 (
            .O(N__16982),
            .I(currentchar_1_6_ns_1_0_cascade_));
    CascadeMux I__3195 (
            .O(N__16979),
            .I(N__16975));
    InMux I__3194 (
            .O(N__16978),
            .I(N__16972));
    InMux I__3193 (
            .O(N__16975),
            .I(N__16969));
    LocalMux I__3192 (
            .O(N__16972),
            .I(N__16966));
    LocalMux I__3191 (
            .O(N__16969),
            .I(N__16961));
    Span4Mux_v I__3190 (
            .O(N__16966),
            .I(N__16961));
    Odrv4 I__3189 (
            .O(N__16961),
            .I(ScreenBuffer_0_1Z0Z_0));
    InMux I__3188 (
            .O(N__16958),
            .I(N__16955));
    LocalMux I__3187 (
            .O(N__16955),
            .I(N__16951));
    InMux I__3186 (
            .O(N__16954),
            .I(N__16948));
    Span4Mux_v I__3185 (
            .O(N__16951),
            .I(N__16945));
    LocalMux I__3184 (
            .O(N__16948),
            .I(ScreenBuffer_1_0Z0Z_4));
    Odrv4 I__3183 (
            .O(N__16945),
            .I(ScreenBuffer_1_0Z0Z_4));
    CascadeMux I__3182 (
            .O(N__16940),
            .I(font_un3_pixel_28_cascade_));
    InMux I__3181 (
            .O(N__16937),
            .I(N__16933));
    InMux I__3180 (
            .O(N__16936),
            .I(N__16930));
    LocalMux I__3179 (
            .O(N__16933),
            .I(un113_pixel_4_0_15__un15_beamyZ0Z_2));
    LocalMux I__3178 (
            .O(N__16930),
            .I(un113_pixel_4_0_15__un15_beamyZ0Z_2));
    InMux I__3177 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__3176 (
            .O(N__16922),
            .I(N__16919));
    Span4Mux_h I__3175 (
            .O(N__16919),
            .I(N__16916));
    Odrv4 I__3174 (
            .O(N__16916),
            .I(un13_beamy));
    CascadeMux I__3173 (
            .O(N__16913),
            .I(font_un61_pixel_cascade_));
    InMux I__3172 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__3171 (
            .O(N__16907),
            .I(un4_row));
    InMux I__3170 (
            .O(N__16904),
            .I(N__16901));
    LocalMux I__3169 (
            .O(N__16901),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0));
    CascadeMux I__3168 (
            .O(N__16898),
            .I(N__16895));
    InMux I__3167 (
            .O(N__16895),
            .I(N__16892));
    LocalMux I__3166 (
            .O(N__16892),
            .I(N__16889));
    Span4Mux_v I__3165 (
            .O(N__16889),
            .I(N__16885));
    InMux I__3164 (
            .O(N__16888),
            .I(N__16882));
    Odrv4 I__3163 (
            .O(N__16885),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    LocalMux I__3162 (
            .O(N__16882),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    InMux I__3161 (
            .O(N__16877),
            .I(N__16871));
    InMux I__3160 (
            .O(N__16876),
            .I(N__16871));
    LocalMux I__3159 (
            .O(N__16871),
            .I(charx_23));
    InMux I__3158 (
            .O(N__16868),
            .I(N__16865));
    LocalMux I__3157 (
            .O(N__16865),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3));
    CascadeMux I__3156 (
            .O(N__16862),
            .I(N__16859));
    InMux I__3155 (
            .O(N__16859),
            .I(N__16856));
    LocalMux I__3154 (
            .O(N__16856),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0));
    InMux I__3153 (
            .O(N__16853),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__3152 (
            .O(N__16850),
            .I(N__16847));
    LocalMux I__3151 (
            .O(N__16847),
            .I(charx_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__3150 (
            .O(N__16844),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__3149 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__3148 (
            .O(N__16838),
            .I(un113_pixel_4_0_15__un18_beamylto9Z0Z_2));
    InMux I__3147 (
            .O(N__16835),
            .I(N__16830));
    InMux I__3146 (
            .O(N__16834),
            .I(N__16827));
    InMux I__3145 (
            .O(N__16833),
            .I(N__16824));
    LocalMux I__3144 (
            .O(N__16830),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    LocalMux I__3143 (
            .O(N__16827),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    LocalMux I__3142 (
            .O(N__16824),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    InMux I__3141 (
            .O(N__16817),
            .I(N__16811));
    InMux I__3140 (
            .O(N__16816),
            .I(N__16811));
    LocalMux I__3139 (
            .O(N__16811),
            .I(charx_if_generate_plus_mult1_un33_sum_i_5));
    InMux I__3138 (
            .O(N__16808),
            .I(N__16796));
    InMux I__3137 (
            .O(N__16807),
            .I(N__16796));
    InMux I__3136 (
            .O(N__16806),
            .I(N__16796));
    InMux I__3135 (
            .O(N__16805),
            .I(N__16796));
    LocalMux I__3134 (
            .O(N__16796),
            .I(un1_beamx_2));
    InMux I__3133 (
            .O(N__16793),
            .I(N__16790));
    LocalMux I__3132 (
            .O(N__16790),
            .I(charx_i_24));
    CascadeMux I__3131 (
            .O(N__16787),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_));
    CascadeMux I__3130 (
            .O(N__16784),
            .I(N__16781));
    InMux I__3129 (
            .O(N__16781),
            .I(N__16778));
    LocalMux I__3128 (
            .O(N__16778),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328));
    InMux I__3127 (
            .O(N__16775),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2));
    CascadeMux I__3126 (
            .O(N__16772),
            .I(N__16769));
    InMux I__3125 (
            .O(N__16769),
            .I(N__16766));
    LocalMux I__3124 (
            .O(N__16766),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538));
    InMux I__3123 (
            .O(N__16763),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_3));
    CascadeMux I__3122 (
            .O(N__16760),
            .I(N__16757));
    InMux I__3121 (
            .O(N__16757),
            .I(N__16754));
    LocalMux I__3120 (
            .O(N__16754),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO));
    InMux I__3119 (
            .O(N__16751),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4));
    InMux I__3118 (
            .O(N__16748),
            .I(N__16742));
    InMux I__3117 (
            .O(N__16747),
            .I(N__16742));
    LocalMux I__3116 (
            .O(N__16742),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    InMux I__3115 (
            .O(N__16739),
            .I(N__16735));
    InMux I__3114 (
            .O(N__16738),
            .I(N__16732));
    LocalMux I__3113 (
            .O(N__16735),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    LocalMux I__3112 (
            .O(N__16732),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    CascadeMux I__3111 (
            .O(N__16727),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_));
    InMux I__3110 (
            .O(N__16724),
            .I(N__16721));
    LocalMux I__3109 (
            .O(N__16721),
            .I(charx_if_generate_plus_mult1_un26_sum_i_5));
    CascadeMux I__3108 (
            .O(N__16718),
            .I(N__16715));
    InMux I__3107 (
            .O(N__16715),
            .I(N__16712));
    LocalMux I__3106 (
            .O(N__16712),
            .I(charx_if_generate_plus_mult1_un33_sum_i));
    InMux I__3105 (
            .O(N__16709),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1));
    CascadeMux I__3104 (
            .O(N__16706),
            .I(N__16703));
    InMux I__3103 (
            .O(N__16703),
            .I(N__16700));
    LocalMux I__3102 (
            .O(N__16700),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0));
    InMux I__3101 (
            .O(N__16697),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__3100 (
            .O(N__16694),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1));
    InMux I__3099 (
            .O(N__16691),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__3098 (
            .O(N__16688),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__3097 (
            .O(N__16685),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4));
    InMux I__3096 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__3095 (
            .O(N__16679),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_0));
    InMux I__3094 (
            .O(N__16676),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1));
    InMux I__3093 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__3092 (
            .O(N__16670),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__3091 (
            .O(N__16667),
            .I(N__16664));
    InMux I__3090 (
            .O(N__16664),
            .I(N__16661));
    LocalMux I__3089 (
            .O(N__16661),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0));
    InMux I__3088 (
            .O(N__16658),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__3087 (
            .O(N__16655),
            .I(N__16652));
    InMux I__3086 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__3085 (
            .O(N__16649),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91));
    InMux I__3084 (
            .O(N__16646),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__3083 (
            .O(N__16643),
            .I(N__16640));
    LocalMux I__3082 (
            .O(N__16640),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__3081 (
            .O(N__16637),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__3080 (
            .O(N__16634),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__3079 (
            .O(N__16631),
            .I(N__16626));
    InMux I__3078 (
            .O(N__16630),
            .I(N__16621));
    InMux I__3077 (
            .O(N__16629),
            .I(N__16621));
    LocalMux I__3076 (
            .O(N__16626),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1));
    LocalMux I__3075 (
            .O(N__16621),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1));
    InMux I__3074 (
            .O(N__16616),
            .I(N__16613));
    LocalMux I__3073 (
            .O(N__16613),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0));
    CascadeMux I__3072 (
            .O(N__16610),
            .I(N__16607));
    InMux I__3071 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__3070 (
            .O(N__16604),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i));
    CascadeMux I__3069 (
            .O(N__16601),
            .I(N__16598));
    InMux I__3068 (
            .O(N__16598),
            .I(N__16595));
    LocalMux I__3067 (
            .O(N__16595),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__3066 (
            .O(N__16592),
            .I(N__16589));
    LocalMux I__3065 (
            .O(N__16589),
            .I(N__16586));
    Span4Mux_v I__3064 (
            .O(N__16586),
            .I(N__16581));
    InMux I__3063 (
            .O(N__16585),
            .I(N__16578));
    InMux I__3062 (
            .O(N__16584),
            .I(N__16574));
    Span4Mux_h I__3061 (
            .O(N__16581),
            .I(N__16569));
    LocalMux I__3060 (
            .O(N__16578),
            .I(N__16569));
    InMux I__3059 (
            .O(N__16577),
            .I(N__16566));
    LocalMux I__3058 (
            .O(N__16574),
            .I(voltage_3Z0Z_2));
    Odrv4 I__3057 (
            .O(N__16569),
            .I(voltage_3Z0Z_2));
    LocalMux I__3056 (
            .O(N__16566),
            .I(voltage_3Z0Z_2));
    InMux I__3055 (
            .O(N__16559),
            .I(N__16556));
    LocalMux I__3054 (
            .O(N__16556),
            .I(N__16551));
    InMux I__3053 (
            .O(N__16555),
            .I(N__16548));
    CascadeMux I__3052 (
            .O(N__16554),
            .I(N__16545));
    Span4Mux_v I__3051 (
            .O(N__16551),
            .I(N__16538));
    LocalMux I__3050 (
            .O(N__16548),
            .I(N__16538));
    InMux I__3049 (
            .O(N__16545),
            .I(N__16535));
    InMux I__3048 (
            .O(N__16544),
            .I(N__16530));
    InMux I__3047 (
            .O(N__16543),
            .I(N__16530));
    Span4Mux_h I__3046 (
            .O(N__16538),
            .I(N__16527));
    LocalMux I__3045 (
            .O(N__16535),
            .I(voltage_0Z0Z_2));
    LocalMux I__3044 (
            .O(N__16530),
            .I(voltage_0Z0Z_2));
    Odrv4 I__3043 (
            .O(N__16527),
            .I(voltage_0Z0Z_2));
    InMux I__3042 (
            .O(N__16520),
            .I(N__16517));
    LocalMux I__3041 (
            .O(N__16517),
            .I(un1_sclk17_7_1));
    CascadeMux I__3040 (
            .O(N__16514),
            .I(N__16508));
    InMux I__3039 (
            .O(N__16513),
            .I(N__16500));
    InMux I__3038 (
            .O(N__16512),
            .I(N__16500));
    InMux I__3037 (
            .O(N__16511),
            .I(N__16500));
    InMux I__3036 (
            .O(N__16508),
            .I(N__16495));
    InMux I__3035 (
            .O(N__16507),
            .I(N__16492));
    LocalMux I__3034 (
            .O(N__16500),
            .I(N__16489));
    InMux I__3033 (
            .O(N__16499),
            .I(N__16486));
    InMux I__3032 (
            .O(N__16498),
            .I(N__16483));
    LocalMux I__3031 (
            .O(N__16495),
            .I(N__16473));
    LocalMux I__3030 (
            .O(N__16492),
            .I(N__16473));
    Span4Mux_v I__3029 (
            .O(N__16489),
            .I(N__16473));
    LocalMux I__3028 (
            .O(N__16486),
            .I(N__16473));
    LocalMux I__3027 (
            .O(N__16483),
            .I(N__16470));
    InMux I__3026 (
            .O(N__16482),
            .I(N__16467));
    Span4Mux_h I__3025 (
            .O(N__16473),
            .I(N__16463));
    Span4Mux_h I__3024 (
            .O(N__16470),
            .I(N__16458));
    LocalMux I__3023 (
            .O(N__16467),
            .I(N__16458));
    InMux I__3022 (
            .O(N__16466),
            .I(N__16455));
    Odrv4 I__3021 (
            .O(N__16463),
            .I(un5_slaveselect));
    Odrv4 I__3020 (
            .O(N__16458),
            .I(un5_slaveselect));
    LocalMux I__3019 (
            .O(N__16455),
            .I(un5_slaveselect));
    IoInMux I__3018 (
            .O(N__16448),
            .I(N__16445));
    LocalMux I__3017 (
            .O(N__16445),
            .I(N__16442));
    Span4Mux_s2_v I__3016 (
            .O(N__16442),
            .I(N__16438));
    InMux I__3015 (
            .O(N__16441),
            .I(N__16435));
    Odrv4 I__3014 (
            .O(N__16438),
            .I(SDATA2_c));
    LocalMux I__3013 (
            .O(N__16435),
            .I(SDATA2_c));
    CascadeMux I__3012 (
            .O(N__16430),
            .I(un1_sclk17_9_1_cascade_));
    CascadeMux I__3011 (
            .O(N__16427),
            .I(N__16420));
    CascadeMux I__3010 (
            .O(N__16426),
            .I(N__16417));
    CascadeMux I__3009 (
            .O(N__16425),
            .I(N__16414));
    CascadeMux I__3008 (
            .O(N__16424),
            .I(N__16411));
    CascadeMux I__3007 (
            .O(N__16423),
            .I(N__16403));
    InMux I__3006 (
            .O(N__16420),
            .I(N__16394));
    InMux I__3005 (
            .O(N__16417),
            .I(N__16394));
    InMux I__3004 (
            .O(N__16414),
            .I(N__16388));
    InMux I__3003 (
            .O(N__16411),
            .I(N__16388));
    InMux I__3002 (
            .O(N__16410),
            .I(N__16381));
    InMux I__3001 (
            .O(N__16409),
            .I(N__16381));
    InMux I__3000 (
            .O(N__16408),
            .I(N__16381));
    InMux I__2999 (
            .O(N__16407),
            .I(N__16378));
    InMux I__2998 (
            .O(N__16406),
            .I(N__16375));
    InMux I__2997 (
            .O(N__16403),
            .I(N__16366));
    InMux I__2996 (
            .O(N__16402),
            .I(N__16366));
    InMux I__2995 (
            .O(N__16401),
            .I(N__16366));
    InMux I__2994 (
            .O(N__16400),
            .I(N__16366));
    CascadeMux I__2993 (
            .O(N__16399),
            .I(N__16363));
    LocalMux I__2992 (
            .O(N__16394),
            .I(N__16357));
    InMux I__2991 (
            .O(N__16393),
            .I(N__16354));
    LocalMux I__2990 (
            .O(N__16388),
            .I(N__16351));
    LocalMux I__2989 (
            .O(N__16381),
            .I(N__16348));
    LocalMux I__2988 (
            .O(N__16378),
            .I(N__16341));
    LocalMux I__2987 (
            .O(N__16375),
            .I(N__16336));
    LocalMux I__2986 (
            .O(N__16366),
            .I(N__16336));
    InMux I__2985 (
            .O(N__16363),
            .I(N__16333));
    InMux I__2984 (
            .O(N__16362),
            .I(N__16328));
    InMux I__2983 (
            .O(N__16361),
            .I(N__16328));
    InMux I__2982 (
            .O(N__16360),
            .I(N__16325));
    Span4Mux_v I__2981 (
            .O(N__16357),
            .I(N__16316));
    LocalMux I__2980 (
            .O(N__16354),
            .I(N__16316));
    Span4Mux_s3_v I__2979 (
            .O(N__16351),
            .I(N__16316));
    Span4Mux_s3_v I__2978 (
            .O(N__16348),
            .I(N__16316));
    InMux I__2977 (
            .O(N__16347),
            .I(N__16311));
    InMux I__2976 (
            .O(N__16346),
            .I(N__16311));
    InMux I__2975 (
            .O(N__16345),
            .I(N__16306));
    InMux I__2974 (
            .O(N__16344),
            .I(N__16306));
    Span4Mux_v I__2973 (
            .O(N__16341),
            .I(N__16297));
    Span4Mux_s3_v I__2972 (
            .O(N__16336),
            .I(N__16297));
    LocalMux I__2971 (
            .O(N__16333),
            .I(N__16297));
    LocalMux I__2970 (
            .O(N__16328),
            .I(N__16297));
    LocalMux I__2969 (
            .O(N__16325),
            .I(counterZ0Z_3));
    Odrv4 I__2968 (
            .O(N__16316),
            .I(counterZ0Z_3));
    LocalMux I__2967 (
            .O(N__16311),
            .I(counterZ0Z_3));
    LocalMux I__2966 (
            .O(N__16306),
            .I(counterZ0Z_3));
    Odrv4 I__2965 (
            .O(N__16297),
            .I(counterZ0Z_3));
    CascadeMux I__2964 (
            .O(N__16286),
            .I(N__16279));
    InMux I__2963 (
            .O(N__16285),
            .I(N__16270));
    CascadeMux I__2962 (
            .O(N__16284),
            .I(N__16262));
    CascadeMux I__2961 (
            .O(N__16283),
            .I(N__16252));
    InMux I__2960 (
            .O(N__16282),
            .I(N__16234));
    InMux I__2959 (
            .O(N__16279),
            .I(N__16234));
    InMux I__2958 (
            .O(N__16278),
            .I(N__16234));
    InMux I__2957 (
            .O(N__16277),
            .I(N__16231));
    InMux I__2956 (
            .O(N__16276),
            .I(N__16224));
    InMux I__2955 (
            .O(N__16275),
            .I(N__16224));
    InMux I__2954 (
            .O(N__16274),
            .I(N__16224));
    InMux I__2953 (
            .O(N__16273),
            .I(N__16218));
    LocalMux I__2952 (
            .O(N__16270),
            .I(N__16209));
    InMux I__2951 (
            .O(N__16269),
            .I(N__16204));
    InMux I__2950 (
            .O(N__16268),
            .I(N__16204));
    InMux I__2949 (
            .O(N__16267),
            .I(N__16201));
    InMux I__2948 (
            .O(N__16266),
            .I(N__16198));
    InMux I__2947 (
            .O(N__16265),
            .I(N__16189));
    InMux I__2946 (
            .O(N__16262),
            .I(N__16189));
    InMux I__2945 (
            .O(N__16261),
            .I(N__16189));
    InMux I__2944 (
            .O(N__16260),
            .I(N__16189));
    InMux I__2943 (
            .O(N__16259),
            .I(N__16182));
    InMux I__2942 (
            .O(N__16258),
            .I(N__16182));
    InMux I__2941 (
            .O(N__16257),
            .I(N__16182));
    InMux I__2940 (
            .O(N__16256),
            .I(N__16174));
    InMux I__2939 (
            .O(N__16255),
            .I(N__16174));
    InMux I__2938 (
            .O(N__16252),
            .I(N__16174));
    InMux I__2937 (
            .O(N__16251),
            .I(N__16167));
    InMux I__2936 (
            .O(N__16250),
            .I(N__16167));
    InMux I__2935 (
            .O(N__16249),
            .I(N__16167));
    InMux I__2934 (
            .O(N__16248),
            .I(N__16160));
    InMux I__2933 (
            .O(N__16247),
            .I(N__16160));
    InMux I__2932 (
            .O(N__16246),
            .I(N__16160));
    InMux I__2931 (
            .O(N__16245),
            .I(N__16157));
    InMux I__2930 (
            .O(N__16244),
            .I(N__16154));
    InMux I__2929 (
            .O(N__16243),
            .I(N__16151));
    CascadeMux I__2928 (
            .O(N__16242),
            .I(N__16147));
    CascadeMux I__2927 (
            .O(N__16241),
            .I(N__16144));
    LocalMux I__2926 (
            .O(N__16234),
            .I(N__16141));
    LocalMux I__2925 (
            .O(N__16231),
            .I(N__16138));
    LocalMux I__2924 (
            .O(N__16224),
            .I(N__16135));
    InMux I__2923 (
            .O(N__16223),
            .I(N__16128));
    InMux I__2922 (
            .O(N__16222),
            .I(N__16128));
    InMux I__2921 (
            .O(N__16221),
            .I(N__16128));
    LocalMux I__2920 (
            .O(N__16218),
            .I(N__16125));
    InMux I__2919 (
            .O(N__16217),
            .I(N__16118));
    InMux I__2918 (
            .O(N__16216),
            .I(N__16118));
    InMux I__2917 (
            .O(N__16215),
            .I(N__16118));
    InMux I__2916 (
            .O(N__16214),
            .I(N__16113));
    InMux I__2915 (
            .O(N__16213),
            .I(N__16113));
    InMux I__2914 (
            .O(N__16212),
            .I(N__16110));
    Span4Mux_s3_h I__2913 (
            .O(N__16209),
            .I(N__16106));
    LocalMux I__2912 (
            .O(N__16204),
            .I(N__16101));
    LocalMux I__2911 (
            .O(N__16201),
            .I(N__16101));
    LocalMux I__2910 (
            .O(N__16198),
            .I(N__16098));
    LocalMux I__2909 (
            .O(N__16189),
            .I(N__16093));
    LocalMux I__2908 (
            .O(N__16182),
            .I(N__16093));
    InMux I__2907 (
            .O(N__16181),
            .I(N__16090));
    LocalMux I__2906 (
            .O(N__16174),
            .I(N__16085));
    LocalMux I__2905 (
            .O(N__16167),
            .I(N__16085));
    LocalMux I__2904 (
            .O(N__16160),
            .I(N__16080));
    LocalMux I__2903 (
            .O(N__16157),
            .I(N__16080));
    LocalMux I__2902 (
            .O(N__16154),
            .I(N__16075));
    LocalMux I__2901 (
            .O(N__16151),
            .I(N__16075));
    InMux I__2900 (
            .O(N__16150),
            .I(N__16072));
    InMux I__2899 (
            .O(N__16147),
            .I(N__16069));
    InMux I__2898 (
            .O(N__16144),
            .I(N__16066));
    Span4Mux_s3_h I__2897 (
            .O(N__16141),
            .I(N__16061));
    Span4Mux_s3_h I__2896 (
            .O(N__16138),
            .I(N__16061));
    Span4Mux_v I__2895 (
            .O(N__16135),
            .I(N__16054));
    LocalMux I__2894 (
            .O(N__16128),
            .I(N__16054));
    Span4Mux_s2_h I__2893 (
            .O(N__16125),
            .I(N__16054));
    LocalMux I__2892 (
            .O(N__16118),
            .I(N__16051));
    LocalMux I__2891 (
            .O(N__16113),
            .I(N__16048));
    LocalMux I__2890 (
            .O(N__16110),
            .I(N__16045));
    InMux I__2889 (
            .O(N__16109),
            .I(N__16042));
    Span4Mux_v I__2888 (
            .O(N__16106),
            .I(N__16037));
    Span4Mux_s3_h I__2887 (
            .O(N__16101),
            .I(N__16037));
    Span4Mux_h I__2886 (
            .O(N__16098),
            .I(N__16026));
    Span4Mux_s3_h I__2885 (
            .O(N__16093),
            .I(N__16026));
    LocalMux I__2884 (
            .O(N__16090),
            .I(N__16026));
    Span4Mux_s3_h I__2883 (
            .O(N__16085),
            .I(N__16026));
    Span4Mux_h I__2882 (
            .O(N__16080),
            .I(N__16026));
    Span12Mux_s3_h I__2881 (
            .O(N__16075),
            .I(N__16023));
    LocalMux I__2880 (
            .O(N__16072),
            .I(counterZ0Z_0));
    LocalMux I__2879 (
            .O(N__16069),
            .I(counterZ0Z_0));
    LocalMux I__2878 (
            .O(N__16066),
            .I(counterZ0Z_0));
    Odrv4 I__2877 (
            .O(N__16061),
            .I(counterZ0Z_0));
    Odrv4 I__2876 (
            .O(N__16054),
            .I(counterZ0Z_0));
    Odrv4 I__2875 (
            .O(N__16051),
            .I(counterZ0Z_0));
    Odrv12 I__2874 (
            .O(N__16048),
            .I(counterZ0Z_0));
    Odrv4 I__2873 (
            .O(N__16045),
            .I(counterZ0Z_0));
    LocalMux I__2872 (
            .O(N__16042),
            .I(counterZ0Z_0));
    Odrv4 I__2871 (
            .O(N__16037),
            .I(counterZ0Z_0));
    Odrv4 I__2870 (
            .O(N__16026),
            .I(counterZ0Z_0));
    Odrv12 I__2869 (
            .O(N__16023),
            .I(counterZ0Z_0));
    CascadeMux I__2868 (
            .O(N__15998),
            .I(N__15985));
    CascadeMux I__2867 (
            .O(N__15997),
            .I(N__15982));
    InMux I__2866 (
            .O(N__15996),
            .I(N__15971));
    InMux I__2865 (
            .O(N__15995),
            .I(N__15964));
    InMux I__2864 (
            .O(N__15994),
            .I(N__15964));
    InMux I__2863 (
            .O(N__15993),
            .I(N__15964));
    InMux I__2862 (
            .O(N__15992),
            .I(N__15959));
    InMux I__2861 (
            .O(N__15991),
            .I(N__15959));
    InMux I__2860 (
            .O(N__15990),
            .I(N__15952));
    InMux I__2859 (
            .O(N__15989),
            .I(N__15952));
    InMux I__2858 (
            .O(N__15988),
            .I(N__15952));
    InMux I__2857 (
            .O(N__15985),
            .I(N__15947));
    InMux I__2856 (
            .O(N__15982),
            .I(N__15947));
    InMux I__2855 (
            .O(N__15981),
            .I(N__15938));
    InMux I__2854 (
            .O(N__15980),
            .I(N__15938));
    InMux I__2853 (
            .O(N__15979),
            .I(N__15938));
    InMux I__2852 (
            .O(N__15978),
            .I(N__15938));
    InMux I__2851 (
            .O(N__15977),
            .I(N__15930));
    InMux I__2850 (
            .O(N__15976),
            .I(N__15930));
    CascadeMux I__2849 (
            .O(N__15975),
            .I(N__15927));
    CascadeMux I__2848 (
            .O(N__15974),
            .I(N__15924));
    LocalMux I__2847 (
            .O(N__15971),
            .I(N__15918));
    LocalMux I__2846 (
            .O(N__15964),
            .I(N__15918));
    LocalMux I__2845 (
            .O(N__15959),
            .I(N__15913));
    LocalMux I__2844 (
            .O(N__15952),
            .I(N__15913));
    LocalMux I__2843 (
            .O(N__15947),
            .I(N__15910));
    LocalMux I__2842 (
            .O(N__15938),
            .I(N__15907));
    InMux I__2841 (
            .O(N__15937),
            .I(N__15902));
    InMux I__2840 (
            .O(N__15936),
            .I(N__15902));
    InMux I__2839 (
            .O(N__15935),
            .I(N__15899));
    LocalMux I__2838 (
            .O(N__15930),
            .I(N__15896));
    InMux I__2837 (
            .O(N__15927),
            .I(N__15893));
    InMux I__2836 (
            .O(N__15924),
            .I(N__15890));
    InMux I__2835 (
            .O(N__15923),
            .I(N__15887));
    Span4Mux_s3_v I__2834 (
            .O(N__15918),
            .I(N__15876));
    Span4Mux_s3_v I__2833 (
            .O(N__15913),
            .I(N__15876));
    Span4Mux_s3_v I__2832 (
            .O(N__15910),
            .I(N__15876));
    Span4Mux_v I__2831 (
            .O(N__15907),
            .I(N__15876));
    LocalMux I__2830 (
            .O(N__15902),
            .I(N__15876));
    LocalMux I__2829 (
            .O(N__15899),
            .I(counterZ0Z_2));
    Odrv12 I__2828 (
            .O(N__15896),
            .I(counterZ0Z_2));
    LocalMux I__2827 (
            .O(N__15893),
            .I(counterZ0Z_2));
    LocalMux I__2826 (
            .O(N__15890),
            .I(counterZ0Z_2));
    LocalMux I__2825 (
            .O(N__15887),
            .I(counterZ0Z_2));
    Odrv4 I__2824 (
            .O(N__15876),
            .I(counterZ0Z_2));
    CascadeMux I__2823 (
            .O(N__15863),
            .I(N__15858));
    InMux I__2822 (
            .O(N__15862),
            .I(N__15851));
    CascadeMux I__2821 (
            .O(N__15861),
            .I(N__15848));
    InMux I__2820 (
            .O(N__15858),
            .I(N__15845));
    CascadeMux I__2819 (
            .O(N__15857),
            .I(N__15842));
    CascadeMux I__2818 (
            .O(N__15856),
            .I(N__15838));
    CascadeMux I__2817 (
            .O(N__15855),
            .I(N__15833));
    CascadeMux I__2816 (
            .O(N__15854),
            .I(N__15829));
    LocalMux I__2815 (
            .O(N__15851),
            .I(N__15826));
    InMux I__2814 (
            .O(N__15848),
            .I(N__15823));
    LocalMux I__2813 (
            .O(N__15845),
            .I(N__15807));
    InMux I__2812 (
            .O(N__15842),
            .I(N__15804));
    InMux I__2811 (
            .O(N__15841),
            .I(N__15797));
    InMux I__2810 (
            .O(N__15838),
            .I(N__15797));
    InMux I__2809 (
            .O(N__15837),
            .I(N__15797));
    InMux I__2808 (
            .O(N__15836),
            .I(N__15794));
    InMux I__2807 (
            .O(N__15833),
            .I(N__15787));
    InMux I__2806 (
            .O(N__15832),
            .I(N__15787));
    InMux I__2805 (
            .O(N__15829),
            .I(N__15787));
    Span4Mux_v I__2804 (
            .O(N__15826),
            .I(N__15782));
    LocalMux I__2803 (
            .O(N__15823),
            .I(N__15782));
    InMux I__2802 (
            .O(N__15822),
            .I(N__15773));
    InMux I__2801 (
            .O(N__15821),
            .I(N__15773));
    InMux I__2800 (
            .O(N__15820),
            .I(N__15773));
    InMux I__2799 (
            .O(N__15819),
            .I(N__15773));
    InMux I__2798 (
            .O(N__15818),
            .I(N__15770));
    InMux I__2797 (
            .O(N__15817),
            .I(N__15767));
    CascadeMux I__2796 (
            .O(N__15816),
            .I(N__15760));
    CascadeMux I__2795 (
            .O(N__15815),
            .I(N__15757));
    InMux I__2794 (
            .O(N__15814),
            .I(N__15751));
    CascadeMux I__2793 (
            .O(N__15813),
            .I(N__15746));
    CascadeMux I__2792 (
            .O(N__15812),
            .I(N__15743));
    CascadeMux I__2791 (
            .O(N__15811),
            .I(N__15736));
    InMux I__2790 (
            .O(N__15810),
            .I(N__15730));
    Span4Mux_v I__2789 (
            .O(N__15807),
            .I(N__15723));
    LocalMux I__2788 (
            .O(N__15804),
            .I(N__15723));
    LocalMux I__2787 (
            .O(N__15797),
            .I(N__15723));
    LocalMux I__2786 (
            .O(N__15794),
            .I(N__15715));
    LocalMux I__2785 (
            .O(N__15787),
            .I(N__15708));
    Span4Mux_s3_v I__2784 (
            .O(N__15782),
            .I(N__15708));
    LocalMux I__2783 (
            .O(N__15773),
            .I(N__15708));
    LocalMux I__2782 (
            .O(N__15770),
            .I(N__15703));
    LocalMux I__2781 (
            .O(N__15767),
            .I(N__15703));
    InMux I__2780 (
            .O(N__15766),
            .I(N__15694));
    InMux I__2779 (
            .O(N__15765),
            .I(N__15694));
    InMux I__2778 (
            .O(N__15764),
            .I(N__15694));
    InMux I__2777 (
            .O(N__15763),
            .I(N__15694));
    InMux I__2776 (
            .O(N__15760),
            .I(N__15689));
    InMux I__2775 (
            .O(N__15757),
            .I(N__15689));
    CascadeMux I__2774 (
            .O(N__15756),
            .I(N__15685));
    CascadeMux I__2773 (
            .O(N__15755),
            .I(N__15681));
    CascadeMux I__2772 (
            .O(N__15754),
            .I(N__15678));
    LocalMux I__2771 (
            .O(N__15751),
            .I(N__15675));
    InMux I__2770 (
            .O(N__15750),
            .I(N__15672));
    InMux I__2769 (
            .O(N__15749),
            .I(N__15665));
    InMux I__2768 (
            .O(N__15746),
            .I(N__15665));
    InMux I__2767 (
            .O(N__15743),
            .I(N__15665));
    InMux I__2766 (
            .O(N__15742),
            .I(N__15659));
    InMux I__2765 (
            .O(N__15741),
            .I(N__15659));
    InMux I__2764 (
            .O(N__15740),
            .I(N__15650));
    InMux I__2763 (
            .O(N__15739),
            .I(N__15650));
    InMux I__2762 (
            .O(N__15736),
            .I(N__15650));
    InMux I__2761 (
            .O(N__15735),
            .I(N__15650));
    CascadeMux I__2760 (
            .O(N__15734),
            .I(N__15647));
    CascadeMux I__2759 (
            .O(N__15733),
            .I(N__15644));
    LocalMux I__2758 (
            .O(N__15730),
            .I(N__15636));
    Span4Mux_s3_v I__2757 (
            .O(N__15723),
            .I(N__15636));
    InMux I__2756 (
            .O(N__15722),
            .I(N__15631));
    InMux I__2755 (
            .O(N__15721),
            .I(N__15631));
    InMux I__2754 (
            .O(N__15720),
            .I(N__15624));
    InMux I__2753 (
            .O(N__15719),
            .I(N__15624));
    InMux I__2752 (
            .O(N__15718),
            .I(N__15624));
    Span4Mux_h I__2751 (
            .O(N__15715),
            .I(N__15615));
    Span4Mux_v I__2750 (
            .O(N__15708),
            .I(N__15615));
    Span4Mux_v I__2749 (
            .O(N__15703),
            .I(N__15615));
    LocalMux I__2748 (
            .O(N__15694),
            .I(N__15615));
    LocalMux I__2747 (
            .O(N__15689),
            .I(N__15612));
    InMux I__2746 (
            .O(N__15688),
            .I(N__15607));
    InMux I__2745 (
            .O(N__15685),
            .I(N__15607));
    InMux I__2744 (
            .O(N__15684),
            .I(N__15604));
    InMux I__2743 (
            .O(N__15681),
            .I(N__15601));
    InMux I__2742 (
            .O(N__15678),
            .I(N__15598));
    Span4Mux_v I__2741 (
            .O(N__15675),
            .I(N__15591));
    LocalMux I__2740 (
            .O(N__15672),
            .I(N__15591));
    LocalMux I__2739 (
            .O(N__15665),
            .I(N__15591));
    InMux I__2738 (
            .O(N__15664),
            .I(N__15588));
    LocalMux I__2737 (
            .O(N__15659),
            .I(N__15583));
    LocalMux I__2736 (
            .O(N__15650),
            .I(N__15583));
    InMux I__2735 (
            .O(N__15647),
            .I(N__15572));
    InMux I__2734 (
            .O(N__15644),
            .I(N__15572));
    InMux I__2733 (
            .O(N__15643),
            .I(N__15572));
    InMux I__2732 (
            .O(N__15642),
            .I(N__15572));
    InMux I__2731 (
            .O(N__15641),
            .I(N__15572));
    Span4Mux_h I__2730 (
            .O(N__15636),
            .I(N__15567));
    LocalMux I__2729 (
            .O(N__15631),
            .I(N__15567));
    LocalMux I__2728 (
            .O(N__15624),
            .I(N__15562));
    Span4Mux_h I__2727 (
            .O(N__15615),
            .I(N__15562));
    Odrv4 I__2726 (
            .O(N__15612),
            .I(counterZ0Z_1));
    LocalMux I__2725 (
            .O(N__15607),
            .I(counterZ0Z_1));
    LocalMux I__2724 (
            .O(N__15604),
            .I(counterZ0Z_1));
    LocalMux I__2723 (
            .O(N__15601),
            .I(counterZ0Z_1));
    LocalMux I__2722 (
            .O(N__15598),
            .I(counterZ0Z_1));
    Odrv4 I__2721 (
            .O(N__15591),
            .I(counterZ0Z_1));
    LocalMux I__2720 (
            .O(N__15588),
            .I(counterZ0Z_1));
    Odrv4 I__2719 (
            .O(N__15583),
            .I(counterZ0Z_1));
    LocalMux I__2718 (
            .O(N__15572),
            .I(counterZ0Z_1));
    Odrv4 I__2717 (
            .O(N__15567),
            .I(counterZ0Z_1));
    Odrv4 I__2716 (
            .O(N__15562),
            .I(counterZ0Z_1));
    InMux I__2715 (
            .O(N__15539),
            .I(N__15536));
    LocalMux I__2714 (
            .O(N__15536),
            .I(un1_sclk17_4_1));
    InMux I__2713 (
            .O(N__15533),
            .I(N__15529));
    InMux I__2712 (
            .O(N__15532),
            .I(N__15526));
    LocalMux I__2711 (
            .O(N__15529),
            .I(N_1505));
    LocalMux I__2710 (
            .O(N__15526),
            .I(N_1505));
    InMux I__2709 (
            .O(N__15521),
            .I(N__15516));
    InMux I__2708 (
            .O(N__15520),
            .I(N__15513));
    CascadeMux I__2707 (
            .O(N__15519),
            .I(N__15509));
    LocalMux I__2706 (
            .O(N__15516),
            .I(N__15506));
    LocalMux I__2705 (
            .O(N__15513),
            .I(N__15503));
    InMux I__2704 (
            .O(N__15512),
            .I(N__15498));
    InMux I__2703 (
            .O(N__15509),
            .I(N__15498));
    Span4Mux_h I__2702 (
            .O(N__15506),
            .I(N__15495));
    Span4Mux_h I__2701 (
            .O(N__15503),
            .I(N__15492));
    LocalMux I__2700 (
            .O(N__15498),
            .I(N_1509));
    Odrv4 I__2699 (
            .O(N__15495),
            .I(N_1509));
    Odrv4 I__2698 (
            .O(N__15492),
            .I(N_1509));
    CascadeMux I__2697 (
            .O(N__15485),
            .I(N__15482));
    InMux I__2696 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__2695 (
            .O(N__15479),
            .I(N__15476));
    Odrv4 I__2694 (
            .O(N__15476),
            .I(un42_cry_2_c_RNOZ0));
    CascadeMux I__2693 (
            .O(N__15473),
            .I(un1_sclk17_6_1_cascade_));
    CascadeMux I__2692 (
            .O(N__15470),
            .I(un1_sclk17_3_1_cascade_));
    InMux I__2691 (
            .O(N__15467),
            .I(N__15464));
    LocalMux I__2690 (
            .O(N__15464),
            .I(N__15461));
    Odrv12 I__2689 (
            .O(N__15461),
            .I(ScreenBuffer_0_0_1_sqmuxa_0));
    InMux I__2688 (
            .O(N__15458),
            .I(N__15454));
    InMux I__2687 (
            .O(N__15457),
            .I(N__15451));
    LocalMux I__2686 (
            .O(N__15454),
            .I(slaveselect_RNILOQCZ0Z2));
    LocalMux I__2685 (
            .O(N__15451),
            .I(slaveselect_RNILOQCZ0Z2));
    CascadeMux I__2684 (
            .O(N__15446),
            .I(un1_sclk17_8_0_0_cascade_));
    CascadeMux I__2683 (
            .O(N__15443),
            .I(N__15440));
    InMux I__2682 (
            .O(N__15440),
            .I(N__15437));
    LocalMux I__2681 (
            .O(N__15437),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3));
    InMux I__2680 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__2679 (
            .O(N__15431),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5));
    InMux I__2678 (
            .O(N__15428),
            .I(N__15425));
    LocalMux I__2677 (
            .O(N__15425),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO));
    InMux I__2676 (
            .O(N__15422),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4));
    InMux I__2675 (
            .O(N__15419),
            .I(N__15413));
    InMux I__2674 (
            .O(N__15418),
            .I(N__15413));
    LocalMux I__2673 (
            .O(N__15413),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO));
    CascadeMux I__2672 (
            .O(N__15410),
            .I(N__15406));
    InMux I__2671 (
            .O(N__15409),
            .I(N__15398));
    InMux I__2670 (
            .O(N__15406),
            .I(N__15398));
    InMux I__2669 (
            .O(N__15405),
            .I(N__15398));
    LocalMux I__2668 (
            .O(N__15398),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803));
    InMux I__2667 (
            .O(N__15395),
            .I(N__15392));
    LocalMux I__2666 (
            .O(N__15392),
            .I(N__15386));
    InMux I__2665 (
            .O(N__15391),
            .I(N__15381));
    InMux I__2664 (
            .O(N__15390),
            .I(N__15381));
    CascadeMux I__2663 (
            .O(N__15389),
            .I(N__15376));
    Span4Mux_h I__2662 (
            .O(N__15386),
            .I(N__15372));
    LocalMux I__2661 (
            .O(N__15381),
            .I(N__15369));
    InMux I__2660 (
            .O(N__15380),
            .I(N__15366));
    InMux I__2659 (
            .O(N__15379),
            .I(N__15363));
    InMux I__2658 (
            .O(N__15376),
            .I(N__15358));
    InMux I__2657 (
            .O(N__15375),
            .I(N__15358));
    Span4Mux_v I__2656 (
            .O(N__15372),
            .I(N__15353));
    Span4Mux_h I__2655 (
            .O(N__15369),
            .I(N__15353));
    LocalMux I__2654 (
            .O(N__15366),
            .I(voltage_2Z0Z_0));
    LocalMux I__2653 (
            .O(N__15363),
            .I(voltage_2Z0Z_0));
    LocalMux I__2652 (
            .O(N__15358),
            .I(voltage_2Z0Z_0));
    Odrv4 I__2651 (
            .O(N__15353),
            .I(voltage_2Z0Z_0));
    InMux I__2650 (
            .O(N__15344),
            .I(N__15340));
    InMux I__2649 (
            .O(N__15343),
            .I(N__15336));
    LocalMux I__2648 (
            .O(N__15340),
            .I(N__15333));
    InMux I__2647 (
            .O(N__15339),
            .I(N__15330));
    LocalMux I__2646 (
            .O(N__15336),
            .I(N__15325));
    Span4Mux_v I__2645 (
            .O(N__15333),
            .I(N__15322));
    LocalMux I__2644 (
            .O(N__15330),
            .I(N__15319));
    InMux I__2643 (
            .O(N__15329),
            .I(N__15314));
    InMux I__2642 (
            .O(N__15328),
            .I(N__15314));
    Odrv12 I__2641 (
            .O(N__15325),
            .I(voltage_1Z0Z_0));
    Odrv4 I__2640 (
            .O(N__15322),
            .I(voltage_1Z0Z_0));
    Odrv4 I__2639 (
            .O(N__15319),
            .I(voltage_1Z0Z_0));
    LocalMux I__2638 (
            .O(N__15314),
            .I(voltage_1Z0Z_0));
    CascadeMux I__2637 (
            .O(N__15305),
            .I(N__15302));
    InMux I__2636 (
            .O(N__15302),
            .I(N__15298));
    InMux I__2635 (
            .O(N__15301),
            .I(N__15295));
    LocalMux I__2634 (
            .O(N__15298),
            .I(N__15290));
    LocalMux I__2633 (
            .O(N__15295),
            .I(N__15287));
    InMux I__2632 (
            .O(N__15294),
            .I(N__15283));
    InMux I__2631 (
            .O(N__15293),
            .I(N__15280));
    Span4Mux_v I__2630 (
            .O(N__15290),
            .I(N__15275));
    Span4Mux_s1_h I__2629 (
            .O(N__15287),
            .I(N__15275));
    InMux I__2628 (
            .O(N__15286),
            .I(N__15272));
    LocalMux I__2627 (
            .O(N__15283),
            .I(voltage_2Z0Z_2));
    LocalMux I__2626 (
            .O(N__15280),
            .I(voltage_2Z0Z_2));
    Odrv4 I__2625 (
            .O(N__15275),
            .I(voltage_2Z0Z_2));
    LocalMux I__2624 (
            .O(N__15272),
            .I(voltage_2Z0Z_2));
    InMux I__2623 (
            .O(N__15263),
            .I(N__15258));
    CascadeMux I__2622 (
            .O(N__15262),
            .I(N__15255));
    InMux I__2621 (
            .O(N__15261),
            .I(N__15252));
    LocalMux I__2620 (
            .O(N__15258),
            .I(N__15249));
    InMux I__2619 (
            .O(N__15255),
            .I(N__15246));
    LocalMux I__2618 (
            .O(N__15252),
            .I(N__15242));
    Span4Mux_v I__2617 (
            .O(N__15249),
            .I(N__15239));
    LocalMux I__2616 (
            .O(N__15246),
            .I(N__15236));
    InMux I__2615 (
            .O(N__15245),
            .I(N__15233));
    Odrv12 I__2614 (
            .O(N__15242),
            .I(voltage_1Z0Z_2));
    Odrv4 I__2613 (
            .O(N__15239),
            .I(voltage_1Z0Z_2));
    Odrv12 I__2612 (
            .O(N__15236),
            .I(voltage_1Z0Z_2));
    LocalMux I__2611 (
            .O(N__15233),
            .I(voltage_1Z0Z_2));
    InMux I__2610 (
            .O(N__15224),
            .I(N__15220));
    InMux I__2609 (
            .O(N__15223),
            .I(N__15216));
    LocalMux I__2608 (
            .O(N__15220),
            .I(N__15213));
    CascadeMux I__2607 (
            .O(N__15219),
            .I(N__15210));
    LocalMux I__2606 (
            .O(N__15216),
            .I(N__15206));
    Span4Mux_h I__2605 (
            .O(N__15213),
            .I(N__15202));
    InMux I__2604 (
            .O(N__15210),
            .I(N__15197));
    InMux I__2603 (
            .O(N__15209),
            .I(N__15197));
    Span4Mux_v I__2602 (
            .O(N__15206),
            .I(N__15194));
    InMux I__2601 (
            .O(N__15205),
            .I(N__15191));
    Span4Mux_v I__2600 (
            .O(N__15202),
            .I(N__15188));
    LocalMux I__2599 (
            .O(N__15197),
            .I(N__15185));
    Odrv4 I__2598 (
            .O(N__15194),
            .I(voltage_2Z0Z_3));
    LocalMux I__2597 (
            .O(N__15191),
            .I(voltage_2Z0Z_3));
    Odrv4 I__2596 (
            .O(N__15188),
            .I(voltage_2Z0Z_3));
    Odrv4 I__2595 (
            .O(N__15185),
            .I(voltage_2Z0Z_3));
    InMux I__2594 (
            .O(N__15176),
            .I(N__15172));
    InMux I__2593 (
            .O(N__15175),
            .I(N__15169));
    LocalMux I__2592 (
            .O(N__15172),
            .I(N__15164));
    LocalMux I__2591 (
            .O(N__15169),
            .I(N__15164));
    Span4Mux_v I__2590 (
            .O(N__15164),
            .I(N__15159));
    InMux I__2589 (
            .O(N__15163),
            .I(N__15156));
    InMux I__2588 (
            .O(N__15162),
            .I(N__15153));
    Odrv4 I__2587 (
            .O(N__15159),
            .I(voltage_1Z0Z_3));
    LocalMux I__2586 (
            .O(N__15156),
            .I(voltage_1Z0Z_3));
    LocalMux I__2585 (
            .O(N__15153),
            .I(voltage_1Z0Z_3));
    InMux I__2584 (
            .O(N__15146),
            .I(N__15143));
    LocalMux I__2583 (
            .O(N__15143),
            .I(N__15139));
    InMux I__2582 (
            .O(N__15142),
            .I(N__15136));
    Span4Mux_s2_h I__2581 (
            .O(N__15139),
            .I(N__15130));
    LocalMux I__2580 (
            .O(N__15136),
            .I(N__15130));
    InMux I__2579 (
            .O(N__15135),
            .I(N__15124));
    Span4Mux_v I__2578 (
            .O(N__15130),
            .I(N__15121));
    InMux I__2577 (
            .O(N__15129),
            .I(N__15116));
    InMux I__2576 (
            .O(N__15128),
            .I(N__15116));
    InMux I__2575 (
            .O(N__15127),
            .I(N__15113));
    LocalMux I__2574 (
            .O(N__15124),
            .I(voltage_2Z0Z_1));
    Odrv4 I__2573 (
            .O(N__15121),
            .I(voltage_2Z0Z_1));
    LocalMux I__2572 (
            .O(N__15116),
            .I(voltage_2Z0Z_1));
    LocalMux I__2571 (
            .O(N__15113),
            .I(voltage_2Z0Z_1));
    InMux I__2570 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__2569 (
            .O(N__15101),
            .I(N__15096));
    InMux I__2568 (
            .O(N__15100),
            .I(N__15093));
    InMux I__2567 (
            .O(N__15099),
            .I(N__15090));
    Span4Mux_v I__2566 (
            .O(N__15096),
            .I(N__15087));
    LocalMux I__2565 (
            .O(N__15093),
            .I(N__15083));
    LocalMux I__2564 (
            .O(N__15090),
            .I(N__15078));
    Span4Mux_s2_h I__2563 (
            .O(N__15087),
            .I(N__15078));
    InMux I__2562 (
            .O(N__15086),
            .I(N__15075));
    Odrv4 I__2561 (
            .O(N__15083),
            .I(voltage_1Z0Z_1));
    Odrv4 I__2560 (
            .O(N__15078),
            .I(voltage_1Z0Z_1));
    LocalMux I__2559 (
            .O(N__15075),
            .I(voltage_1Z0Z_1));
    CEMux I__2558 (
            .O(N__15068),
            .I(N__15065));
    LocalMux I__2557 (
            .O(N__15065),
            .I(N__15062));
    Span4Mux_h I__2556 (
            .O(N__15062),
            .I(N__15059));
    Odrv4 I__2555 (
            .O(N__15059),
            .I(un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0));
    InMux I__2554 (
            .O(N__15056),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1));
    InMux I__2553 (
            .O(N__15053),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2));
    InMux I__2552 (
            .O(N__15050),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3));
    InMux I__2551 (
            .O(N__15047),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4));
    CascadeMux I__2550 (
            .O(N__15044),
            .I(N__15041));
    InMux I__2549 (
            .O(N__15041),
            .I(N__15038));
    LocalMux I__2548 (
            .O(N__15038),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_i));
    InMux I__2547 (
            .O(N__15035),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1));
    InMux I__2546 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__2545 (
            .O(N__15029),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3));
    InMux I__2544 (
            .O(N__15026),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2));
    InMux I__2543 (
            .O(N__15023),
            .I(N__15020));
    LocalMux I__2542 (
            .O(N__15020),
            .I(N__15017));
    Odrv4 I__2541 (
            .O(N__15017),
            .I(un13_beamy_0));
    InMux I__2540 (
            .O(N__15014),
            .I(N__15011));
    LocalMux I__2539 (
            .O(N__15011),
            .I(N__15008));
    Odrv4 I__2538 (
            .O(N__15008),
            .I(chessboardpixel_un174_pixel));
    CascadeMux I__2537 (
            .O(N__15005),
            .I(un4_row_cascade_));
    InMux I__2536 (
            .O(N__15002),
            .I(N__14999));
    LocalMux I__2535 (
            .O(N__14999),
            .I(N__14995));
    InMux I__2534 (
            .O(N__14998),
            .I(N__14992));
    Span4Mux_v I__2533 (
            .O(N__14995),
            .I(N__14984));
    LocalMux I__2532 (
            .O(N__14992),
            .I(N__14984));
    InMux I__2531 (
            .O(N__14991),
            .I(N__14980));
    InMux I__2530 (
            .O(N__14990),
            .I(N__14977));
    InMux I__2529 (
            .O(N__14989),
            .I(N__14974));
    Span4Mux_v I__2528 (
            .O(N__14984),
            .I(N__14969));
    InMux I__2527 (
            .O(N__14983),
            .I(N__14966));
    LocalMux I__2526 (
            .O(N__14980),
            .I(N__14963));
    LocalMux I__2525 (
            .O(N__14977),
            .I(N__14958));
    LocalMux I__2524 (
            .O(N__14974),
            .I(N__14958));
    InMux I__2523 (
            .O(N__14973),
            .I(N__14955));
    InMux I__2522 (
            .O(N__14972),
            .I(N__14952));
    Sp12to4 I__2521 (
            .O(N__14969),
            .I(N__14947));
    LocalMux I__2520 (
            .O(N__14966),
            .I(N__14947));
    Span4Mux_v I__2519 (
            .O(N__14963),
            .I(N__14942));
    Span4Mux_v I__2518 (
            .O(N__14958),
            .I(N__14942));
    LocalMux I__2517 (
            .O(N__14955),
            .I(N__14939));
    LocalMux I__2516 (
            .O(N__14952),
            .I(beamYZ0Z_9));
    Odrv12 I__2515 (
            .O(N__14947),
            .I(beamYZ0Z_9));
    Odrv4 I__2514 (
            .O(N__14942),
            .I(beamYZ0Z_9));
    Odrv4 I__2513 (
            .O(N__14939),
            .I(beamYZ0Z_9));
    CascadeMux I__2512 (
            .O(N__14930),
            .I(N__14926));
    CascadeMux I__2511 (
            .O(N__14929),
            .I(N__14922));
    InMux I__2510 (
            .O(N__14926),
            .I(N__14917));
    InMux I__2509 (
            .O(N__14925),
            .I(N__14914));
    InMux I__2508 (
            .O(N__14922),
            .I(N__14911));
    InMux I__2507 (
            .O(N__14921),
            .I(N__14908));
    InMux I__2506 (
            .O(N__14920),
            .I(N__14905));
    LocalMux I__2505 (
            .O(N__14917),
            .I(N__14898));
    LocalMux I__2504 (
            .O(N__14914),
            .I(N__14898));
    LocalMux I__2503 (
            .O(N__14911),
            .I(N__14898));
    LocalMux I__2502 (
            .O(N__14908),
            .I(N__14893));
    LocalMux I__2501 (
            .O(N__14905),
            .I(N__14893));
    Span4Mux_v I__2500 (
            .O(N__14898),
            .I(N__14884));
    Span4Mux_v I__2499 (
            .O(N__14893),
            .I(N__14884));
    InMux I__2498 (
            .O(N__14892),
            .I(N__14881));
    InMux I__2497 (
            .O(N__14891),
            .I(N__14878));
    CascadeMux I__2496 (
            .O(N__14890),
            .I(N__14874));
    InMux I__2495 (
            .O(N__14889),
            .I(N__14871));
    Sp12to4 I__2494 (
            .O(N__14884),
            .I(N__14866));
    LocalMux I__2493 (
            .O(N__14881),
            .I(N__14866));
    LocalMux I__2492 (
            .O(N__14878),
            .I(N__14863));
    InMux I__2491 (
            .O(N__14877),
            .I(N__14860));
    InMux I__2490 (
            .O(N__14874),
            .I(N__14857));
    LocalMux I__2489 (
            .O(N__14871),
            .I(beamYZ0Z_8));
    Odrv12 I__2488 (
            .O(N__14866),
            .I(beamYZ0Z_8));
    Odrv4 I__2487 (
            .O(N__14863),
            .I(beamYZ0Z_8));
    LocalMux I__2486 (
            .O(N__14860),
            .I(beamYZ0Z_8));
    LocalMux I__2485 (
            .O(N__14857),
            .I(beamYZ0Z_8));
    CascadeMux I__2484 (
            .O(N__14846),
            .I(N__14842));
    CascadeMux I__2483 (
            .O(N__14845),
            .I(N__14839));
    InMux I__2482 (
            .O(N__14842),
            .I(N__14834));
    InMux I__2481 (
            .O(N__14839),
            .I(N__14831));
    InMux I__2480 (
            .O(N__14838),
            .I(N__14828));
    InMux I__2479 (
            .O(N__14837),
            .I(N__14825));
    LocalMux I__2478 (
            .O(N__14834),
            .I(N__14821));
    LocalMux I__2477 (
            .O(N__14831),
            .I(N__14818));
    LocalMux I__2476 (
            .O(N__14828),
            .I(N__14813));
    LocalMux I__2475 (
            .O(N__14825),
            .I(N__14813));
    InMux I__2474 (
            .O(N__14824),
            .I(N__14806));
    Span4Mux_h I__2473 (
            .O(N__14821),
            .I(N__14803));
    Span4Mux_h I__2472 (
            .O(N__14818),
            .I(N__14800));
    Span4Mux_v I__2471 (
            .O(N__14813),
            .I(N__14797));
    InMux I__2470 (
            .O(N__14812),
            .I(N__14794));
    InMux I__2469 (
            .O(N__14811),
            .I(N__14791));
    CascadeMux I__2468 (
            .O(N__14810),
            .I(N__14786));
    InMux I__2467 (
            .O(N__14809),
            .I(N__14777));
    LocalMux I__2466 (
            .O(N__14806),
            .I(N__14774));
    Span4Mux_h I__2465 (
            .O(N__14803),
            .I(N__14771));
    Span4Mux_h I__2464 (
            .O(N__14800),
            .I(N__14768));
    Sp12to4 I__2463 (
            .O(N__14797),
            .I(N__14761));
    LocalMux I__2462 (
            .O(N__14794),
            .I(N__14761));
    LocalMux I__2461 (
            .O(N__14791),
            .I(N__14761));
    InMux I__2460 (
            .O(N__14790),
            .I(N__14756));
    InMux I__2459 (
            .O(N__14789),
            .I(N__14756));
    InMux I__2458 (
            .O(N__14786),
            .I(N__14751));
    InMux I__2457 (
            .O(N__14785),
            .I(N__14751));
    InMux I__2456 (
            .O(N__14784),
            .I(N__14746));
    InMux I__2455 (
            .O(N__14783),
            .I(N__14746));
    InMux I__2454 (
            .O(N__14782),
            .I(N__14739));
    InMux I__2453 (
            .O(N__14781),
            .I(N__14739));
    InMux I__2452 (
            .O(N__14780),
            .I(N__14739));
    LocalMux I__2451 (
            .O(N__14777),
            .I(beamYZ0Z_7));
    Odrv4 I__2450 (
            .O(N__14774),
            .I(beamYZ0Z_7));
    Odrv4 I__2449 (
            .O(N__14771),
            .I(beamYZ0Z_7));
    Odrv4 I__2448 (
            .O(N__14768),
            .I(beamYZ0Z_7));
    Odrv12 I__2447 (
            .O(N__14761),
            .I(beamYZ0Z_7));
    LocalMux I__2446 (
            .O(N__14756),
            .I(beamYZ0Z_7));
    LocalMux I__2445 (
            .O(N__14751),
            .I(beamYZ0Z_7));
    LocalMux I__2444 (
            .O(N__14746),
            .I(beamYZ0Z_7));
    LocalMux I__2443 (
            .O(N__14739),
            .I(beamYZ0Z_7));
    InMux I__2442 (
            .O(N__14720),
            .I(N__14717));
    LocalMux I__2441 (
            .O(N__14717),
            .I(un4_beamylt8_0));
    InMux I__2440 (
            .O(N__14714),
            .I(N__14711));
    LocalMux I__2439 (
            .O(N__14711),
            .I(un4_beamy_0));
    InMux I__2438 (
            .O(N__14708),
            .I(N__14705));
    LocalMux I__2437 (
            .O(N__14705),
            .I(un113_pixel_4_0_15__un8_beamylto9Z0Z_1));
    CascadeMux I__2436 (
            .O(N__14702),
            .I(N__14697));
    CascadeMux I__2435 (
            .O(N__14701),
            .I(N__14691));
    InMux I__2434 (
            .O(N__14700),
            .I(N__14684));
    InMux I__2433 (
            .O(N__14697),
            .I(N__14681));
    InMux I__2432 (
            .O(N__14696),
            .I(N__14678));
    InMux I__2431 (
            .O(N__14695),
            .I(N__14675));
    InMux I__2430 (
            .O(N__14694),
            .I(N__14672));
    InMux I__2429 (
            .O(N__14691),
            .I(N__14669));
    InMux I__2428 (
            .O(N__14690),
            .I(N__14662));
    InMux I__2427 (
            .O(N__14689),
            .I(N__14662));
    InMux I__2426 (
            .O(N__14688),
            .I(N__14662));
    InMux I__2425 (
            .O(N__14687),
            .I(N__14654));
    LocalMux I__2424 (
            .O(N__14684),
            .I(N__14651));
    LocalMux I__2423 (
            .O(N__14681),
            .I(N__14648));
    LocalMux I__2422 (
            .O(N__14678),
            .I(N__14645));
    LocalMux I__2421 (
            .O(N__14675),
            .I(N__14640));
    LocalMux I__2420 (
            .O(N__14672),
            .I(N__14640));
    LocalMux I__2419 (
            .O(N__14669),
            .I(N__14637));
    LocalMux I__2418 (
            .O(N__14662),
            .I(N__14634));
    InMux I__2417 (
            .O(N__14661),
            .I(N__14631));
    CascadeMux I__2416 (
            .O(N__14660),
            .I(N__14627));
    CascadeMux I__2415 (
            .O(N__14659),
            .I(N__14624));
    CascadeMux I__2414 (
            .O(N__14658),
            .I(N__14618));
    InMux I__2413 (
            .O(N__14657),
            .I(N__14614));
    LocalMux I__2412 (
            .O(N__14654),
            .I(N__14611));
    Span12Mux_s5_v I__2411 (
            .O(N__14651),
            .I(N__14606));
    Span12Mux_s10_v I__2410 (
            .O(N__14648),
            .I(N__14606));
    Span4Mux_v I__2409 (
            .O(N__14645),
            .I(N__14601));
    Span4Mux_v I__2408 (
            .O(N__14640),
            .I(N__14601));
    Span4Mux_v I__2407 (
            .O(N__14637),
            .I(N__14596));
    Span4Mux_v I__2406 (
            .O(N__14634),
            .I(N__14596));
    LocalMux I__2405 (
            .O(N__14631),
            .I(N__14593));
    InMux I__2404 (
            .O(N__14630),
            .I(N__14588));
    InMux I__2403 (
            .O(N__14627),
            .I(N__14588));
    InMux I__2402 (
            .O(N__14624),
            .I(N__14585));
    InMux I__2401 (
            .O(N__14623),
            .I(N__14580));
    InMux I__2400 (
            .O(N__14622),
            .I(N__14580));
    InMux I__2399 (
            .O(N__14621),
            .I(N__14573));
    InMux I__2398 (
            .O(N__14618),
            .I(N__14573));
    InMux I__2397 (
            .O(N__14617),
            .I(N__14573));
    LocalMux I__2396 (
            .O(N__14614),
            .I(beamYZ0Z_4));
    Odrv4 I__2395 (
            .O(N__14611),
            .I(beamYZ0Z_4));
    Odrv12 I__2394 (
            .O(N__14606),
            .I(beamYZ0Z_4));
    Odrv4 I__2393 (
            .O(N__14601),
            .I(beamYZ0Z_4));
    Odrv4 I__2392 (
            .O(N__14596),
            .I(beamYZ0Z_4));
    Odrv4 I__2391 (
            .O(N__14593),
            .I(beamYZ0Z_4));
    LocalMux I__2390 (
            .O(N__14588),
            .I(beamYZ0Z_4));
    LocalMux I__2389 (
            .O(N__14585),
            .I(beamYZ0Z_4));
    LocalMux I__2388 (
            .O(N__14580),
            .I(beamYZ0Z_4));
    LocalMux I__2387 (
            .O(N__14573),
            .I(beamYZ0Z_4));
    CascadeMux I__2386 (
            .O(N__14552),
            .I(N__14549));
    InMux I__2385 (
            .O(N__14549),
            .I(N__14546));
    LocalMux I__2384 (
            .O(N__14546),
            .I(N__14543));
    Odrv4 I__2383 (
            .O(N__14543),
            .I(un8_beamy));
    CascadeMux I__2382 (
            .O(N__14540),
            .I(N__14537));
    InMux I__2381 (
            .O(N__14537),
            .I(N__14534));
    LocalMux I__2380 (
            .O(N__14534),
            .I(N_6_i));
    CascadeMux I__2379 (
            .O(N__14531),
            .I(N_6_i_cascade_));
    InMux I__2378 (
            .O(N__14528),
            .I(N__14525));
    LocalMux I__2377 (
            .O(N__14525),
            .I(N__14522));
    Span4Mux_h I__2376 (
            .O(N__14522),
            .I(N__14514));
    InMux I__2375 (
            .O(N__14521),
            .I(N__14511));
    InMux I__2374 (
            .O(N__14520),
            .I(N__14502));
    InMux I__2373 (
            .O(N__14519),
            .I(N__14502));
    InMux I__2372 (
            .O(N__14518),
            .I(N__14502));
    InMux I__2371 (
            .O(N__14517),
            .I(N__14502));
    Odrv4 I__2370 (
            .O(N__14514),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3));
    LocalMux I__2369 (
            .O(N__14511),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3));
    LocalMux I__2368 (
            .O(N__14502),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3));
    InMux I__2367 (
            .O(N__14495),
            .I(N__14491));
    InMux I__2366 (
            .O(N__14494),
            .I(N__14488));
    LocalMux I__2365 (
            .O(N__14491),
            .I(N__14482));
    LocalMux I__2364 (
            .O(N__14488),
            .I(N__14482));
    CascadeMux I__2363 (
            .O(N__14487),
            .I(N__14473));
    Span4Mux_v I__2362 (
            .O(N__14482),
            .I(N__14466));
    InMux I__2361 (
            .O(N__14481),
            .I(N__14459));
    InMux I__2360 (
            .O(N__14480),
            .I(N__14459));
    InMux I__2359 (
            .O(N__14479),
            .I(N__14459));
    InMux I__2358 (
            .O(N__14478),
            .I(N__14454));
    InMux I__2357 (
            .O(N__14477),
            .I(N__14454));
    InMux I__2356 (
            .O(N__14476),
            .I(N__14451));
    InMux I__2355 (
            .O(N__14473),
            .I(N__14442));
    InMux I__2354 (
            .O(N__14472),
            .I(N__14442));
    InMux I__2353 (
            .O(N__14471),
            .I(N__14442));
    InMux I__2352 (
            .O(N__14470),
            .I(N__14442));
    InMux I__2351 (
            .O(N__14469),
            .I(N__14437));
    Sp12to4 I__2350 (
            .O(N__14466),
            .I(N__14430));
    LocalMux I__2349 (
            .O(N__14459),
            .I(N__14430));
    LocalMux I__2348 (
            .O(N__14454),
            .I(N__14430));
    LocalMux I__2347 (
            .O(N__14451),
            .I(N__14425));
    LocalMux I__2346 (
            .O(N__14442),
            .I(N__14425));
    InMux I__2345 (
            .O(N__14441),
            .I(N__14422));
    InMux I__2344 (
            .O(N__14440),
            .I(N__14414));
    LocalMux I__2343 (
            .O(N__14437),
            .I(N__14411));
    Span12Mux_s11_h I__2342 (
            .O(N__14430),
            .I(N__14408));
    Span4Mux_v I__2341 (
            .O(N__14425),
            .I(N__14403));
    LocalMux I__2340 (
            .O(N__14422),
            .I(N__14403));
    InMux I__2339 (
            .O(N__14421),
            .I(N__14400));
    InMux I__2338 (
            .O(N__14420),
            .I(N__14395));
    InMux I__2337 (
            .O(N__14419),
            .I(N__14395));
    InMux I__2336 (
            .O(N__14418),
            .I(N__14392));
    InMux I__2335 (
            .O(N__14417),
            .I(N__14389));
    LocalMux I__2334 (
            .O(N__14414),
            .I(beamYZ0Z_3));
    Odrv4 I__2333 (
            .O(N__14411),
            .I(beamYZ0Z_3));
    Odrv12 I__2332 (
            .O(N__14408),
            .I(beamYZ0Z_3));
    Odrv4 I__2331 (
            .O(N__14403),
            .I(beamYZ0Z_3));
    LocalMux I__2330 (
            .O(N__14400),
            .I(beamYZ0Z_3));
    LocalMux I__2329 (
            .O(N__14395),
            .I(beamYZ0Z_3));
    LocalMux I__2328 (
            .O(N__14392),
            .I(beamYZ0Z_3));
    LocalMux I__2327 (
            .O(N__14389),
            .I(beamYZ0Z_3));
    InMux I__2326 (
            .O(N__14372),
            .I(N__14367));
    InMux I__2325 (
            .O(N__14371),
            .I(N__14364));
    InMux I__2324 (
            .O(N__14370),
            .I(N__14361));
    LocalMux I__2323 (
            .O(N__14367),
            .I(un4_beamylt6));
    LocalMux I__2322 (
            .O(N__14364),
            .I(un4_beamylt6));
    LocalMux I__2321 (
            .O(N__14361),
            .I(un4_beamylt6));
    InMux I__2320 (
            .O(N__14354),
            .I(N__14351));
    LocalMux I__2319 (
            .O(N__14351),
            .I(N__14348));
    Odrv4 I__2318 (
            .O(N__14348),
            .I(if_m1_ns));
    CascadeMux I__2317 (
            .O(N__14345),
            .I(if_m2_2_cascade_));
    InMux I__2316 (
            .O(N__14342),
            .I(N__14339));
    LocalMux I__2315 (
            .O(N__14339),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5_0));
    InMux I__2314 (
            .O(N__14336),
            .I(N__14330));
    InMux I__2313 (
            .O(N__14335),
            .I(N__14330));
    LocalMux I__2312 (
            .O(N__14330),
            .I(un18_beamylt4));
    InMux I__2311 (
            .O(N__14327),
            .I(N__14324));
    LocalMux I__2310 (
            .O(N__14324),
            .I(un113_pixel_4_0_15__un4_rowZ0Z_2));
    InMux I__2309 (
            .O(N__14321),
            .I(N__14318));
    LocalMux I__2308 (
            .O(N__14318),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    CascadeMux I__2307 (
            .O(N__14315),
            .I(N__14312));
    InMux I__2306 (
            .O(N__14312),
            .I(N__14307));
    CascadeMux I__2305 (
            .O(N__14311),
            .I(N__14304));
    CascadeMux I__2304 (
            .O(N__14310),
            .I(N__14300));
    LocalMux I__2303 (
            .O(N__14307),
            .I(N__14294));
    InMux I__2302 (
            .O(N__14304),
            .I(N__14289));
    InMux I__2301 (
            .O(N__14303),
            .I(N__14289));
    InMux I__2300 (
            .O(N__14300),
            .I(N__14284));
    InMux I__2299 (
            .O(N__14299),
            .I(N__14284));
    CascadeMux I__2298 (
            .O(N__14298),
            .I(N__14281));
    CascadeMux I__2297 (
            .O(N__14297),
            .I(N__14278));
    Span4Mux_h I__2296 (
            .O(N__14294),
            .I(N__14273));
    LocalMux I__2295 (
            .O(N__14289),
            .I(N__14273));
    LocalMux I__2294 (
            .O(N__14284),
            .I(N__14270));
    InMux I__2293 (
            .O(N__14281),
            .I(N__14265));
    InMux I__2292 (
            .O(N__14278),
            .I(N__14265));
    Span4Mux_v I__2291 (
            .O(N__14273),
            .I(N__14260));
    Span4Mux_h I__2290 (
            .O(N__14270),
            .I(N__14260));
    LocalMux I__2289 (
            .O(N__14265),
            .I(N__14257));
    Span4Mux_h I__2288 (
            .O(N__14260),
            .I(N__14254));
    Odrv4 I__2287 (
            .O(N__14257),
            .I(r_N_6));
    Odrv4 I__2286 (
            .O(N__14254),
            .I(r_N_6));
    InMux I__2285 (
            .O(N__14249),
            .I(N__14246));
    LocalMux I__2284 (
            .O(N__14246),
            .I(un113_pixel_4_0_15__un3_beamxZ0Z_7));
    CascadeMux I__2283 (
            .O(N__14243),
            .I(un1_beamxlt10_0_cascade_));
    IoInMux I__2282 (
            .O(N__14240),
            .I(N__14237));
    LocalMux I__2281 (
            .O(N__14237),
            .I(N__14234));
    IoSpan4Mux I__2280 (
            .O(N__14234),
            .I(N__14231));
    Span4Mux_s3_v I__2279 (
            .O(N__14231),
            .I(N__14228));
    Odrv4 I__2278 (
            .O(N__14228),
            .I(HSync_c));
    InMux I__2277 (
            .O(N__14225),
            .I(N__14222));
    LocalMux I__2276 (
            .O(N__14222),
            .I(un18_beamylt10_0));
    InMux I__2275 (
            .O(N__14219),
            .I(N__14216));
    LocalMux I__2274 (
            .O(N__14216),
            .I(if_generate_plus_mult1_un82_sum_axbxc5_0_x1));
    InMux I__2273 (
            .O(N__14213),
            .I(N__14210));
    LocalMux I__2272 (
            .O(N__14210),
            .I(if_generate_plus_mult1_un82_sum_axbxc5_0_x0));
    InMux I__2271 (
            .O(N__14207),
            .I(N__14204));
    LocalMux I__2270 (
            .O(N__14204),
            .I(N__14199));
    InMux I__2269 (
            .O(N__14203),
            .I(N__14196));
    InMux I__2268 (
            .O(N__14202),
            .I(N__14193));
    Odrv4 I__2267 (
            .O(N__14199),
            .I(un1_beamy_4));
    LocalMux I__2266 (
            .O(N__14196),
            .I(un1_beamy_4));
    LocalMux I__2265 (
            .O(N__14193),
            .I(un1_beamy_4));
    InMux I__2264 (
            .O(N__14186),
            .I(N__14181));
    InMux I__2263 (
            .O(N__14185),
            .I(N__14176));
    InMux I__2262 (
            .O(N__14184),
            .I(N__14176));
    LocalMux I__2261 (
            .O(N__14181),
            .I(N__14171));
    LocalMux I__2260 (
            .O(N__14176),
            .I(N__14171));
    Span4Mux_h I__2259 (
            .O(N__14171),
            .I(N__14168));
    Odrv4 I__2258 (
            .O(N__14168),
            .I(row_1_if_generate_plus_mult1_un68_sum_i_5));
    CascadeMux I__2257 (
            .O(N__14165),
            .I(N__14162));
    InMux I__2256 (
            .O(N__14162),
            .I(N__14159));
    LocalMux I__2255 (
            .O(N__14159),
            .I(un113_pixel_4_0_15__un4_rowZ0Z_5));
    InMux I__2254 (
            .O(N__14156),
            .I(N__14153));
    LocalMux I__2253 (
            .O(N__14153),
            .I(un113_pixel_4_0_15__un5_beamx_2Z0Z_0));
    CascadeMux I__2252 (
            .O(N__14150),
            .I(un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_));
    InMux I__2251 (
            .O(N__14147),
            .I(N__14139));
    InMux I__2250 (
            .O(N__14146),
            .I(N__14139));
    InMux I__2249 (
            .O(N__14145),
            .I(N__14136));
    InMux I__2248 (
            .O(N__14144),
            .I(N__14133));
    LocalMux I__2247 (
            .O(N__14139),
            .I(N__14126));
    LocalMux I__2246 (
            .O(N__14136),
            .I(N__14126));
    LocalMux I__2245 (
            .O(N__14133),
            .I(N__14126));
    Span4Mux_v I__2244 (
            .O(N__14126),
            .I(N__14122));
    InMux I__2243 (
            .O(N__14125),
            .I(N__14119));
    Span4Mux_h I__2242 (
            .O(N__14122),
            .I(N__14116));
    LocalMux I__2241 (
            .O(N__14119),
            .I(un5_beamx_0));
    Odrv4 I__2240 (
            .O(N__14116),
            .I(un5_beamx_0));
    CascadeMux I__2239 (
            .O(N__14111),
            .I(un5_beamx_0_cascade_));
    CascadeMux I__2238 (
            .O(N__14108),
            .I(un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_));
    InMux I__2237 (
            .O(N__14105),
            .I(N__14102));
    LocalMux I__2236 (
            .O(N__14102),
            .I(un13_beamylt6_0));
    CascadeMux I__2235 (
            .O(N__14099),
            .I(un13_beamylt6_0_cascade_));
    CascadeMux I__2234 (
            .O(N__14096),
            .I(N__14093));
    InMux I__2233 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__2232 (
            .O(N__14090),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2));
    InMux I__2231 (
            .O(N__14087),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__2230 (
            .O(N__14084),
            .I(N__14081));
    LocalMux I__2229 (
            .O(N__14081),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__2228 (
            .O(N__14078),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__2227 (
            .O(N__14075),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__2226 (
            .O(N__14072),
            .I(N__14067));
    InMux I__2225 (
            .O(N__14071),
            .I(N__14062));
    InMux I__2224 (
            .O(N__14070),
            .I(N__14062));
    LocalMux I__2223 (
            .O(N__14067),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63));
    LocalMux I__2222 (
            .O(N__14062),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63));
    InMux I__2221 (
            .O(N__14057),
            .I(N__14051));
    InMux I__2220 (
            .O(N__14056),
            .I(N__14051));
    LocalMux I__2219 (
            .O(N__14051),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__2218 (
            .O(N__14048),
            .I(N__14045));
    InMux I__2217 (
            .O(N__14045),
            .I(N__14042));
    LocalMux I__2216 (
            .O(N__14042),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__2215 (
            .O(N__14039),
            .I(N__14029));
    InMux I__2214 (
            .O(N__14038),
            .I(N__14025));
    InMux I__2213 (
            .O(N__14037),
            .I(N__14022));
    CascadeMux I__2212 (
            .O(N__14036),
            .I(N__14017));
    InMux I__2211 (
            .O(N__14035),
            .I(N__14012));
    InMux I__2210 (
            .O(N__14034),
            .I(N__14012));
    InMux I__2209 (
            .O(N__14033),
            .I(N__14009));
    InMux I__2208 (
            .O(N__14032),
            .I(N__14004));
    InMux I__2207 (
            .O(N__14029),
            .I(N__14004));
    CascadeMux I__2206 (
            .O(N__14028),
            .I(N__13998));
    LocalMux I__2205 (
            .O(N__14025),
            .I(N__13993));
    LocalMux I__2204 (
            .O(N__14022),
            .I(N__13990));
    InMux I__2203 (
            .O(N__14021),
            .I(N__13983));
    InMux I__2202 (
            .O(N__14020),
            .I(N__13983));
    InMux I__2201 (
            .O(N__14017),
            .I(N__13983));
    LocalMux I__2200 (
            .O(N__14012),
            .I(N__13976));
    LocalMux I__2199 (
            .O(N__14009),
            .I(N__13976));
    LocalMux I__2198 (
            .O(N__14004),
            .I(N__13976));
    InMux I__2197 (
            .O(N__14003),
            .I(N__13971));
    InMux I__2196 (
            .O(N__14002),
            .I(N__13971));
    InMux I__2195 (
            .O(N__14001),
            .I(N__13966));
    InMux I__2194 (
            .O(N__13998),
            .I(N__13966));
    CascadeMux I__2193 (
            .O(N__13997),
            .I(N__13962));
    InMux I__2192 (
            .O(N__13996),
            .I(N__13959));
    Span4Mux_h I__2191 (
            .O(N__13993),
            .I(N__13952));
    Span4Mux_v I__2190 (
            .O(N__13990),
            .I(N__13952));
    LocalMux I__2189 (
            .O(N__13983),
            .I(N__13952));
    Span12Mux_s11_h I__2188 (
            .O(N__13976),
            .I(N__13947));
    LocalMux I__2187 (
            .O(N__13971),
            .I(N__13947));
    LocalMux I__2186 (
            .O(N__13966),
            .I(N__13944));
    InMux I__2185 (
            .O(N__13965),
            .I(N__13939));
    InMux I__2184 (
            .O(N__13962),
            .I(N__13939));
    LocalMux I__2183 (
            .O(N__13959),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2182 (
            .O(N__13952),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum));
    Odrv12 I__2181 (
            .O(N__13947),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2180 (
            .O(N__13944),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum));
    LocalMux I__2179 (
            .O(N__13939),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum));
    CascadeMux I__2178 (
            .O(N__13928),
            .I(N__13925));
    InMux I__2177 (
            .O(N__13925),
            .I(N__13918));
    InMux I__2176 (
            .O(N__13924),
            .I(N__13915));
    InMux I__2175 (
            .O(N__13923),
            .I(N__13912));
    InMux I__2174 (
            .O(N__13922),
            .I(N__13907));
    InMux I__2173 (
            .O(N__13921),
            .I(N__13907));
    LocalMux I__2172 (
            .O(N__13918),
            .I(counterZ0Z_9));
    LocalMux I__2171 (
            .O(N__13915),
            .I(counterZ0Z_9));
    LocalMux I__2170 (
            .O(N__13912),
            .I(counterZ0Z_9));
    LocalMux I__2169 (
            .O(N__13907),
            .I(counterZ0Z_9));
    InMux I__2168 (
            .O(N__13898),
            .I(N__13892));
    InMux I__2167 (
            .O(N__13897),
            .I(N__13889));
    InMux I__2166 (
            .O(N__13896),
            .I(N__13884));
    InMux I__2165 (
            .O(N__13895),
            .I(N__13884));
    LocalMux I__2164 (
            .O(N__13892),
            .I(counterZ0Z_7));
    LocalMux I__2163 (
            .O(N__13889),
            .I(counterZ0Z_7));
    LocalMux I__2162 (
            .O(N__13884),
            .I(counterZ0Z_7));
    CascadeMux I__2161 (
            .O(N__13877),
            .I(un1_counter_1lto9_2_cascade_));
    InMux I__2160 (
            .O(N__13874),
            .I(N__13871));
    LocalMux I__2159 (
            .O(N__13871),
            .I(un10_slaveselectlt4));
    InMux I__2158 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__2157 (
            .O(N__13865),
            .I(N__13856));
    InMux I__2156 (
            .O(N__13864),
            .I(N__13852));
    InMux I__2155 (
            .O(N__13863),
            .I(N__13849));
    InMux I__2154 (
            .O(N__13862),
            .I(N__13846));
    InMux I__2153 (
            .O(N__13861),
            .I(N__13843));
    InMux I__2152 (
            .O(N__13860),
            .I(N__13840));
    InMux I__2151 (
            .O(N__13859),
            .I(N__13837));
    Span4Mux_s3_h I__2150 (
            .O(N__13856),
            .I(N__13834));
    InMux I__2149 (
            .O(N__13855),
            .I(N__13831));
    LocalMux I__2148 (
            .O(N__13852),
            .I(N__13826));
    LocalMux I__2147 (
            .O(N__13849),
            .I(N__13826));
    LocalMux I__2146 (
            .O(N__13846),
            .I(counterZ0Z_4));
    LocalMux I__2145 (
            .O(N__13843),
            .I(counterZ0Z_4));
    LocalMux I__2144 (
            .O(N__13840),
            .I(counterZ0Z_4));
    LocalMux I__2143 (
            .O(N__13837),
            .I(counterZ0Z_4));
    Odrv4 I__2142 (
            .O(N__13834),
            .I(counterZ0Z_4));
    LocalMux I__2141 (
            .O(N__13831),
            .I(counterZ0Z_4));
    Odrv12 I__2140 (
            .O(N__13826),
            .I(counterZ0Z_4));
    InMux I__2139 (
            .O(N__13811),
            .I(N__13807));
    InMux I__2138 (
            .O(N__13810),
            .I(N__13804));
    LocalMux I__2137 (
            .O(N__13807),
            .I(un1_counter_1lt9));
    LocalMux I__2136 (
            .O(N__13804),
            .I(un1_counter_1lt9));
    InMux I__2135 (
            .O(N__13799),
            .I(N__13796));
    LocalMux I__2134 (
            .O(N__13796),
            .I(N__13790));
    InMux I__2133 (
            .O(N__13795),
            .I(N__13787));
    InMux I__2132 (
            .O(N__13794),
            .I(N__13784));
    InMux I__2131 (
            .O(N__13793),
            .I(N__13781));
    Odrv4 I__2130 (
            .O(N__13790),
            .I(counterZ0Z_6));
    LocalMux I__2129 (
            .O(N__13787),
            .I(counterZ0Z_6));
    LocalMux I__2128 (
            .O(N__13784),
            .I(counterZ0Z_6));
    LocalMux I__2127 (
            .O(N__13781),
            .I(counterZ0Z_6));
    InMux I__2126 (
            .O(N__13772),
            .I(N__13768));
    InMux I__2125 (
            .O(N__13771),
            .I(N__13760));
    LocalMux I__2124 (
            .O(N__13768),
            .I(N__13757));
    InMux I__2123 (
            .O(N__13767),
            .I(N__13754));
    InMux I__2122 (
            .O(N__13766),
            .I(N__13751));
    InMux I__2121 (
            .O(N__13765),
            .I(N__13748));
    InMux I__2120 (
            .O(N__13764),
            .I(N__13745));
    InMux I__2119 (
            .O(N__13763),
            .I(N__13742));
    LocalMux I__2118 (
            .O(N__13760),
            .I(N__13739));
    Odrv4 I__2117 (
            .O(N__13757),
            .I(counterZ0Z_5));
    LocalMux I__2116 (
            .O(N__13754),
            .I(counterZ0Z_5));
    LocalMux I__2115 (
            .O(N__13751),
            .I(counterZ0Z_5));
    LocalMux I__2114 (
            .O(N__13748),
            .I(counterZ0Z_5));
    LocalMux I__2113 (
            .O(N__13745),
            .I(counterZ0Z_5));
    LocalMux I__2112 (
            .O(N__13742),
            .I(counterZ0Z_5));
    Odrv4 I__2111 (
            .O(N__13739),
            .I(counterZ0Z_5));
    InMux I__2110 (
            .O(N__13724),
            .I(N__13721));
    LocalMux I__2109 (
            .O(N__13721),
            .I(N__13714));
    InMux I__2108 (
            .O(N__13720),
            .I(N__13711));
    InMux I__2107 (
            .O(N__13719),
            .I(N__13708));
    InMux I__2106 (
            .O(N__13718),
            .I(N__13703));
    InMux I__2105 (
            .O(N__13717),
            .I(N__13703));
    Odrv4 I__2104 (
            .O(N__13714),
            .I(counterZ0Z_8));
    LocalMux I__2103 (
            .O(N__13711),
            .I(counterZ0Z_8));
    LocalMux I__2102 (
            .O(N__13708),
            .I(counterZ0Z_8));
    LocalMux I__2101 (
            .O(N__13703),
            .I(counterZ0Z_8));
    InMux I__2100 (
            .O(N__13694),
            .I(N__13691));
    LocalMux I__2099 (
            .O(N__13691),
            .I(N__13688));
    Odrv4 I__2098 (
            .O(N__13688),
            .I(slaveselect_1lto9_4));
    InMux I__2097 (
            .O(N__13685),
            .I(N__13682));
    LocalMux I__2096 (
            .O(N__13682),
            .I(slaveselect_1lto9_3));
    IoInMux I__2095 (
            .O(N__13679),
            .I(N__13675));
    IoInMux I__2094 (
            .O(N__13678),
            .I(N__13672));
    LocalMux I__2093 (
            .O(N__13675),
            .I(N__13667));
    LocalMux I__2092 (
            .O(N__13672),
            .I(N__13667));
    IoSpan4Mux I__2091 (
            .O(N__13667),
            .I(N__13664));
    Span4Mux_s3_h I__2090 (
            .O(N__13664),
            .I(N__13661));
    Odrv4 I__2089 (
            .O(N__13661),
            .I(SCLK1_0_i));
    CascadeMux I__2088 (
            .O(N__13658),
            .I(N__13655));
    InMux I__2087 (
            .O(N__13655),
            .I(N__13652));
    LocalMux I__2086 (
            .O(N__13652),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1));
    InMux I__2085 (
            .O(N__13649),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__2084 (
            .O(N__13646),
            .I(un1_sclk17_0_0_cascade_));
    InMux I__2083 (
            .O(N__13643),
            .I(N__13639));
    InMux I__2082 (
            .O(N__13642),
            .I(N__13636));
    LocalMux I__2081 (
            .O(N__13639),
            .I(N__13633));
    LocalMux I__2080 (
            .O(N__13636),
            .I(un39_0_3));
    Odrv12 I__2079 (
            .O(N__13633),
            .I(un39_0_3));
    CascadeMux I__2078 (
            .O(N__13628),
            .I(un39_0_3_cascade_));
    InMux I__2077 (
            .O(N__13625),
            .I(N__13622));
    LocalMux I__2076 (
            .O(N__13622),
            .I(N__13619));
    Odrv4 I__2075 (
            .O(N__13619),
            .I(un5_slaveselect_1));
    CascadeMux I__2074 (
            .O(N__13616),
            .I(un5_slaveselect_1_cascade_));
    InMux I__2073 (
            .O(N__13613),
            .I(N__13608));
    InMux I__2072 (
            .O(N__13612),
            .I(N__13603));
    InMux I__2071 (
            .O(N__13611),
            .I(N__13603));
    LocalMux I__2070 (
            .O(N__13608),
            .I(ScreenBuffer_1_122_1));
    LocalMux I__2069 (
            .O(N__13603),
            .I(ScreenBuffer_1_122_1));
    InMux I__2068 (
            .O(N__13598),
            .I(N__13591));
    InMux I__2067 (
            .O(N__13597),
            .I(N__13588));
    InMux I__2066 (
            .O(N__13596),
            .I(N__13581));
    InMux I__2065 (
            .O(N__13595),
            .I(N__13581));
    InMux I__2064 (
            .O(N__13594),
            .I(N__13581));
    LocalMux I__2063 (
            .O(N__13591),
            .I(N__13578));
    LocalMux I__2062 (
            .O(N__13588),
            .I(un39_0_6));
    LocalMux I__2061 (
            .O(N__13581),
            .I(un39_0_6));
    Odrv4 I__2060 (
            .O(N__13578),
            .I(un39_0_6));
    InMux I__2059 (
            .O(N__13571),
            .I(N__13568));
    LocalMux I__2058 (
            .O(N__13568),
            .I(ScreenBuffer_1_2_1_sqmuxa));
    CascadeMux I__2057 (
            .O(N__13565),
            .I(ScreenBuffer_1_2_1_sqmuxa_cascade_));
    InMux I__2056 (
            .O(N__13562),
            .I(N__13558));
    InMux I__2055 (
            .O(N__13561),
            .I(N__13550));
    LocalMux I__2054 (
            .O(N__13558),
            .I(N__13547));
    InMux I__2053 (
            .O(N__13557),
            .I(N__13540));
    InMux I__2052 (
            .O(N__13556),
            .I(N__13540));
    InMux I__2051 (
            .O(N__13555),
            .I(N__13540));
    InMux I__2050 (
            .O(N__13554),
            .I(N__13537));
    InMux I__2049 (
            .O(N__13553),
            .I(N__13534));
    LocalMux I__2048 (
            .O(N__13550),
            .I(N__13527));
    Span4Mux_h I__2047 (
            .O(N__13547),
            .I(N__13527));
    LocalMux I__2046 (
            .O(N__13540),
            .I(N__13527));
    LocalMux I__2045 (
            .O(N__13537),
            .I(un10_slaveselect));
    LocalMux I__2044 (
            .O(N__13534),
            .I(un10_slaveselect));
    Odrv4 I__2043 (
            .O(N__13527),
            .I(un10_slaveselect));
    CascadeMux I__2042 (
            .O(N__13520),
            .I(slaveselect_RNILOQC2Z0Z_0_cascade_));
    InMux I__2041 (
            .O(N__13517),
            .I(N__13513));
    InMux I__2040 (
            .O(N__13516),
            .I(N__13510));
    LocalMux I__2039 (
            .O(N__13513),
            .I(N__13507));
    LocalMux I__2038 (
            .O(N__13510),
            .I(N__13503));
    Span4Mux_h I__2037 (
            .O(N__13507),
            .I(N__13500));
    InMux I__2036 (
            .O(N__13506),
            .I(N__13497));
    Odrv4 I__2035 (
            .O(N__13503),
            .I(Z_decfrac4_2));
    Odrv4 I__2034 (
            .O(N__13500),
            .I(Z_decfrac4_2));
    LocalMux I__2033 (
            .O(N__13497),
            .I(Z_decfrac4_2));
    CascadeMux I__2032 (
            .O(N__13490),
            .I(ScreenBuffer_1_122_1_cascade_));
    InMux I__2031 (
            .O(N__13487),
            .I(N__13481));
    InMux I__2030 (
            .O(N__13486),
            .I(N__13481));
    LocalMux I__2029 (
            .O(N__13481),
            .I(ScreenBuffer_1_3_1_sqmuxa));
    InMux I__2028 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__2027 (
            .O(N__13475),
            .I(N__13472));
    Odrv4 I__2026 (
            .O(N__13472),
            .I(ScreenBuffer_1_0_1_sqmuxa));
    InMux I__2025 (
            .O(N__13469),
            .I(N__13462));
    InMux I__2024 (
            .O(N__13468),
            .I(N__13462));
    InMux I__2023 (
            .O(N__13467),
            .I(N__13459));
    LocalMux I__2022 (
            .O(N__13462),
            .I(N__13456));
    LocalMux I__2021 (
            .O(N__13459),
            .I(Z_decfrac4));
    Odrv4 I__2020 (
            .O(N__13456),
            .I(Z_decfrac4));
    InMux I__2019 (
            .O(N__13451),
            .I(N__13448));
    LocalMux I__2018 (
            .O(N__13448),
            .I(N__13445));
    Odrv4 I__2017 (
            .O(N__13445),
            .I(voltage_2_9_iv_0_0));
    CascadeMux I__2016 (
            .O(N__13442),
            .I(un1_voltage_2_1_axb_0_cascade_));
    InMux I__2015 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__2014 (
            .O(N__13436),
            .I(voltage_2_9_iv_0_2));
    InMux I__2013 (
            .O(N__13433),
            .I(N__13430));
    LocalMux I__2012 (
            .O(N__13430),
            .I(N__13427));
    Span4Mux_h I__2011 (
            .O(N__13427),
            .I(N__13424));
    Odrv4 I__2010 (
            .O(N__13424),
            .I(voltage_2_RNO_0Z0Z_2));
    InMux I__2009 (
            .O(N__13421),
            .I(N__13418));
    LocalMux I__2008 (
            .O(N__13418),
            .I(N__13415));
    Span4Mux_v I__2007 (
            .O(N__13415),
            .I(N__13409));
    InMux I__2006 (
            .O(N__13414),
            .I(N__13402));
    InMux I__2005 (
            .O(N__13413),
            .I(N__13402));
    InMux I__2004 (
            .O(N__13412),
            .I(N__13402));
    Odrv4 I__2003 (
            .O(N__13409),
            .I(un1_voltage_012_3_0));
    LocalMux I__2002 (
            .O(N__13402),
            .I(un1_voltage_012_3_0));
    InMux I__2001 (
            .O(N__13397),
            .I(N__13394));
    LocalMux I__2000 (
            .O(N__13394),
            .I(N__13391));
    Odrv4 I__1999 (
            .O(N__13391),
            .I(voltage_2_9_iv_0_1));
    InMux I__1998 (
            .O(N__13388),
            .I(N__13385));
    LocalMux I__1997 (
            .O(N__13385),
            .I(N__13382));
    Span4Mux_h I__1996 (
            .O(N__13382),
            .I(N__13379));
    Odrv4 I__1995 (
            .O(N__13379),
            .I(voltage_2_RNO_0Z0Z_1));
    InMux I__1994 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__1993 (
            .O(N__13373),
            .I(un42_cry_1_c_RNOZ0));
    InMux I__1992 (
            .O(N__13370),
            .I(N__13367));
    LocalMux I__1991 (
            .O(N__13367),
            .I(N__13364));
    Span4Mux_h I__1990 (
            .O(N__13364),
            .I(N__13361));
    Odrv4 I__1989 (
            .O(N__13361),
            .I(counter_RNIGLLH1Z0Z_0));
    InMux I__1988 (
            .O(N__13358),
            .I(N__13355));
    LocalMux I__1987 (
            .O(N__13355),
            .I(voltage_011_0));
    InMux I__1986 (
            .O(N__13352),
            .I(un42_cry_3));
    CascadeMux I__1985 (
            .O(N__13349),
            .I(N__13344));
    CascadeMux I__1984 (
            .O(N__13348),
            .I(N__13340));
    CascadeMux I__1983 (
            .O(N__13347),
            .I(N__13337));
    InMux I__1982 (
            .O(N__13344),
            .I(N__13331));
    InMux I__1981 (
            .O(N__13343),
            .I(N__13331));
    InMux I__1980 (
            .O(N__13340),
            .I(N__13326));
    InMux I__1979 (
            .O(N__13337),
            .I(N__13326));
    InMux I__1978 (
            .O(N__13336),
            .I(N__13323));
    LocalMux I__1977 (
            .O(N__13331),
            .I(N__13320));
    LocalMux I__1976 (
            .O(N__13326),
            .I(N__13317));
    LocalMux I__1975 (
            .O(N__13323),
            .I(voltage_011));
    Odrv12 I__1974 (
            .O(N__13320),
            .I(voltage_011));
    Odrv4 I__1973 (
            .O(N__13317),
            .I(voltage_011));
    InMux I__1972 (
            .O(N__13310),
            .I(N__13302));
    InMux I__1971 (
            .O(N__13309),
            .I(N__13297));
    InMux I__1970 (
            .O(N__13308),
            .I(N__13297));
    InMux I__1969 (
            .O(N__13307),
            .I(N__13294));
    InMux I__1968 (
            .O(N__13306),
            .I(N__13289));
    InMux I__1967 (
            .O(N__13305),
            .I(N__13289));
    LocalMux I__1966 (
            .O(N__13302),
            .I(N__13286));
    LocalMux I__1965 (
            .O(N__13297),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3));
    LocalMux I__1964 (
            .O(N__13294),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3));
    LocalMux I__1963 (
            .O(N__13289),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3));
    Odrv4 I__1962 (
            .O(N__13286),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3));
    CascadeMux I__1961 (
            .O(N__13277),
            .I(N__13273));
    InMux I__1960 (
            .O(N__13276),
            .I(N__13259));
    InMux I__1959 (
            .O(N__13273),
            .I(N__13256));
    InMux I__1958 (
            .O(N__13272),
            .I(N__13251));
    InMux I__1957 (
            .O(N__13271),
            .I(N__13251));
    InMux I__1956 (
            .O(N__13270),
            .I(N__13248));
    InMux I__1955 (
            .O(N__13269),
            .I(N__13239));
    InMux I__1954 (
            .O(N__13268),
            .I(N__13239));
    InMux I__1953 (
            .O(N__13267),
            .I(N__13239));
    InMux I__1952 (
            .O(N__13266),
            .I(N__13239));
    InMux I__1951 (
            .O(N__13265),
            .I(N__13232));
    InMux I__1950 (
            .O(N__13264),
            .I(N__13232));
    InMux I__1949 (
            .O(N__13263),
            .I(N__13232));
    InMux I__1948 (
            .O(N__13262),
            .I(N__13226));
    LocalMux I__1947 (
            .O(N__13259),
            .I(N__13223));
    LocalMux I__1946 (
            .O(N__13256),
            .I(N__13212));
    LocalMux I__1945 (
            .O(N__13251),
            .I(N__13212));
    LocalMux I__1944 (
            .O(N__13248),
            .I(N__13212));
    LocalMux I__1943 (
            .O(N__13239),
            .I(N__13212));
    LocalMux I__1942 (
            .O(N__13232),
            .I(N__13212));
    InMux I__1941 (
            .O(N__13231),
            .I(N__13208));
    InMux I__1940 (
            .O(N__13230),
            .I(N__13203));
    InMux I__1939 (
            .O(N__13229),
            .I(N__13203));
    LocalMux I__1938 (
            .O(N__13226),
            .I(N__13196));
    Span4Mux_s3_v I__1937 (
            .O(N__13223),
            .I(N__13196));
    Span4Mux_v I__1936 (
            .O(N__13212),
            .I(N__13196));
    InMux I__1935 (
            .O(N__13211),
            .I(N__13193));
    LocalMux I__1934 (
            .O(N__13208),
            .I(N__13190));
    LocalMux I__1933 (
            .O(N__13203),
            .I(N__13187));
    Span4Mux_h I__1932 (
            .O(N__13196),
            .I(N__13182));
    LocalMux I__1931 (
            .O(N__13193),
            .I(N__13182));
    Odrv12 I__1930 (
            .O(N__13190),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1929 (
            .O(N__13187),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1928 (
            .O(N__13182),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum));
    InMux I__1927 (
            .O(N__13175),
            .I(N__13171));
    InMux I__1926 (
            .O(N__13174),
            .I(N__13168));
    LocalMux I__1925 (
            .O(N__13171),
            .I(beamY_RNIV42D31Z0Z_6));
    LocalMux I__1924 (
            .O(N__13168),
            .I(beamY_RNIV42D31Z0Z_6));
    CascadeMux I__1923 (
            .O(N__13163),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_));
    InMux I__1922 (
            .O(N__13160),
            .I(N__13153));
    InMux I__1921 (
            .O(N__13159),
            .I(N__13150));
    InMux I__1920 (
            .O(N__13158),
            .I(N__13147));
    InMux I__1919 (
            .O(N__13157),
            .I(N__13142));
    InMux I__1918 (
            .O(N__13156),
            .I(N__13142));
    LocalMux I__1917 (
            .O(N__13153),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__1916 (
            .O(N__13150),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__1915 (
            .O(N__13147),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__1914 (
            .O(N__13142),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    InMux I__1913 (
            .O(N__13133),
            .I(N__13130));
    LocalMux I__1912 (
            .O(N__13130),
            .I(un113_pixel_3_0_11__g0_0_x2_0Z0Z_0));
    CEMux I__1911 (
            .O(N__13127),
            .I(N__13124));
    LocalMux I__1910 (
            .O(N__13124),
            .I(N__13121));
    Odrv4 I__1909 (
            .O(N__13121),
            .I(un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0));
    InMux I__1908 (
            .O(N__13118),
            .I(N__13114));
    InMux I__1907 (
            .O(N__13117),
            .I(N__13111));
    LocalMux I__1906 (
            .O(N__13114),
            .I(N__13108));
    LocalMux I__1905 (
            .O(N__13111),
            .I(N__13103));
    Span4Mux_h I__1904 (
            .O(N__13108),
            .I(N__13103));
    Odrv4 I__1903 (
            .O(N__13103),
            .I(N_1520));
    CascadeMux I__1902 (
            .O(N__13100),
            .I(N__13097));
    InMux I__1901 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__1900 (
            .O(N__13094),
            .I(N__13091));
    Span4Mux_s2_h I__1899 (
            .O(N__13091),
            .I(N__13088));
    Span4Mux_v I__1898 (
            .O(N__13088),
            .I(N__13085));
    Odrv4 I__1897 (
            .O(N__13085),
            .I(un1_voltage_2_1_cry_0_c_RNOZ0));
    InMux I__1896 (
            .O(N__13082),
            .I(N__13079));
    LocalMux I__1895 (
            .O(N__13079),
            .I(N__13076));
    Odrv4 I__1894 (
            .O(N__13076),
            .I(if_generate_plus_mult1_un75_sum_c5_x0));
    CascadeMux I__1893 (
            .O(N__13073),
            .I(if_generate_plus_mult1_un75_sum_c5_x1_cascade_));
    InMux I__1892 (
            .O(N__13070),
            .I(N__13065));
    InMux I__1891 (
            .O(N__13069),
            .I(N__13060));
    InMux I__1890 (
            .O(N__13068),
            .I(N__13060));
    LocalMux I__1889 (
            .O(N__13065),
            .I(beamY_RNIPNEA3_0Z0Z_6));
    LocalMux I__1888 (
            .O(N__13060),
            .I(beamY_RNIPNEA3_0Z0Z_6));
    InMux I__1887 (
            .O(N__13055),
            .I(N__13049));
    InMux I__1886 (
            .O(N__13054),
            .I(N__13049));
    LocalMux I__1885 (
            .O(N__13049),
            .I(beamY_RNI0K169Z0Z_6));
    InMux I__1884 (
            .O(N__13046),
            .I(N__13041));
    InMux I__1883 (
            .O(N__13045),
            .I(N__13036));
    InMux I__1882 (
            .O(N__13044),
            .I(N__13036));
    LocalMux I__1881 (
            .O(N__13041),
            .I(N__13033));
    LocalMux I__1880 (
            .O(N__13036),
            .I(N__13030));
    Odrv4 I__1879 (
            .O(N__13033),
            .I(chary_if_generate_plus_mult1_un61_sum_c4));
    Odrv4 I__1878 (
            .O(N__13030),
            .I(chary_if_generate_plus_mult1_un61_sum_c4));
    InMux I__1877 (
            .O(N__13025),
            .I(N__13022));
    LocalMux I__1876 (
            .O(N__13022),
            .I(N__13019));
    Odrv4 I__1875 (
            .O(N__13019),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9));
    CascadeMux I__1874 (
            .O(N__13016),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_));
    InMux I__1873 (
            .O(N__13013),
            .I(N__13008));
    InMux I__1872 (
            .O(N__13012),
            .I(N__13005));
    InMux I__1871 (
            .O(N__13011),
            .I(N__13002));
    LocalMux I__1870 (
            .O(N__13008),
            .I(N__12998));
    LocalMux I__1869 (
            .O(N__13005),
            .I(N__12993));
    LocalMux I__1868 (
            .O(N__13002),
            .I(N__12993));
    InMux I__1867 (
            .O(N__13001),
            .I(N__12990));
    Span4Mux_h I__1866 (
            .O(N__12998),
            .I(N__12981));
    Span4Mux_v I__1865 (
            .O(N__12993),
            .I(N__12981));
    LocalMux I__1864 (
            .O(N__12990),
            .I(N__12981));
    CascadeMux I__1863 (
            .O(N__12989),
            .I(N__12974));
    InMux I__1862 (
            .O(N__12988),
            .I(N__12967));
    Span4Mux_h I__1861 (
            .O(N__12981),
            .I(N__12964));
    InMux I__1860 (
            .O(N__12980),
            .I(N__12959));
    InMux I__1859 (
            .O(N__12979),
            .I(N__12959));
    InMux I__1858 (
            .O(N__12978),
            .I(N__12954));
    InMux I__1857 (
            .O(N__12977),
            .I(N__12954));
    InMux I__1856 (
            .O(N__12974),
            .I(N__12949));
    InMux I__1855 (
            .O(N__12973),
            .I(N__12949));
    InMux I__1854 (
            .O(N__12972),
            .I(N__12942));
    InMux I__1853 (
            .O(N__12971),
            .I(N__12942));
    InMux I__1852 (
            .O(N__12970),
            .I(N__12942));
    LocalMux I__1851 (
            .O(N__12967),
            .I(beamYZ0Z_6));
    Odrv4 I__1850 (
            .O(N__12964),
            .I(beamYZ0Z_6));
    LocalMux I__1849 (
            .O(N__12959),
            .I(beamYZ0Z_6));
    LocalMux I__1848 (
            .O(N__12954),
            .I(beamYZ0Z_6));
    LocalMux I__1847 (
            .O(N__12949),
            .I(beamYZ0Z_6));
    LocalMux I__1846 (
            .O(N__12942),
            .I(beamYZ0Z_6));
    CascadeMux I__1845 (
            .O(N__12929),
            .I(N__12925));
    CascadeMux I__1844 (
            .O(N__12928),
            .I(N__12922));
    InMux I__1843 (
            .O(N__12925),
            .I(N__12918));
    InMux I__1842 (
            .O(N__12922),
            .I(N__12915));
    InMux I__1841 (
            .O(N__12921),
            .I(N__12912));
    LocalMux I__1840 (
            .O(N__12918),
            .I(N__12908));
    LocalMux I__1839 (
            .O(N__12915),
            .I(N__12903));
    LocalMux I__1838 (
            .O(N__12912),
            .I(N__12903));
    InMux I__1837 (
            .O(N__12911),
            .I(N__12900));
    Span4Mux_h I__1836 (
            .O(N__12908),
            .I(N__12891));
    Span4Mux_v I__1835 (
            .O(N__12903),
            .I(N__12891));
    LocalMux I__1834 (
            .O(N__12900),
            .I(N__12891));
    CascadeMux I__1833 (
            .O(N__12899),
            .I(N__12887));
    InMux I__1832 (
            .O(N__12898),
            .I(N__12876));
    Span4Mux_h I__1831 (
            .O(N__12891),
            .I(N__12873));
    InMux I__1830 (
            .O(N__12890),
            .I(N__12866));
    InMux I__1829 (
            .O(N__12887),
            .I(N__12866));
    InMux I__1828 (
            .O(N__12886),
            .I(N__12866));
    InMux I__1827 (
            .O(N__12885),
            .I(N__12861));
    InMux I__1826 (
            .O(N__12884),
            .I(N__12861));
    InMux I__1825 (
            .O(N__12883),
            .I(N__12856));
    InMux I__1824 (
            .O(N__12882),
            .I(N__12856));
    InMux I__1823 (
            .O(N__12881),
            .I(N__12849));
    InMux I__1822 (
            .O(N__12880),
            .I(N__12849));
    InMux I__1821 (
            .O(N__12879),
            .I(N__12849));
    LocalMux I__1820 (
            .O(N__12876),
            .I(beamYZ0Z_5));
    Odrv4 I__1819 (
            .O(N__12873),
            .I(beamYZ0Z_5));
    LocalMux I__1818 (
            .O(N__12866),
            .I(beamYZ0Z_5));
    LocalMux I__1817 (
            .O(N__12861),
            .I(beamYZ0Z_5));
    LocalMux I__1816 (
            .O(N__12856),
            .I(beamYZ0Z_5));
    LocalMux I__1815 (
            .O(N__12849),
            .I(beamYZ0Z_5));
    InMux I__1814 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__1813 (
            .O(N__12833),
            .I(chary_if_generate_plus_mult1_un75_sum_c5_N_9));
    CascadeMux I__1812 (
            .O(N__12830),
            .I(beamY_RNIPLAE31Z0Z_4_cascade_));
    InMux I__1811 (
            .O(N__12827),
            .I(N__12824));
    LocalMux I__1810 (
            .O(N__12824),
            .I(chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0));
    CascadeMux I__1809 (
            .O(N__12821),
            .I(N__12814));
    InMux I__1808 (
            .O(N__12820),
            .I(N__12806));
    InMux I__1807 (
            .O(N__12819),
            .I(N__12806));
    InMux I__1806 (
            .O(N__12818),
            .I(N__12806));
    InMux I__1805 (
            .O(N__12817),
            .I(N__12803));
    InMux I__1804 (
            .O(N__12814),
            .I(N__12798));
    InMux I__1803 (
            .O(N__12813),
            .I(N__12798));
    LocalMux I__1802 (
            .O(N__12806),
            .I(beamY_RNIV42D31_0Z0Z_6));
    LocalMux I__1801 (
            .O(N__12803),
            .I(beamY_RNIV42D31_0Z0Z_6));
    LocalMux I__1800 (
            .O(N__12798),
            .I(beamY_RNIV42D31_0Z0Z_6));
    InMux I__1799 (
            .O(N__12791),
            .I(N__12788));
    LocalMux I__1798 (
            .O(N__12788),
            .I(un113_pixel_3_0_11__N_4_i_0));
    InMux I__1797 (
            .O(N__12785),
            .I(N__12782));
    LocalMux I__1796 (
            .O(N__12782),
            .I(g1_0_0));
    CascadeMux I__1795 (
            .O(N__12779),
            .I(row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_));
    CascadeMux I__1794 (
            .O(N__12776),
            .I(N__12772));
    CascadeMux I__1793 (
            .O(N__12775),
            .I(N__12769));
    InMux I__1792 (
            .O(N__12772),
            .I(N__12765));
    InMux I__1791 (
            .O(N__12769),
            .I(N__12762));
    CascadeMux I__1790 (
            .O(N__12768),
            .I(N__12758));
    LocalMux I__1789 (
            .O(N__12765),
            .I(N__12753));
    LocalMux I__1788 (
            .O(N__12762),
            .I(N__12753));
    CascadeMux I__1787 (
            .O(N__12761),
            .I(N__12750));
    InMux I__1786 (
            .O(N__12758),
            .I(N__12746));
    Span4Mux_h I__1785 (
            .O(N__12753),
            .I(N__12742));
    InMux I__1784 (
            .O(N__12750),
            .I(N__12737));
    InMux I__1783 (
            .O(N__12749),
            .I(N__12737));
    LocalMux I__1782 (
            .O(N__12746),
            .I(N__12734));
    InMux I__1781 (
            .O(N__12745),
            .I(N__12731));
    Odrv4 I__1780 (
            .O(N__12742),
            .I(un5_visibley_c5));
    LocalMux I__1779 (
            .O(N__12737),
            .I(un5_visibley_c5));
    Odrv4 I__1778 (
            .O(N__12734),
            .I(un5_visibley_c5));
    LocalMux I__1777 (
            .O(N__12731),
            .I(un5_visibley_c5));
    CascadeMux I__1776 (
            .O(N__12722),
            .I(N__12716));
    InMux I__1775 (
            .O(N__12721),
            .I(N__12711));
    InMux I__1774 (
            .O(N__12720),
            .I(N__12711));
    InMux I__1773 (
            .O(N__12719),
            .I(N__12708));
    InMux I__1772 (
            .O(N__12716),
            .I(N__12705));
    LocalMux I__1771 (
            .O(N__12711),
            .I(N__12702));
    LocalMux I__1770 (
            .O(N__12708),
            .I(beamY_RNIJNLCZ0Z_9));
    LocalMux I__1769 (
            .O(N__12705),
            .I(beamY_RNIJNLCZ0Z_9));
    Odrv4 I__1768 (
            .O(N__12702),
            .I(beamY_RNIJNLCZ0Z_9));
    CascadeMux I__1767 (
            .O(N__12695),
            .I(beamY_RNIJNLCZ0Z_9_cascade_));
    InMux I__1766 (
            .O(N__12692),
            .I(N__12682));
    InMux I__1765 (
            .O(N__12691),
            .I(N__12682));
    InMux I__1764 (
            .O(N__12690),
            .I(N__12679));
    InMux I__1763 (
            .O(N__12689),
            .I(N__12673));
    InMux I__1762 (
            .O(N__12688),
            .I(N__12670));
    InMux I__1761 (
            .O(N__12687),
            .I(N__12665));
    LocalMux I__1760 (
            .O(N__12682),
            .I(N__12660));
    LocalMux I__1759 (
            .O(N__12679),
            .I(N__12657));
    InMux I__1758 (
            .O(N__12678),
            .I(N__12650));
    InMux I__1757 (
            .O(N__12677),
            .I(N__12650));
    InMux I__1756 (
            .O(N__12676),
            .I(N__12650));
    LocalMux I__1755 (
            .O(N__12673),
            .I(N__12645));
    LocalMux I__1754 (
            .O(N__12670),
            .I(N__12645));
    InMux I__1753 (
            .O(N__12669),
            .I(N__12640));
    InMux I__1752 (
            .O(N__12668),
            .I(N__12640));
    LocalMux I__1751 (
            .O(N__12665),
            .I(N__12637));
    CascadeMux I__1750 (
            .O(N__12664),
            .I(N__12633));
    CascadeMux I__1749 (
            .O(N__12663),
            .I(N__12628));
    Span4Mux_v I__1748 (
            .O(N__12660),
            .I(N__12618));
    Span4Mux_v I__1747 (
            .O(N__12657),
            .I(N__12618));
    LocalMux I__1746 (
            .O(N__12650),
            .I(N__12618));
    Span4Mux_s1_v I__1745 (
            .O(N__12645),
            .I(N__12615));
    LocalMux I__1744 (
            .O(N__12640),
            .I(N__12612));
    Span4Mux_h I__1743 (
            .O(N__12637),
            .I(N__12609));
    InMux I__1742 (
            .O(N__12636),
            .I(N__12606));
    InMux I__1741 (
            .O(N__12633),
            .I(N__12597));
    InMux I__1740 (
            .O(N__12632),
            .I(N__12597));
    InMux I__1739 (
            .O(N__12631),
            .I(N__12597));
    InMux I__1738 (
            .O(N__12628),
            .I(N__12597));
    InMux I__1737 (
            .O(N__12627),
            .I(N__12590));
    InMux I__1736 (
            .O(N__12626),
            .I(N__12590));
    InMux I__1735 (
            .O(N__12625),
            .I(N__12590));
    Odrv4 I__1734 (
            .O(N__12618),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1733 (
            .O(N__12615),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    Odrv12 I__1732 (
            .O(N__12612),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1731 (
            .O(N__12609),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1730 (
            .O(N__12606),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1729 (
            .O(N__12597),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1728 (
            .O(N__12590),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum));
    CascadeMux I__1727 (
            .O(N__12575),
            .I(N__12571));
    CascadeMux I__1726 (
            .O(N__12574),
            .I(N__12568));
    InMux I__1725 (
            .O(N__12571),
            .I(N__12560));
    InMux I__1724 (
            .O(N__12568),
            .I(N__12560));
    InMux I__1723 (
            .O(N__12567),
            .I(N__12560));
    LocalMux I__1722 (
            .O(N__12560),
            .I(beamY_RNIVGU01Z0Z_9));
    CascadeMux I__1721 (
            .O(N__12557),
            .I(N__12552));
    InMux I__1720 (
            .O(N__12556),
            .I(N__12549));
    InMux I__1719 (
            .O(N__12555),
            .I(N__12546));
    InMux I__1718 (
            .O(N__12552),
            .I(N__12541));
    LocalMux I__1717 (
            .O(N__12549),
            .I(N__12536));
    LocalMux I__1716 (
            .O(N__12546),
            .I(N__12536));
    InMux I__1715 (
            .O(N__12545),
            .I(N__12533));
    InMux I__1714 (
            .O(N__12544),
            .I(N__12530));
    LocalMux I__1713 (
            .O(N__12541),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum));
    Odrv12 I__1712 (
            .O(N__12536),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum));
    LocalMux I__1711 (
            .O(N__12533),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum));
    LocalMux I__1710 (
            .O(N__12530),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum));
    CascadeMux I__1709 (
            .O(N__12521),
            .I(N__12517));
    InMux I__1708 (
            .O(N__12520),
            .I(N__12514));
    InMux I__1707 (
            .O(N__12517),
            .I(N__12511));
    LocalMux I__1706 (
            .O(N__12514),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0));
    LocalMux I__1705 (
            .O(N__12511),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0));
    CascadeMux I__1704 (
            .O(N__12506),
            .I(N__12502));
    InMux I__1703 (
            .O(N__12505),
            .I(N__12496));
    InMux I__1702 (
            .O(N__12502),
            .I(N__12496));
    InMux I__1701 (
            .O(N__12501),
            .I(N__12493));
    LocalMux I__1700 (
            .O(N__12496),
            .I(N__12490));
    LocalMux I__1699 (
            .O(N__12493),
            .I(row_1_if_generate_plus_mult1_un75_sum_ac0_5));
    Odrv4 I__1698 (
            .O(N__12490),
            .I(row_1_if_generate_plus_mult1_un75_sum_ac0_5));
    CascadeMux I__1697 (
            .O(N__12485),
            .I(N__12482));
    InMux I__1696 (
            .O(N__12482),
            .I(N__12474));
    InMux I__1695 (
            .O(N__12481),
            .I(N__12464));
    InMux I__1694 (
            .O(N__12480),
            .I(N__12459));
    InMux I__1693 (
            .O(N__12479),
            .I(N__12459));
    InMux I__1692 (
            .O(N__12478),
            .I(N__12450));
    InMux I__1691 (
            .O(N__12477),
            .I(N__12447));
    LocalMux I__1690 (
            .O(N__12474),
            .I(N__12444));
    InMux I__1689 (
            .O(N__12473),
            .I(N__12439));
    InMux I__1688 (
            .O(N__12472),
            .I(N__12439));
    InMux I__1687 (
            .O(N__12471),
            .I(N__12432));
    InMux I__1686 (
            .O(N__12470),
            .I(N__12432));
    InMux I__1685 (
            .O(N__12469),
            .I(N__12432));
    InMux I__1684 (
            .O(N__12468),
            .I(N__12427));
    InMux I__1683 (
            .O(N__12467),
            .I(N__12427));
    LocalMux I__1682 (
            .O(N__12464),
            .I(N__12422));
    LocalMux I__1681 (
            .O(N__12459),
            .I(N__12422));
    CascadeMux I__1680 (
            .O(N__12458),
            .I(N__12419));
    CascadeMux I__1679 (
            .O(N__12457),
            .I(N__12416));
    CascadeMux I__1678 (
            .O(N__12456),
            .I(N__12412));
    CascadeMux I__1677 (
            .O(N__12455),
            .I(N__12409));
    InMux I__1676 (
            .O(N__12454),
            .I(N__12402));
    InMux I__1675 (
            .O(N__12453),
            .I(N__12402));
    LocalMux I__1674 (
            .O(N__12450),
            .I(N__12397));
    LocalMux I__1673 (
            .O(N__12447),
            .I(N__12397));
    Span4Mux_v I__1672 (
            .O(N__12444),
            .I(N__12394));
    LocalMux I__1671 (
            .O(N__12439),
            .I(N__12391));
    LocalMux I__1670 (
            .O(N__12432),
            .I(N__12386));
    LocalMux I__1669 (
            .O(N__12427),
            .I(N__12386));
    Span4Mux_h I__1668 (
            .O(N__12422),
            .I(N__12383));
    InMux I__1667 (
            .O(N__12419),
            .I(N__12374));
    InMux I__1666 (
            .O(N__12416),
            .I(N__12374));
    InMux I__1665 (
            .O(N__12415),
            .I(N__12374));
    InMux I__1664 (
            .O(N__12412),
            .I(N__12374));
    InMux I__1663 (
            .O(N__12409),
            .I(N__12367));
    InMux I__1662 (
            .O(N__12408),
            .I(N__12367));
    InMux I__1661 (
            .O(N__12407),
            .I(N__12367));
    LocalMux I__1660 (
            .O(N__12402),
            .I(N__12362));
    Span4Mux_h I__1659 (
            .O(N__12397),
            .I(N__12362));
    Odrv4 I__1658 (
            .O(N__12394),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1657 (
            .O(N__12391),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1656 (
            .O(N__12386),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1655 (
            .O(N__12383),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    LocalMux I__1654 (
            .O(N__12374),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    LocalMux I__1653 (
            .O(N__12367),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1652 (
            .O(N__12362),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum));
    InMux I__1651 (
            .O(N__12347),
            .I(N__12344));
    LocalMux I__1650 (
            .O(N__12344),
            .I(N__12341));
    Odrv12 I__1649 (
            .O(N__12341),
            .I(un113_pixel_4_0_15__un1_beamylto9_3));
    IoInMux I__1648 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__1647 (
            .O(N__12335),
            .I(N__12332));
    Span4Mux_s3_v I__1646 (
            .O(N__12332),
            .I(N__12329));
    Odrv4 I__1645 (
            .O(N__12329),
            .I(VSync_c));
    CascadeMux I__1644 (
            .O(N__12326),
            .I(un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_));
    InMux I__1643 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__1642 (
            .O(N__12320),
            .I(N__12317));
    Odrv12 I__1641 (
            .O(N__12317),
            .I(beamY_RNII8O41Z0Z_9));
    InMux I__1640 (
            .O(N__12314),
            .I(N__12311));
    LocalMux I__1639 (
            .O(N__12311),
            .I(un113_pixel_4_0_15__g0_i_a3_0Z0Z_4));
    InMux I__1638 (
            .O(N__12308),
            .I(N__12305));
    LocalMux I__1637 (
            .O(N__12305),
            .I(if_m1_5));
    CascadeMux I__1636 (
            .O(N__12302),
            .I(if_generate_plus_mult1_un54_sum_axbxc5_cascade_));
    InMux I__1635 (
            .O(N__12299),
            .I(N__12294));
    InMux I__1634 (
            .O(N__12298),
            .I(N__12287));
    InMux I__1633 (
            .O(N__12297),
            .I(N__12287));
    LocalMux I__1632 (
            .O(N__12294),
            .I(N__12283));
    InMux I__1631 (
            .O(N__12293),
            .I(N__12278));
    InMux I__1630 (
            .O(N__12292),
            .I(N__12278));
    LocalMux I__1629 (
            .O(N__12287),
            .I(N__12275));
    InMux I__1628 (
            .O(N__12286),
            .I(N__12272));
    Span4Mux_h I__1627 (
            .O(N__12283),
            .I(N__12269));
    LocalMux I__1626 (
            .O(N__12278),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4));
    Odrv12 I__1625 (
            .O(N__12275),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4));
    LocalMux I__1624 (
            .O(N__12272),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4));
    Odrv4 I__1623 (
            .O(N__12269),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4));
    InMux I__1622 (
            .O(N__12260),
            .I(N__12257));
    LocalMux I__1621 (
            .O(N__12257),
            .I(if_generate_plus_mult1_un75_sum_ac0_5_x1));
    CascadeMux I__1620 (
            .O(N__12254),
            .I(row_1_if_i2_mux_0_cascade_));
    InMux I__1619 (
            .O(N__12251),
            .I(N__12248));
    LocalMux I__1618 (
            .O(N__12248),
            .I(if_generate_plus_mult1_un75_sum_ac0_5_x0));
    InMux I__1617 (
            .O(N__12245),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__1616 (
            .O(N__12242),
            .I(N__12236));
    InMux I__1615 (
            .O(N__12241),
            .I(N__12236));
    LocalMux I__1614 (
            .O(N__12236),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579));
    InMux I__1613 (
            .O(N__12233),
            .I(N__12230));
    LocalMux I__1612 (
            .O(N__12230),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4));
    InMux I__1611 (
            .O(N__12227),
            .I(N__12221));
    InMux I__1610 (
            .O(N__12226),
            .I(N__12221));
    LocalMux I__1609 (
            .O(N__12221),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36));
    InMux I__1608 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__1607 (
            .O(N__12215),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0));
    CascadeMux I__1606 (
            .O(N__12212),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_));
    InMux I__1605 (
            .O(N__12209),
            .I(N__12206));
    LocalMux I__1604 (
            .O(N__12206),
            .I(chessboardpixel_un173_pixellt10));
    InMux I__1603 (
            .O(N__12203),
            .I(N__12200));
    LocalMux I__1602 (
            .O(N__12200),
            .I(chessboardpixel_un151_pixel_27));
    CascadeMux I__1601 (
            .O(N__12197),
            .I(chessboardpixel_un177_pixel_26_cascade_));
    InMux I__1600 (
            .O(N__12194),
            .I(N__12188));
    InMux I__1599 (
            .O(N__12193),
            .I(N__12188));
    LocalMux I__1598 (
            .O(N__12188),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0));
    InMux I__1597 (
            .O(N__12185),
            .I(N__12179));
    InMux I__1596 (
            .O(N__12184),
            .I(N__12179));
    LocalMux I__1595 (
            .O(N__12179),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0));
    InMux I__1594 (
            .O(N__12176),
            .I(N__12169));
    InMux I__1593 (
            .O(N__12175),
            .I(N__12162));
    InMux I__1592 (
            .O(N__12174),
            .I(N__12162));
    InMux I__1591 (
            .O(N__12173),
            .I(N__12162));
    InMux I__1590 (
            .O(N__12172),
            .I(N__12159));
    LocalMux I__1589 (
            .O(N__12169),
            .I(beamY_i_2));
    LocalMux I__1588 (
            .O(N__12162),
            .I(beamY_i_2));
    LocalMux I__1587 (
            .O(N__12159),
            .I(beamY_i_2));
    CascadeMux I__1586 (
            .O(N__12152),
            .I(N__12147));
    InMux I__1585 (
            .O(N__12151),
            .I(N__12144));
    InMux I__1584 (
            .O(N__12150),
            .I(N__12139));
    InMux I__1583 (
            .O(N__12147),
            .I(N__12139));
    LocalMux I__1582 (
            .O(N__12144),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0));
    LocalMux I__1581 (
            .O(N__12139),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0));
    CascadeMux I__1580 (
            .O(N__12134),
            .I(un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_));
    InMux I__1579 (
            .O(N__12131),
            .I(N__12128));
    LocalMux I__1578 (
            .O(N__12128),
            .I(chessboardpixel_un199_pixellt10));
    InMux I__1577 (
            .O(N__12125),
            .I(counter_cry_4));
    InMux I__1576 (
            .O(N__12122),
            .I(counter_cry_5));
    InMux I__1575 (
            .O(N__12119),
            .I(counter_cry_6));
    InMux I__1574 (
            .O(N__12116),
            .I(counter_cry_7));
    InMux I__1573 (
            .O(N__12113),
            .I(bfn_4_14_0_));
    SRMux I__1572 (
            .O(N__12110),
            .I(N__12106));
    SRMux I__1571 (
            .O(N__12109),
            .I(N__12103));
    LocalMux I__1570 (
            .O(N__12106),
            .I(N__12099));
    LocalMux I__1569 (
            .O(N__12103),
            .I(N__12096));
    SRMux I__1568 (
            .O(N__12102),
            .I(N__12093));
    Span4Mux_h I__1567 (
            .O(N__12099),
            .I(N__12090));
    Span4Mux_s3_v I__1566 (
            .O(N__12096),
            .I(N__12085));
    LocalMux I__1565 (
            .O(N__12093),
            .I(N__12085));
    Odrv4 I__1564 (
            .O(N__12090),
            .I(un1_counter_i_0));
    Odrv4 I__1563 (
            .O(N__12085),
            .I(un1_counter_i_0));
    InMux I__1562 (
            .O(N__12080),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1561 (
            .O(N__12077),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__1560 (
            .O(N__12074),
            .I(N__12068));
    InMux I__1559 (
            .O(N__12073),
            .I(N__12068));
    LocalMux I__1558 (
            .O(N__12068),
            .I(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__1557 (
            .O(N__12065),
            .I(N__12059));
    InMux I__1556 (
            .O(N__12064),
            .I(N__12059));
    LocalMux I__1555 (
            .O(N__12059),
            .I(slaveselect_RNILOQC2Z0Z_2));
    InMux I__1554 (
            .O(N__12056),
            .I(counter_cry_1));
    InMux I__1553 (
            .O(N__12053),
            .I(counter_cry_2));
    InMux I__1552 (
            .O(N__12050),
            .I(counter_cry_3));
    CascadeMux I__1551 (
            .O(N__12047),
            .I(un1_voltage_012_0_cascade_));
    InMux I__1550 (
            .O(N__12044),
            .I(N__12039));
    CascadeMux I__1549 (
            .O(N__12043),
            .I(N__12035));
    CascadeMux I__1548 (
            .O(N__12042),
            .I(N__12032));
    LocalMux I__1547 (
            .O(N__12039),
            .I(N__12028));
    InMux I__1546 (
            .O(N__12038),
            .I(N__12025));
    InMux I__1545 (
            .O(N__12035),
            .I(N__12022));
    InMux I__1544 (
            .O(N__12032),
            .I(N__12017));
    InMux I__1543 (
            .O(N__12031),
            .I(N__12017));
    Span4Mux_h I__1542 (
            .O(N__12028),
            .I(N__12014));
    LocalMux I__1541 (
            .O(N__12025),
            .I(un74_voltage_0));
    LocalMux I__1540 (
            .O(N__12022),
            .I(un74_voltage_0));
    LocalMux I__1539 (
            .O(N__12017),
            .I(un74_voltage_0));
    Odrv4 I__1538 (
            .O(N__12014),
            .I(un74_voltage_0));
    CascadeMux I__1537 (
            .O(N__12005),
            .I(N__12000));
    InMux I__1536 (
            .O(N__12004),
            .I(N__11997));
    InMux I__1535 (
            .O(N__12003),
            .I(N__11992));
    InMux I__1534 (
            .O(N__12000),
            .I(N__11992));
    LocalMux I__1533 (
            .O(N__11997),
            .I(N__11987));
    LocalMux I__1532 (
            .O(N__11992),
            .I(N__11987));
    Span4Mux_v I__1531 (
            .O(N__11987),
            .I(N__11984));
    Odrv4 I__1530 (
            .O(N__11984),
            .I(N_1153));
    CascadeMux I__1529 (
            .O(N__11981),
            .I(N__11977));
    InMux I__1528 (
            .O(N__11980),
            .I(N__11970));
    InMux I__1527 (
            .O(N__11977),
            .I(N__11970));
    InMux I__1526 (
            .O(N__11976),
            .I(N__11967));
    CascadeMux I__1525 (
            .O(N__11975),
            .I(N__11964));
    LocalMux I__1524 (
            .O(N__11970),
            .I(N__11958));
    LocalMux I__1523 (
            .O(N__11967),
            .I(N__11955));
    InMux I__1522 (
            .O(N__11964),
            .I(N__11952));
    InMux I__1521 (
            .O(N__11963),
            .I(N__11945));
    InMux I__1520 (
            .O(N__11962),
            .I(N__11945));
    InMux I__1519 (
            .O(N__11961),
            .I(N__11945));
    Odrv4 I__1518 (
            .O(N__11958),
            .I(voltage_0_1_sqmuxa_1));
    Odrv4 I__1517 (
            .O(N__11955),
            .I(voltage_0_1_sqmuxa_1));
    LocalMux I__1516 (
            .O(N__11952),
            .I(voltage_0_1_sqmuxa_1));
    LocalMux I__1515 (
            .O(N__11945),
            .I(voltage_0_1_sqmuxa_1));
    CascadeMux I__1514 (
            .O(N__11936),
            .I(N_1153_cascade_));
    InMux I__1513 (
            .O(N__11933),
            .I(N__11928));
    InMux I__1512 (
            .O(N__11932),
            .I(N__11925));
    InMux I__1511 (
            .O(N__11931),
            .I(N__11922));
    LocalMux I__1510 (
            .O(N__11928),
            .I(N__11916));
    LocalMux I__1509 (
            .O(N__11925),
            .I(N__11916));
    LocalMux I__1508 (
            .O(N__11922),
            .I(N__11909));
    InMux I__1507 (
            .O(N__11921),
            .I(N__11906));
    Span4Mux_h I__1506 (
            .O(N__11916),
            .I(N__11903));
    InMux I__1505 (
            .O(N__11915),
            .I(N__11898));
    InMux I__1504 (
            .O(N__11914),
            .I(N__11898));
    InMux I__1503 (
            .O(N__11913),
            .I(N__11893));
    InMux I__1502 (
            .O(N__11912),
            .I(N__11893));
    Odrv4 I__1501 (
            .O(N__11909),
            .I(voltage_3_1_sqmuxa));
    LocalMux I__1500 (
            .O(N__11906),
            .I(voltage_3_1_sqmuxa));
    Odrv4 I__1499 (
            .O(N__11903),
            .I(voltage_3_1_sqmuxa));
    LocalMux I__1498 (
            .O(N__11898),
            .I(voltage_3_1_sqmuxa));
    LocalMux I__1497 (
            .O(N__11893),
            .I(voltage_3_1_sqmuxa));
    InMux I__1496 (
            .O(N__11882),
            .I(N__11879));
    LocalMux I__1495 (
            .O(N__11879),
            .I(N__11876));
    Span4Mux_v I__1494 (
            .O(N__11876),
            .I(N__11873));
    Span4Mux_h I__1493 (
            .O(N__11873),
            .I(N__11870));
    Odrv4 I__1492 (
            .O(N__11870),
            .I(voltage_3_RNO_0Z0Z_1));
    CascadeMux I__1491 (
            .O(N__11867),
            .I(voltage_3_9_iv_0_1_cascade_));
    InMux I__1490 (
            .O(N__11864),
            .I(N__11853));
    InMux I__1489 (
            .O(N__11863),
            .I(N__11853));
    InMux I__1488 (
            .O(N__11862),
            .I(N__11848));
    InMux I__1487 (
            .O(N__11861),
            .I(N__11848));
    InMux I__1486 (
            .O(N__11860),
            .I(N__11841));
    InMux I__1485 (
            .O(N__11859),
            .I(N__11841));
    InMux I__1484 (
            .O(N__11858),
            .I(N__11841));
    LocalMux I__1483 (
            .O(N__11853),
            .I(N__11836));
    LocalMux I__1482 (
            .O(N__11848),
            .I(N__11833));
    LocalMux I__1481 (
            .O(N__11841),
            .I(N__11830));
    InMux I__1480 (
            .O(N__11840),
            .I(N__11825));
    InMux I__1479 (
            .O(N__11839),
            .I(N__11825));
    Span4Mux_s3_h I__1478 (
            .O(N__11836),
            .I(N__11822));
    Span4Mux_v I__1477 (
            .O(N__11833),
            .I(N__11819));
    Span4Mux_s3_h I__1476 (
            .O(N__11830),
            .I(N__11816));
    LocalMux I__1475 (
            .O(N__11825),
            .I(un1_voltage_012_0));
    Odrv4 I__1474 (
            .O(N__11822),
            .I(un1_voltage_012_0));
    Odrv4 I__1473 (
            .O(N__11819),
            .I(un1_voltage_012_0));
    Odrv4 I__1472 (
            .O(N__11816),
            .I(un1_voltage_012_0));
    InMux I__1471 (
            .O(N__11807),
            .I(N__11804));
    LocalMux I__1470 (
            .O(N__11804),
            .I(N__11801));
    Odrv4 I__1469 (
            .O(N__11801),
            .I(voltage_1_9_iv_0_1));
    CascadeMux I__1468 (
            .O(N__11798),
            .I(N__11795));
    InMux I__1467 (
            .O(N__11795),
            .I(N__11792));
    LocalMux I__1466 (
            .O(N__11792),
            .I(N__11789));
    Span4Mux_v I__1465 (
            .O(N__11789),
            .I(N__11786));
    Odrv4 I__1464 (
            .O(N__11786),
            .I(voltage_1_RNO_0Z0Z_1));
    CascadeMux I__1463 (
            .O(N__11783),
            .I(N_1504_cascade_));
    InMux I__1462 (
            .O(N__11780),
            .I(N__11777));
    LocalMux I__1461 (
            .O(N__11777),
            .I(N_1504));
    InMux I__1460 (
            .O(N__11774),
            .I(N__11766));
    InMux I__1459 (
            .O(N__11773),
            .I(N__11766));
    InMux I__1458 (
            .O(N__11772),
            .I(N__11762));
    InMux I__1457 (
            .O(N__11771),
            .I(N__11758));
    LocalMux I__1456 (
            .O(N__11766),
            .I(N__11755));
    InMux I__1455 (
            .O(N__11765),
            .I(N__11752));
    LocalMux I__1454 (
            .O(N__11762),
            .I(N__11749));
    InMux I__1453 (
            .O(N__11761),
            .I(N__11746));
    LocalMux I__1452 (
            .O(N__11758),
            .I(N__11743));
    Span4Mux_s3_h I__1451 (
            .O(N__11755),
            .I(N__11740));
    LocalMux I__1450 (
            .O(N__11752),
            .I(N__11735));
    Span4Mux_s3_h I__1449 (
            .O(N__11749),
            .I(N__11735));
    LocalMux I__1448 (
            .O(N__11746),
            .I(counter_RNI8DLH1Z0Z_0));
    Odrv4 I__1447 (
            .O(N__11743),
            .I(counter_RNI8DLH1Z0Z_0));
    Odrv4 I__1446 (
            .O(N__11740),
            .I(counter_RNI8DLH1Z0Z_0));
    Odrv4 I__1445 (
            .O(N__11735),
            .I(counter_RNI8DLH1Z0Z_0));
    InMux I__1444 (
            .O(N__11726),
            .I(N__11721));
    CascadeMux I__1443 (
            .O(N__11725),
            .I(N__11718));
    CascadeMux I__1442 (
            .O(N__11724),
            .I(N__11715));
    LocalMux I__1441 (
            .O(N__11721),
            .I(N__11711));
    InMux I__1440 (
            .O(N__11718),
            .I(N__11704));
    InMux I__1439 (
            .O(N__11715),
            .I(N__11704));
    InMux I__1438 (
            .O(N__11714),
            .I(N__11704));
    Odrv4 I__1437 (
            .O(N__11711),
            .I(N_1508));
    LocalMux I__1436 (
            .O(N__11704),
            .I(N_1508));
    InMux I__1435 (
            .O(N__11699),
            .I(N__11690));
    InMux I__1434 (
            .O(N__11698),
            .I(N__11690));
    InMux I__1433 (
            .O(N__11697),
            .I(N__11690));
    LocalMux I__1432 (
            .O(N__11690),
            .I(N__11687));
    Odrv12 I__1431 (
            .O(N__11687),
            .I(N_1159_i));
    InMux I__1430 (
            .O(N__11684),
            .I(N__11681));
    LocalMux I__1429 (
            .O(N__11681),
            .I(N__11675));
    InMux I__1428 (
            .O(N__11680),
            .I(N__11668));
    InMux I__1427 (
            .O(N__11679),
            .I(N__11668));
    InMux I__1426 (
            .O(N__11678),
            .I(N__11668));
    Span4Mux_h I__1425 (
            .O(N__11675),
            .I(N__11665));
    LocalMux I__1424 (
            .O(N__11668),
            .I(N_1154));
    Odrv4 I__1423 (
            .O(N__11665),
            .I(N_1154));
    CascadeMux I__1422 (
            .O(N__11660),
            .I(N_1159_i_cascade_));
    CascadeMux I__1421 (
            .O(N__11657),
            .I(N__11652));
    InMux I__1420 (
            .O(N__11656),
            .I(N__11649));
    InMux I__1419 (
            .O(N__11655),
            .I(N__11646));
    InMux I__1418 (
            .O(N__11652),
            .I(N__11639));
    LocalMux I__1417 (
            .O(N__11649),
            .I(N__11634));
    LocalMux I__1416 (
            .O(N__11646),
            .I(N__11634));
    InMux I__1415 (
            .O(N__11645),
            .I(N__11631));
    InMux I__1414 (
            .O(N__11644),
            .I(N__11624));
    InMux I__1413 (
            .O(N__11643),
            .I(N__11624));
    InMux I__1412 (
            .O(N__11642),
            .I(N__11624));
    LocalMux I__1411 (
            .O(N__11639),
            .I(N__11619));
    Span4Mux_h I__1410 (
            .O(N__11634),
            .I(N__11619));
    LocalMux I__1409 (
            .O(N__11631),
            .I(voltage_2_1_sqmuxa));
    LocalMux I__1408 (
            .O(N__11624),
            .I(voltage_2_1_sqmuxa));
    Odrv4 I__1407 (
            .O(N__11619),
            .I(voltage_2_1_sqmuxa));
    IoInMux I__1406 (
            .O(N__11612),
            .I(N__11609));
    LocalMux I__1405 (
            .O(N__11609),
            .I(N__11606));
    Span4Mux_s3_h I__1404 (
            .O(N__11606),
            .I(N__11603));
    Odrv4 I__1403 (
            .O(N__11603),
            .I(voltage_0_0_sqmuxa_1));
    InMux I__1402 (
            .O(N__11600),
            .I(N__11597));
    LocalMux I__1401 (
            .O(N__11597),
            .I(slaveselect_RNILOQC2Z0Z_1));
    CascadeMux I__1400 (
            .O(N__11594),
            .I(slaveselect_RNILOQC2Z0Z_1_cascade_));
    InMux I__1399 (
            .O(N__11591),
            .I(N__11588));
    LocalMux I__1398 (
            .O(N__11588),
            .I(N__11584));
    InMux I__1397 (
            .O(N__11587),
            .I(N__11581));
    Span4Mux_v I__1396 (
            .O(N__11584),
            .I(N__11578));
    LocalMux I__1395 (
            .O(N__11581),
            .I(counter_RNICHLH1Z0Z_0));
    Odrv4 I__1394 (
            .O(N__11578),
            .I(counter_RNICHLH1Z0Z_0));
    InMux I__1393 (
            .O(N__11573),
            .I(N__11570));
    LocalMux I__1392 (
            .O(N__11570),
            .I(un5_visibley_0_29));
    CascadeMux I__1391 (
            .O(N__11567),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_));
    CascadeMux I__1390 (
            .O(N__11564),
            .I(if_m1_x1_cascade_));
    InMux I__1389 (
            .O(N__11561),
            .I(N__11557));
    InMux I__1388 (
            .O(N__11560),
            .I(N__11553));
    LocalMux I__1387 (
            .O(N__11557),
            .I(N__11550));
    InMux I__1386 (
            .O(N__11556),
            .I(N__11547));
    LocalMux I__1385 (
            .O(N__11553),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    Odrv4 I__1384 (
            .O(N__11550),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    LocalMux I__1383 (
            .O(N__11547),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    InMux I__1382 (
            .O(N__11540),
            .I(N__11534));
    InMux I__1381 (
            .O(N__11539),
            .I(N__11534));
    LocalMux I__1380 (
            .O(N__11534),
            .I(N__11531));
    Span4Mux_h I__1379 (
            .O(N__11531),
            .I(N__11523));
    InMux I__1378 (
            .O(N__11530),
            .I(N__11516));
    InMux I__1377 (
            .O(N__11529),
            .I(N__11516));
    InMux I__1376 (
            .O(N__11528),
            .I(N__11516));
    InMux I__1375 (
            .O(N__11527),
            .I(N__11511));
    InMux I__1374 (
            .O(N__11526),
            .I(N__11511));
    Odrv4 I__1373 (
            .O(N__11523),
            .I(row_1_if_generate_plus_mult1_un61_sum_axb4_i));
    LocalMux I__1372 (
            .O(N__11516),
            .I(row_1_if_generate_plus_mult1_un61_sum_axb4_i));
    LocalMux I__1371 (
            .O(N__11511),
            .I(row_1_if_generate_plus_mult1_un61_sum_axb4_i));
    InMux I__1370 (
            .O(N__11504),
            .I(N__11501));
    LocalMux I__1369 (
            .O(N__11501),
            .I(if_m1_x0));
    InMux I__1368 (
            .O(N__11498),
            .I(N__11495));
    LocalMux I__1367 (
            .O(N__11495),
            .I(un113_pixel_3_0_11__g1_0));
    CascadeMux I__1366 (
            .O(N__11492),
            .I(chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_));
    IoInMux I__1365 (
            .O(N__11489),
            .I(N__11486));
    LocalMux I__1364 (
            .O(N__11486),
            .I(N__11483));
    Span4Mux_s3_h I__1363 (
            .O(N__11483),
            .I(N__11480));
    Span4Mux_v I__1362 (
            .O(N__11480),
            .I(N__11477));
    Odrv4 I__1361 (
            .O(N__11477),
            .I(GB_BUFFER_Clock12MHz_c_g_THRU_CO));
    CascadeMux I__1360 (
            .O(N__11474),
            .I(beamY_RNIQTGS2Z0Z_8_cascade_));
    CascadeMux I__1359 (
            .O(N__11471),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_));
    CascadeMux I__1358 (
            .O(N__11468),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_cascade_));
    InMux I__1357 (
            .O(N__11465),
            .I(N__11459));
    InMux I__1356 (
            .O(N__11464),
            .I(N__11459));
    LocalMux I__1355 (
            .O(N__11459),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0));
    CascadeMux I__1354 (
            .O(N__11456),
            .I(N__11451));
    InMux I__1353 (
            .O(N__11455),
            .I(N__11438));
    InMux I__1352 (
            .O(N__11454),
            .I(N__11438));
    InMux I__1351 (
            .O(N__11451),
            .I(N__11438));
    InMux I__1350 (
            .O(N__11450),
            .I(N__11438));
    InMux I__1349 (
            .O(N__11449),
            .I(N__11438));
    LocalMux I__1348 (
            .O(N__11438),
            .I(beamY_RNIQTGS2Z0Z_8));
    InMux I__1347 (
            .O(N__11435),
            .I(N__11429));
    InMux I__1346 (
            .O(N__11434),
            .I(N__11429));
    LocalMux I__1345 (
            .O(N__11429),
            .I(chary_if_generate_plus_mult1_un54_sum_c4));
    CascadeMux I__1344 (
            .O(N__11426),
            .I(beamY_RNI0K169Z0Z_6_cascade_));
    InMux I__1343 (
            .O(N__11423),
            .I(N__11420));
    LocalMux I__1342 (
            .O(N__11420),
            .I(chary_if_generate_plus_mult1_un61_sum_c4_3_1));
    CascadeMux I__1341 (
            .O(N__11417),
            .I(chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_));
    CascadeMux I__1340 (
            .O(N__11414),
            .I(N__11410));
    InMux I__1339 (
            .O(N__11413),
            .I(N__11405));
    InMux I__1338 (
            .O(N__11410),
            .I(N__11405));
    LocalMux I__1337 (
            .O(N__11405),
            .I(N__11401));
    InMux I__1336 (
            .O(N__11404),
            .I(N__11398));
    Odrv4 I__1335 (
            .O(N__11401),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0));
    LocalMux I__1334 (
            .O(N__11398),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0));
    InMux I__1333 (
            .O(N__11393),
            .I(N__11390));
    LocalMux I__1332 (
            .O(N__11390),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_2));
    CascadeMux I__1331 (
            .O(N__11387),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_));
    InMux I__1330 (
            .O(N__11384),
            .I(N__11378));
    InMux I__1329 (
            .O(N__11383),
            .I(N__11378));
    LocalMux I__1328 (
            .O(N__11378),
            .I(N__11374));
    InMux I__1327 (
            .O(N__11377),
            .I(N__11371));
    Span4Mux_h I__1326 (
            .O(N__11374),
            .I(N__11368));
    LocalMux I__1325 (
            .O(N__11371),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0));
    Odrv4 I__1324 (
            .O(N__11368),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0));
    CascadeMux I__1323 (
            .O(N__11363),
            .I(N__11360));
    InMux I__1322 (
            .O(N__11360),
            .I(N__11353));
    InMux I__1321 (
            .O(N__11359),
            .I(N__11353));
    InMux I__1320 (
            .O(N__11358),
            .I(N__11350));
    LocalMux I__1319 (
            .O(N__11353),
            .I(N__11347));
    LocalMux I__1318 (
            .O(N__11350),
            .I(N__11344));
    Span4Mux_h I__1317 (
            .O(N__11347),
            .I(N__11341));
    Odrv4 I__1316 (
            .O(N__11344),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0));
    Odrv4 I__1315 (
            .O(N__11341),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0));
    InMux I__1314 (
            .O(N__11336),
            .I(N__11331));
    InMux I__1313 (
            .O(N__11335),
            .I(N__11326));
    InMux I__1312 (
            .O(N__11334),
            .I(N__11326));
    LocalMux I__1311 (
            .O(N__11331),
            .I(N__11323));
    LocalMux I__1310 (
            .O(N__11326),
            .I(N__11320));
    Odrv12 I__1309 (
            .O(N__11323),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0));
    Odrv12 I__1308 (
            .O(N__11320),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0));
    CascadeMux I__1307 (
            .O(N__11315),
            .I(N__11312));
    InMux I__1306 (
            .O(N__11312),
            .I(N__11309));
    LocalMux I__1305 (
            .O(N__11309),
            .I(beamY_RNIFS4TZ0Z_7));
    CascadeMux I__1304 (
            .O(N__11306),
            .I(beamY_RNIFS4TZ0Z_7_cascade_));
    CascadeMux I__1303 (
            .O(N__11303),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_));
    InMux I__1302 (
            .O(N__11300),
            .I(N__11297));
    LocalMux I__1301 (
            .O(N__11297),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__1300 (
            .O(N__11294),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6));
    CascadeMux I__1299 (
            .O(N__11291),
            .I(N__11288));
    InMux I__1298 (
            .O(N__11288),
            .I(N__11285));
    LocalMux I__1297 (
            .O(N__11285),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0));
    CascadeMux I__1296 (
            .O(N__11282),
            .I(N__11279));
    InMux I__1295 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__1294 (
            .O(N__11276),
            .I(N__11273));
    Odrv4 I__1293 (
            .O(N__11273),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__1292 (
            .O(N__11270),
            .I(N__11267));
    LocalMux I__1291 (
            .O(N__11267),
            .I(N__11264));
    Span4Mux_h I__1290 (
            .O(N__11264),
            .I(N__11260));
    InMux I__1289 (
            .O(N__11263),
            .I(N__11257));
    Odrv4 I__1288 (
            .O(N__11260),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0));
    LocalMux I__1287 (
            .O(N__11257),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0));
    InMux I__1286 (
            .O(N__11252),
            .I(N__11249));
    LocalMux I__1285 (
            .O(N__11249),
            .I(N__11242));
    InMux I__1284 (
            .O(N__11248),
            .I(N__11239));
    InMux I__1283 (
            .O(N__11247),
            .I(N__11236));
    InMux I__1282 (
            .O(N__11246),
            .I(N__11231));
    InMux I__1281 (
            .O(N__11245),
            .I(N__11231));
    Odrv4 I__1280 (
            .O(N__11242),
            .I(un5_visibley_c2));
    LocalMux I__1279 (
            .O(N__11239),
            .I(un5_visibley_c2));
    LocalMux I__1278 (
            .O(N__11236),
            .I(un5_visibley_c2));
    LocalMux I__1277 (
            .O(N__11231),
            .I(un5_visibley_c2));
    CascadeMux I__1276 (
            .O(N__11222),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_));
    InMux I__1275 (
            .O(N__11219),
            .I(N__11216));
    LocalMux I__1274 (
            .O(N__11216),
            .I(beamY_RNIEDF31Z0Z_6));
    CascadeMux I__1273 (
            .O(N__11213),
            .I(chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_));
    CascadeMux I__1272 (
            .O(N__11210),
            .I(N__11207));
    InMux I__1271 (
            .O(N__11207),
            .I(N__11204));
    LocalMux I__1270 (
            .O(N__11204),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246));
    InMux I__1269 (
            .O(N__11201),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1268 (
            .O(N__11198),
            .I(N__11195));
    LocalMux I__1267 (
            .O(N__11195),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__1266 (
            .O(N__11192),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__1265 (
            .O(N__11189),
            .I(N__11184));
    InMux I__1264 (
            .O(N__11188),
            .I(N__11179));
    InMux I__1263 (
            .O(N__11187),
            .I(N__11170));
    InMux I__1262 (
            .O(N__11184),
            .I(N__11170));
    InMux I__1261 (
            .O(N__11183),
            .I(N__11170));
    InMux I__1260 (
            .O(N__11182),
            .I(N__11170));
    LocalMux I__1259 (
            .O(N__11179),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8));
    LocalMux I__1258 (
            .O(N__11170),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8));
    InMux I__1257 (
            .O(N__11165),
            .I(N__11162));
    LocalMux I__1256 (
            .O(N__11162),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__1255 (
            .O(N__11159),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__1254 (
            .O(N__11156),
            .I(N__11153));
    InMux I__1253 (
            .O(N__11153),
            .I(N__11150));
    LocalMux I__1252 (
            .O(N__11150),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79));
    InMux I__1251 (
            .O(N__11147),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    CascadeMux I__1250 (
            .O(N__11144),
            .I(N__11141));
    InMux I__1249 (
            .O(N__11141),
            .I(N__11138));
    LocalMux I__1248 (
            .O(N__11138),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0));
    InMux I__1247 (
            .O(N__11135),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1246 (
            .O(N__11132),
            .I(N__11129));
    InMux I__1245 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__1244 (
            .O(N__11126),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0));
    InMux I__1243 (
            .O(N__11123),
            .I(N__11114));
    InMux I__1242 (
            .O(N__11122),
            .I(N__11114));
    InMux I__1241 (
            .O(N__11121),
            .I(N__11111));
    InMux I__1240 (
            .O(N__11120),
            .I(N__11106));
    InMux I__1239 (
            .O(N__11119),
            .I(N__11106));
    LocalMux I__1238 (
            .O(N__11114),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0));
    LocalMux I__1237 (
            .O(N__11111),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0));
    LocalMux I__1236 (
            .O(N__11106),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0));
    InMux I__1235 (
            .O(N__11099),
            .I(N__11096));
    LocalMux I__1234 (
            .O(N__11096),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7));
    CascadeMux I__1233 (
            .O(N__11093),
            .I(N__11090));
    InMux I__1232 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__1231 (
            .O(N__11087),
            .I(N__11084));
    Odrv12 I__1230 (
            .O(N__11084),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1));
    InMux I__1229 (
            .O(N__11081),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__1228 (
            .O(N__11078),
            .I(N__11075));
    InMux I__1227 (
            .O(N__11075),
            .I(N__11072));
    LocalMux I__1226 (
            .O(N__11072),
            .I(N__11069));
    Odrv4 I__1225 (
            .O(N__11069),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2));
    InMux I__1224 (
            .O(N__11066),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__1223 (
            .O(N__11063),
            .I(N__11060));
    InMux I__1222 (
            .O(N__11060),
            .I(N__11057));
    LocalMux I__1221 (
            .O(N__11057),
            .I(N__11054));
    Odrv4 I__1220 (
            .O(N__11054),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513));
    InMux I__1219 (
            .O(N__11051),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1218 (
            .O(N__11048),
            .I(N__11045));
    LocalMux I__1217 (
            .O(N__11045),
            .I(N__11042));
    Odrv4 I__1216 (
            .O(N__11042),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__1215 (
            .O(N__11039),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1214 (
            .O(N__11036),
            .I(N__11029));
    InMux I__1213 (
            .O(N__11035),
            .I(N__11022));
    InMux I__1212 (
            .O(N__11034),
            .I(N__11022));
    InMux I__1211 (
            .O(N__11033),
            .I(N__11022));
    InMux I__1210 (
            .O(N__11032),
            .I(N__11019));
    LocalMux I__1209 (
            .O(N__11029),
            .I(N__11014));
    LocalMux I__1208 (
            .O(N__11022),
            .I(N__11014));
    LocalMux I__1207 (
            .O(N__11019),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73));
    Odrv4 I__1206 (
            .O(N__11014),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73));
    InMux I__1205 (
            .O(N__11009),
            .I(N__11006));
    LocalMux I__1204 (
            .O(N__11006),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__1203 (
            .O(N__11003),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1202 (
            .O(N__11000),
            .I(N__10997));
    LocalMux I__1201 (
            .O(N__10997),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404));
    InMux I__1200 (
            .O(N__10994),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__1199 (
            .O(N__10991),
            .I(N__10988));
    InMux I__1198 (
            .O(N__10988),
            .I(N__10985));
    LocalMux I__1197 (
            .O(N__10985),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45));
    InMux I__1196 (
            .O(N__10982),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__1195 (
            .O(N__10979),
            .I(N__10976));
    LocalMux I__1194 (
            .O(N__10976),
            .I(counter_RNI2RBA2Z0Z_3));
    InMux I__1193 (
            .O(N__10973),
            .I(un1_voltage_2_1_cry_1));
    InMux I__1192 (
            .O(N__10970),
            .I(N__10967));
    LocalMux I__1191 (
            .O(N__10967),
            .I(un1_voltage_2_1_axb_3));
    CascadeMux I__1190 (
            .O(N__10964),
            .I(N__10961));
    InMux I__1189 (
            .O(N__10961),
            .I(N__10958));
    LocalMux I__1188 (
            .O(N__10958),
            .I(N__10955));
    Odrv4 I__1187 (
            .O(N__10955),
            .I(voltage_2_9_iv_0_3));
    InMux I__1186 (
            .O(N__10952),
            .I(un1_voltage_2_1_cry_2));
    InMux I__1185 (
            .O(N__10949),
            .I(N__10941));
    InMux I__1184 (
            .O(N__10948),
            .I(N__10941));
    InMux I__1183 (
            .O(N__10947),
            .I(N__10936));
    InMux I__1182 (
            .O(N__10946),
            .I(N__10936));
    LocalMux I__1181 (
            .O(N__10941),
            .I(N__10933));
    LocalMux I__1180 (
            .O(N__10936),
            .I(N_46_1));
    Odrv4 I__1179 (
            .O(N__10933),
            .I(N_46_1));
    CascadeMux I__1178 (
            .O(N__10928),
            .I(un1_sclk17_2_1_cascade_));
    CascadeMux I__1177 (
            .O(N__10925),
            .I(un1_sclk17_1_1_cascade_));
    CascadeMux I__1176 (
            .O(N__10922),
            .I(N__10919));
    InMux I__1175 (
            .O(N__10919),
            .I(N__10916));
    LocalMux I__1174 (
            .O(N__10916),
            .I(N__10913));
    Odrv12 I__1173 (
            .O(N__10913),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__1172 (
            .O(N__10910),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__1171 (
            .O(N__10907),
            .I(N__10904));
    InMux I__1170 (
            .O(N__10904),
            .I(N__10901));
    LocalMux I__1169 (
            .O(N__10901),
            .I(counter_RNILOUG2Z0Z_3));
    InMux I__1168 (
            .O(N__10898),
            .I(un1_voltage_1_1_cry_0));
    InMux I__1167 (
            .O(N__10895),
            .I(N__10892));
    LocalMux I__1166 (
            .O(N__10892),
            .I(counter_RNIT58K2Z0Z_2));
    InMux I__1165 (
            .O(N__10889),
            .I(N__10886));
    LocalMux I__1164 (
            .O(N__10886),
            .I(N__10883));
    Odrv12 I__1163 (
            .O(N__10883),
            .I(voltage_1_RNO_0Z0Z_2));
    InMux I__1162 (
            .O(N__10880),
            .I(un1_voltage_1_1_cry_1));
    InMux I__1161 (
            .O(N__10877),
            .I(un1_voltage_1_1_cry_2));
    InMux I__1160 (
            .O(N__10874),
            .I(N__10871));
    LocalMux I__1159 (
            .O(N__10871),
            .I(voltage_1_RNO_0Z0Z_3));
    CascadeMux I__1158 (
            .O(N__10868),
            .I(un6_slaveselectlto9_1_cascade_));
    CascadeMux I__1157 (
            .O(N__10865),
            .I(un6_slaveselect_0_cascade_));
    InMux I__1156 (
            .O(N__10862),
            .I(N__10859));
    LocalMux I__1155 (
            .O(N__10859),
            .I(un3_slaveselectlt9));
    CascadeMux I__1154 (
            .O(N__10856),
            .I(N__10853));
    InMux I__1153 (
            .O(N__10853),
            .I(N__10850));
    LocalMux I__1152 (
            .O(N__10850),
            .I(N__10847));
    Odrv4 I__1151 (
            .O(N__10847),
            .I(voltage_2_RNIKG123Z0Z_1));
    InMux I__1150 (
            .O(N__10844),
            .I(un1_voltage_2_1_cry_0));
    CascadeMux I__1149 (
            .O(N__10841),
            .I(voltage_1_1_sqmuxa_cascade_));
    InMux I__1148 (
            .O(N__10838),
            .I(N__10835));
    LocalMux I__1147 (
            .O(N__10835),
            .I(voltage_1_9_iv_0_3));
    InMux I__1146 (
            .O(N__10832),
            .I(N__10829));
    LocalMux I__1145 (
            .O(N__10829),
            .I(voltage_3_RNO_0Z0Z_3));
    InMux I__1144 (
            .O(N__10826),
            .I(N__10823));
    LocalMux I__1143 (
            .O(N__10823),
            .I(voltage_3_9_iv_0_3));
    InMux I__1142 (
            .O(N__10820),
            .I(N__10817));
    LocalMux I__1141 (
            .O(N__10817),
            .I(N__10813));
    InMux I__1140 (
            .O(N__10816),
            .I(N__10810));
    Odrv4 I__1139 (
            .O(N__10813),
            .I(N_1510));
    LocalMux I__1138 (
            .O(N__10810),
            .I(N_1510));
    CascadeMux I__1137 (
            .O(N__10805),
            .I(N_1506_cascade_));
    CascadeMux I__1136 (
            .O(N__10802),
            .I(counter_RNIGLLH1Z0Z_0_cascade_));
    InMux I__1135 (
            .O(N__10799),
            .I(N__10796));
    LocalMux I__1134 (
            .O(N__10796),
            .I(N__10790));
    InMux I__1133 (
            .O(N__10795),
            .I(N__10783));
    InMux I__1132 (
            .O(N__10794),
            .I(N__10783));
    InMux I__1131 (
            .O(N__10793),
            .I(N__10783));
    Odrv4 I__1130 (
            .O(N__10790),
            .I(N_2063));
    LocalMux I__1129 (
            .O(N__10783),
            .I(N_2063));
    InMux I__1128 (
            .O(N__10778),
            .I(N__10775));
    LocalMux I__1127 (
            .O(N__10775),
            .I(N__10772));
    Odrv4 I__1126 (
            .O(N__10772),
            .I(N_1522));
    CascadeMux I__1125 (
            .O(N__10769),
            .I(N__10766));
    InMux I__1124 (
            .O(N__10766),
            .I(N__10763));
    LocalMux I__1123 (
            .O(N__10763),
            .I(N__10760));
    Odrv4 I__1122 (
            .O(N__10760),
            .I(un1_voltage_1_1_cry_0_0_c_RNOZ0));
    InMux I__1121 (
            .O(N__10757),
            .I(N__10751));
    InMux I__1120 (
            .O(N__10756),
            .I(N__10751));
    LocalMux I__1119 (
            .O(N__10751),
            .I(N_1521));
    InMux I__1118 (
            .O(N__10748),
            .I(N__10743));
    InMux I__1117 (
            .O(N__10747),
            .I(N__10738));
    InMux I__1116 (
            .O(N__10746),
            .I(N__10738));
    LocalMux I__1115 (
            .O(N__10743),
            .I(counter_RNI49LH1_0Z0Z_0));
    LocalMux I__1114 (
            .O(N__10738),
            .I(counter_RNI49LH1_0Z0Z_0));
    InMux I__1113 (
            .O(N__10733),
            .I(N__10730));
    LocalMux I__1112 (
            .O(N__10730),
            .I(voltage_1_9_iv_0_0));
    InMux I__1111 (
            .O(N__10727),
            .I(N__10721));
    InMux I__1110 (
            .O(N__10726),
            .I(N__10721));
    LocalMux I__1109 (
            .O(N__10721),
            .I(CO1_3));
    CascadeMux I__1108 (
            .O(N__10718),
            .I(voltage_2_1_sqmuxa_cascade_));
    InMux I__1107 (
            .O(N__10715),
            .I(N__10706));
    InMux I__1106 (
            .O(N__10714),
            .I(N__10706));
    InMux I__1105 (
            .O(N__10713),
            .I(N__10706));
    LocalMux I__1104 (
            .O(N__10706),
            .I(N_1155));
    CascadeMux I__1103 (
            .O(N__10703),
            .I(N__10699));
    CascadeMux I__1102 (
            .O(N__10702),
            .I(N__10696));
    InMux I__1101 (
            .O(N__10699),
            .I(N__10689));
    InMux I__1100 (
            .O(N__10696),
            .I(N__10689));
    CascadeMux I__1099 (
            .O(N__10695),
            .I(N__10686));
    CascadeMux I__1098 (
            .O(N__10694),
            .I(N__10680));
    LocalMux I__1097 (
            .O(N__10689),
            .I(N__10677));
    InMux I__1096 (
            .O(N__10686),
            .I(N__10674));
    InMux I__1095 (
            .O(N__10685),
            .I(N__10671));
    InMux I__1094 (
            .O(N__10684),
            .I(N__10666));
    InMux I__1093 (
            .O(N__10683),
            .I(N__10666));
    InMux I__1092 (
            .O(N__10680),
            .I(N__10663));
    Odrv12 I__1091 (
            .O(N__10677),
            .I(voltage_1_1_sqmuxa));
    LocalMux I__1090 (
            .O(N__10674),
            .I(voltage_1_1_sqmuxa));
    LocalMux I__1089 (
            .O(N__10671),
            .I(voltage_1_1_sqmuxa));
    LocalMux I__1088 (
            .O(N__10666),
            .I(voltage_1_1_sqmuxa));
    LocalMux I__1087 (
            .O(N__10663),
            .I(voltage_1_1_sqmuxa));
    InMux I__1086 (
            .O(N__10652),
            .I(N__10649));
    LocalMux I__1085 (
            .O(N__10649),
            .I(N__10646));
    Odrv4 I__1084 (
            .O(N__10646),
            .I(voltage_3_RNO_0Z0Z_2));
    CascadeMux I__1083 (
            .O(N__10643),
            .I(voltage_3_9_iv_0_2_cascade_));
    CascadeMux I__1082 (
            .O(N__10640),
            .I(CO2_3_cascade_));
    CascadeMux I__1081 (
            .O(N__10637),
            .I(N_1155_cascade_));
    InMux I__1080 (
            .O(N__10634),
            .I(N__10631));
    LocalMux I__1079 (
            .O(N__10631),
            .I(voltage_0_10_iv_0_3));
    InMux I__1078 (
            .O(N__10628),
            .I(N__10624));
    InMux I__1077 (
            .O(N__10627),
            .I(N__10621));
    LocalMux I__1076 (
            .O(N__10624),
            .I(N_1519));
    LocalMux I__1075 (
            .O(N__10621),
            .I(N_1519));
    InMux I__1074 (
            .O(N__10616),
            .I(N__10613));
    LocalMux I__1073 (
            .O(N__10613),
            .I(if_generate_plus_mult1_un68_sum_axbxc5_x0));
    CascadeMux I__1072 (
            .O(N__10610),
            .I(if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_));
    InMux I__1071 (
            .O(N__10607),
            .I(N__10598));
    InMux I__1070 (
            .O(N__10606),
            .I(N__10598));
    InMux I__1069 (
            .O(N__10605),
            .I(N__10591));
    InMux I__1068 (
            .O(N__10604),
            .I(N__10591));
    InMux I__1067 (
            .O(N__10603),
            .I(N__10591));
    LocalMux I__1066 (
            .O(N__10598),
            .I(N__10586));
    LocalMux I__1065 (
            .O(N__10591),
            .I(N__10586));
    Odrv4 I__1064 (
            .O(N__10586),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8));
    InMux I__1063 (
            .O(N__10583),
            .I(N__10580));
    LocalMux I__1062 (
            .O(N__10580),
            .I(if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0));
    CascadeMux I__1061 (
            .O(N__10577),
            .I(if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_));
    InMux I__1060 (
            .O(N__10574),
            .I(N__10568));
    InMux I__1059 (
            .O(N__10573),
            .I(N__10565));
    InMux I__1058 (
            .O(N__10572),
            .I(N__10560));
    InMux I__1057 (
            .O(N__10571),
            .I(N__10560));
    LocalMux I__1056 (
            .O(N__10568),
            .I(beamY_RNI75QM4Z0Z_5));
    LocalMux I__1055 (
            .O(N__10565),
            .I(beamY_RNI75QM4Z0Z_5));
    LocalMux I__1054 (
            .O(N__10560),
            .I(beamY_RNI75QM4Z0Z_5));
    CascadeMux I__1053 (
            .O(N__10553),
            .I(voltage_0_10_iv_0_2_cascade_));
    InMux I__1052 (
            .O(N__10550),
            .I(N__10547));
    LocalMux I__1051 (
            .O(N__10547),
            .I(voltage_0_RNO_0Z0Z_2));
    CascadeMux I__1050 (
            .O(N__10544),
            .I(voltage_1_9_iv_0_2_cascade_));
    CascadeMux I__1049 (
            .O(N__10541),
            .I(beamY_RNI9425Z0Z_6_cascade_));
    InMux I__1048 (
            .O(N__10538),
            .I(N__10535));
    LocalMux I__1047 (
            .O(N__10535),
            .I(if_generate_plus_mult1_un61_sum_ac0_x0));
    InMux I__1046 (
            .O(N__10532),
            .I(N__10529));
    LocalMux I__1045 (
            .O(N__10529),
            .I(if_generate_plus_mult1_un61_sum_ac0_x1));
    InMux I__1044 (
            .O(N__10526),
            .I(N__10523));
    LocalMux I__1043 (
            .O(N__10523),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0_6));
    InMux I__1042 (
            .O(N__10520),
            .I(N__10517));
    LocalMux I__1041 (
            .O(N__10517),
            .I(N__10514));
    Odrv4 I__1040 (
            .O(N__10514),
            .I(row_1_if_generate_plus_mult1_un61_sum_c4_d));
    CascadeMux I__1039 (
            .O(N__10511),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_));
    CascadeMux I__1038 (
            .O(N__10508),
            .I(beamY_RNI75QM4Z0Z_5_cascade_));
    InMux I__1037 (
            .O(N__10505),
            .I(N__10502));
    LocalMux I__1036 (
            .O(N__10502),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz));
    CascadeMux I__1035 (
            .O(N__10499),
            .I(chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_));
    CascadeMux I__1034 (
            .O(N__10496),
            .I(beamY_RNI9425_0Z0Z_6_cascade_));
    CascadeMux I__1033 (
            .O(N__10493),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_));
    CascadeMux I__1032 (
            .O(N__10490),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_));
    InMux I__1031 (
            .O(N__10487),
            .I(N__10484));
    LocalMux I__1030 (
            .O(N__10484),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__1029 (
            .O(N__10481),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__1028 (
            .O(N__10478),
            .I(N__10475));
    InMux I__1027 (
            .O(N__10475),
            .I(N__10472));
    LocalMux I__1026 (
            .O(N__10472),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0));
    CascadeMux I__1025 (
            .O(N__10469),
            .I(un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_));
    CascadeMux I__1024 (
            .O(N__10466),
            .I(un5_visibley_axbxc7_1_cascade_));
    CascadeMux I__1023 (
            .O(N__10463),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3_cascade_));
    InMux I__1022 (
            .O(N__10460),
            .I(N__10457));
    LocalMux I__1021 (
            .O(N__10457),
            .I(N__10454));
    Odrv12 I__1020 (
            .O(N__10454),
            .I(N_41_i));
    CascadeMux I__1019 (
            .O(N__10451),
            .I(N_41_i_cascade_));
    InMux I__1018 (
            .O(N__10448),
            .I(N__10443));
    InMux I__1017 (
            .O(N__10447),
            .I(N__10438));
    InMux I__1016 (
            .O(N__10446),
            .I(N__10438));
    LocalMux I__1015 (
            .O(N__10443),
            .I(N__10427));
    LocalMux I__1014 (
            .O(N__10438),
            .I(N__10427));
    InMux I__1013 (
            .O(N__10437),
            .I(N__10422));
    InMux I__1012 (
            .O(N__10436),
            .I(N__10422));
    InMux I__1011 (
            .O(N__10435),
            .I(N__10415));
    InMux I__1010 (
            .O(N__10434),
            .I(N__10415));
    InMux I__1009 (
            .O(N__10433),
            .I(N__10415));
    InMux I__1008 (
            .O(N__10432),
            .I(N__10412));
    Odrv12 I__1007 (
            .O(N__10427),
            .I(voltage_0_1_sqmuxa));
    LocalMux I__1006 (
            .O(N__10422),
            .I(voltage_0_1_sqmuxa));
    LocalMux I__1005 (
            .O(N__10415),
            .I(voltage_0_1_sqmuxa));
    LocalMux I__1004 (
            .O(N__10412),
            .I(voltage_0_1_sqmuxa));
    InMux I__1003 (
            .O(N__10403),
            .I(N__10400));
    LocalMux I__1002 (
            .O(N__10400),
            .I(ScreenBuffer_0_1_1_sqmuxa_2));
    InMux I__1001 (
            .O(N__10397),
            .I(N__10394));
    LocalMux I__1000 (
            .O(N__10394),
            .I(N__10391));
    Span4Mux_v I__999 (
            .O(N__10391),
            .I(N__10388));
    Odrv4 I__998 (
            .O(N__10388),
            .I(un4_voltage_2_0__i2_mux));
    InMux I__997 (
            .O(N__10385),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__996 (
            .O(N__10382),
            .I(N__10379));
    LocalMux I__995 (
            .O(N__10379),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31));
    InMux I__994 (
            .O(N__10376),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__993 (
            .O(N__10373),
            .I(N__10369));
    InMux I__992 (
            .O(N__10372),
            .I(N__10360));
    InMux I__991 (
            .O(N__10369),
            .I(N__10360));
    InMux I__990 (
            .O(N__10368),
            .I(N__10360));
    InMux I__989 (
            .O(N__10367),
            .I(N__10357));
    LocalMux I__988 (
            .O(N__10360),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1));
    LocalMux I__987 (
            .O(N__10357),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1));
    CascadeMux I__986 (
            .O(N__10352),
            .I(N__10349));
    InMux I__985 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__984 (
            .O(N__10346),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1));
    InMux I__983 (
            .O(N__10343),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__982 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__981 (
            .O(N__10337),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33));
    CascadeMux I__980 (
            .O(N__10334),
            .I(N__10330));
    InMux I__979 (
            .O(N__10333),
            .I(N__10327));
    InMux I__978 (
            .O(N__10330),
            .I(N__10324));
    LocalMux I__977 (
            .O(N__10327),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1));
    LocalMux I__976 (
            .O(N__10324),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1));
    InMux I__975 (
            .O(N__10319),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    CascadeMux I__974 (
            .O(N__10316),
            .I(un4_voltage_10_9__N_4_cascade_));
    InMux I__973 (
            .O(N__10313),
            .I(N__10310));
    LocalMux I__972 (
            .O(N__10310),
            .I(N__10306));
    InMux I__971 (
            .O(N__10309),
            .I(N__10303));
    Odrv12 I__970 (
            .O(N__10306),
            .I(un4_voltage_2_0__N_5_iZ0));
    LocalMux I__969 (
            .O(N__10303),
            .I(un4_voltage_2_0__N_5_iZ0));
    CascadeMux I__968 (
            .O(N__10298),
            .I(voltage_0_1_sqmuxa_cascade_));
    CascadeMux I__967 (
            .O(N__10295),
            .I(N__10292));
    InMux I__966 (
            .O(N__10292),
            .I(N__10289));
    LocalMux I__965 (
            .O(N__10289),
            .I(N__10286));
    Span4Mux_v I__964 (
            .O(N__10286),
            .I(N__10283));
    Odrv4 I__963 (
            .O(N__10283),
            .I(un1_voltage_0_cry_0_0_c_RNOZ0));
    InMux I__962 (
            .O(N__10280),
            .I(N__10277));
    LocalMux I__961 (
            .O(N__10277),
            .I(N_34_0_i));
    InMux I__960 (
            .O(N__10274),
            .I(un1_voltage_3_1_cry_1));
    InMux I__959 (
            .O(N__10271),
            .I(un1_voltage_3_1_cry_2));
    CascadeMux I__958 (
            .O(N__10268),
            .I(N__10264));
    InMux I__957 (
            .O(N__10267),
            .I(N__10261));
    InMux I__956 (
            .O(N__10264),
            .I(N__10258));
    LocalMux I__955 (
            .O(N__10261),
            .I(ScreenBuffer_0_0_1_sqmuxa));
    LocalMux I__954 (
            .O(N__10258),
            .I(ScreenBuffer_0_0_1_sqmuxa));
    CascadeMux I__953 (
            .O(N__10253),
            .I(un4_voltage_2_0__N_13_mux_iZ0_cascade_));
    CascadeMux I__952 (
            .O(N__10250),
            .I(N__10247));
    InMux I__951 (
            .O(N__10247),
            .I(N__10244));
    LocalMux I__950 (
            .O(N__10244),
            .I(N__10241));
    Odrv12 I__949 (
            .O(N__10241),
            .I(SDATA1_ibuf_RNI098KZ0Z2));
    CascadeMux I__948 (
            .O(N__10238),
            .I(N_35_0_i_cascade_));
    CascadeMux I__947 (
            .O(N__10235),
            .I(un1_voltage_1_1_axb_0_cascade_));
    CascadeMux I__946 (
            .O(N__10232),
            .I(voltage_0_1_sqmuxa_1_cascade_));
    CascadeMux I__945 (
            .O(N__10229),
            .I(voltage_3_9_iv_0_0_cascade_));
    InMux I__944 (
            .O(N__10226),
            .I(N__10222));
    InMux I__943 (
            .O(N__10225),
            .I(N__10219));
    LocalMux I__942 (
            .O(N__10222),
            .I(N_1507));
    LocalMux I__941 (
            .O(N__10219),
            .I(N_1507));
    CascadeMux I__940 (
            .O(N__10214),
            .I(N_1507_cascade_));
    InMux I__939 (
            .O(N__10211),
            .I(N__10208));
    LocalMux I__938 (
            .O(N__10208),
            .I(voltage_3_RNO_0Z0Z_0));
    InMux I__937 (
            .O(N__10205),
            .I(un1_voltage_3_1_cry_0));
    InMux I__936 (
            .O(N__10202),
            .I(un1_voltage_0_cry_2));
    CascadeMux I__935 (
            .O(N__10199),
            .I(N_1503_cascade_));
    InMux I__934 (
            .O(N__10196),
            .I(N__10193));
    LocalMux I__933 (
            .O(N__10193),
            .I(SDATA1_ibuf_RNILOUGZ0Z2));
    InMux I__932 (
            .O(N__10190),
            .I(N__10187));
    LocalMux I__931 (
            .O(N__10187),
            .I(if_generate_plus_mult1_un75_sum_axbxc5_0_x1));
    CascadeMux I__930 (
            .O(N__10184),
            .I(if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_));
    CascadeMux I__929 (
            .O(N__10181),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_));
    InMux I__928 (
            .O(N__10178),
            .I(un1_voltage_0_cry_0));
    InMux I__927 (
            .O(N__10175),
            .I(un1_voltage_0_cry_1));
    InMux I__926 (
            .O(N__10172),
            .I(un20_beamy_cry_1));
    InMux I__925 (
            .O(N__10169),
            .I(un20_beamy_cry_2));
    InMux I__924 (
            .O(N__10166),
            .I(un20_beamy_cry_3));
    InMux I__923 (
            .O(N__10163),
            .I(un20_beamy_cry_4));
    InMux I__922 (
            .O(N__10160),
            .I(un20_beamy_cry_5));
    InMux I__921 (
            .O(N__10157),
            .I(un20_beamy_cry_6));
    InMux I__920 (
            .O(N__10154),
            .I(un20_beamy_cry_7));
    InMux I__919 (
            .O(N__10151),
            .I(bfn_1_7_0_));
    InMux I__918 (
            .O(N__10148),
            .I(N__10145));
    LocalMux I__917 (
            .O(N__10145),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0));
    InMux I__916 (
            .O(N__10142),
            .I(N__10139));
    LocalMux I__915 (
            .O(N__10139),
            .I(beamY_RNISI4A_0Z0Z_9));
    CascadeMux I__914 (
            .O(N__10136),
            .I(beamY_RNIE925Z0Z_6_cascade_));
    InMux I__913 (
            .O(N__10133),
            .I(N__10130));
    LocalMux I__912 (
            .O(N__10130),
            .I(beamY_RNIKOP3_0Z0Z_6));
    CascadeMux I__911 (
            .O(N__10127),
            .I(un5_visibley_c2_cascade_));
    CascadeMux I__910 (
            .O(N__10124),
            .I(N__10120));
    InMux I__909 (
            .O(N__10123),
            .I(N__10117));
    InMux I__908 (
            .O(N__10120),
            .I(N__10114));
    LocalMux I__907 (
            .O(N__10117),
            .I(un5_visibley_c6_0_0_0));
    LocalMux I__906 (
            .O(N__10114),
            .I(un5_visibley_c6_0_0_0));
    InMux I__905 (
            .O(N__10109),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__904 (
            .O(N__10106),
            .I(N__10097));
    InMux I__903 (
            .O(N__10105),
            .I(N__10097));
    InMux I__902 (
            .O(N__10104),
            .I(N__10090));
    InMux I__901 (
            .O(N__10103),
            .I(N__10090));
    InMux I__900 (
            .O(N__10102),
            .I(N__10090));
    LocalMux I__899 (
            .O(N__10097),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0));
    LocalMux I__898 (
            .O(N__10090),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0));
    CascadeMux I__897 (
            .O(N__10085),
            .I(N__10082));
    InMux I__896 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__895 (
            .O(N__10079),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__894 (
            .O(N__10076),
            .I(N__10071));
    InMux I__893 (
            .O(N__10075),
            .I(N__10066));
    InMux I__892 (
            .O(N__10074),
            .I(N__10066));
    LocalMux I__891 (
            .O(N__10071),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__890 (
            .O(N__10066),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    CascadeMux I__889 (
            .O(N__10061),
            .I(N__10058));
    InMux I__888 (
            .O(N__10058),
            .I(N__10055));
    LocalMux I__887 (
            .O(N__10055),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0));
    InMux I__886 (
            .O(N__10052),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__885 (
            .O(N__10049),
            .I(N__10046));
    LocalMux I__884 (
            .O(N__10046),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0));
    InMux I__883 (
            .O(N__10043),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__882 (
            .O(N__10040),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__881 (
            .O(N__10037),
            .I(N__10031));
    InMux I__880 (
            .O(N__10036),
            .I(N__10031));
    LocalMux I__879 (
            .O(N__10031),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__878 (
            .O(N__10028),
            .I(N__10025));
    LocalMux I__877 (
            .O(N__10025),
            .I(beamY_RNITSR8_0Z0Z_8));
    InMux I__876 (
            .O(N__10022),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__875 (
            .O(N__10019),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__874 (
            .O(N__10016),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_));
    CascadeMux I__873 (
            .O(N__10013),
            .I(N__10010));
    InMux I__872 (
            .O(N__10010),
            .I(N__10007));
    LocalMux I__871 (
            .O(N__10007),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7));
    CascadeMux I__870 (
            .O(N__10004),
            .I(N__10001));
    InMux I__869 (
            .O(N__10001),
            .I(N__9998));
    LocalMux I__868 (
            .O(N__9998),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0));
    InMux I__867 (
            .O(N__9995),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__866 (
            .O(N__9992),
            .I(N__9989));
    InMux I__865 (
            .O(N__9989),
            .I(N__9986));
    LocalMux I__864 (
            .O(N__9986),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0));
    InMux I__863 (
            .O(N__9983),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__862 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__861 (
            .O(N__9977),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0));
    InMux I__860 (
            .O(N__9974),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__859 (
            .O(N__9971),
            .I(N__9968));
    InMux I__858 (
            .O(N__9968),
            .I(N__9965));
    LocalMux I__857 (
            .O(N__9965),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__856 (
            .O(N__9962),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    IoInMux I__855 (
            .O(N__9959),
            .I(N__9956));
    LocalMux I__854 (
            .O(N__9956),
            .I(N__9953));
    IoSpan4Mux I__853 (
            .O(N__9953),
            .I(N__9950));
    IoSpan4Mux I__852 (
            .O(N__9950),
            .I(N__9947));
    IoSpan4Mux I__851 (
            .O(N__9947),
            .I(N__9944));
    Odrv4 I__850 (
            .O(N__9944),
            .I(\Clock50MHz.PixelClock ));
    InMux I__849 (
            .O(N__9941),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__848 (
            .O(N__9938),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__847 (
            .O(N__9935),
            .I(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(un20_beamy_cry_8),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(counter_cry_8),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_2_0_));
    defparam IN_MUX_bfv_4_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_1_0_));
    defparam IN_MUX_bfv_2_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_1_0_));
    defparam IN_MUX_bfv_1_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_1_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    ICE_GB slaveselect_RNIO5RB1_0 (
            .USERSIGNALTOGLOBALBUFFER(N__11612),
            .GLOBALBUFFEROUTPUT(voltage_0_0_sqmuxa_1_g));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__9959),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_1_1_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_1_1_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_1_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_1_1_0 (
            .in0(_gnd_net_),
            .in1(N__12688),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_1_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01J31_LC_1_1_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01J31_LC_1_1_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01J31_LC_1_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01J31_LC_1_1_1 (
            .in0(_gnd_net_),
            .in1(N__10103),
            .in2(N__10085),
            .in3(N__9941),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQI1_LC_1_1_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQI1_LC_1_1_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQI1_LC_1_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQI1_LC_1_1_2 (
            .in0(_gnd_net_),
            .in1(N__10105),
            .in2(N__10004),
            .in3(N__9938),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9P1_LC_1_1_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9P1_LC_1_1_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9P1_LC_1_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9P1_LC_1_1_3 (
            .in0(_gnd_net_),
            .in1(N__10104),
            .in2(N__9992),
            .in3(N__9935),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI8SH33_LC_1_1_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI8SH33_LC_1_1_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI8SH33_LC_1_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI8SH33_LC_1_1_4 (
            .in0(N__10367),
            .in1(N__9980),
            .in2(N__10013),
            .in3(N__10022),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25A1_LC_1_1_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25A1_LC_1_1_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25A1_LC_1_1_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25A1_LC_1_1_5 (
            .in0(N__10106),
            .in1(N__10076),
            .in2(N__9971),
            .in3(N__10019),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1),
            .ltout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5ME33_LC_1_1_6.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5ME33_LC_1_1_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5ME33_LC_1_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5ME33_LC_1_1_6 (
            .in0(N__10333),
            .in1(_gnd_net_),
            .in2(N__10016),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_0_LC_1_1_7.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_0_LC_1_1_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_0_LC_1_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_0_LC_1_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10102),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_2_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_2_0 (
            .in0(_gnd_net_),
            .in1(N__14002),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7K_LC_1_2_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7K_LC_1_2_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7K_LC_1_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7K_LC_1_2_1 (
            .in0(_gnd_net_),
            .in1(N__10028),
            .in2(N__21913),
            .in3(N__9995),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQ_LC_1_2_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQ_LC_1_2_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQ_LC_1_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQ_LC_1_2_2 (
            .in0(_gnd_net_),
            .in1(N__21908),
            .in2(N__10061),
            .in3(N__9983),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQ_LC_1_2_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQ_LC_1_2_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQ_LC_1_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQ_LC_1_2_3 (
            .in0(_gnd_net_),
            .in1(N__10049),
            .in2(N__21914),
            .in3(N__9974),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_1_2_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_1_2_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_1_2_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_1_2_4 (
            .in0(_gnd_net_),
            .in1(N__10074),
            .in2(_gnd_net_),
            .in3(N__9962),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_LC_1_2_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_LC_1_2_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_LC_1_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_LC_1_2_5 (
            .in0(_gnd_net_),
            .in1(N__10037),
            .in2(_gnd_net_),
            .in3(N__10109),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_2_6.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_2_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14003),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_1_2_7.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_1_2_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_1_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_1_2_7 (
            .in0(N__10075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10036),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_3_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_3_0 (
            .in0(_gnd_net_),
            .in1(N__10148),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8F_LC_1_3_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8F_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8F_LC_1_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8F_LC_1_3_1 (
            .in0(_gnd_net_),
            .in1(N__10142),
            .in2(N__21887),
            .in3(N__10052),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9F_LC_1_3_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9F_LC_1_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9F_LC_1_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9F_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(N__21866),
            .in2(N__18283),
            .in3(N__10043),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_1_3_3.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_1_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_1_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_1_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10040),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITSR8_0_8_LC_1_3_5.C_ON=1'b0;
    defparam beamY_RNITSR8_0_8_LC_1_3_5.SEQ_MODE=4'b0000;
    defparam beamY_RNITSR8_0_8_LC_1_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNITSR8_0_8_LC_1_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18157),
            .lcout(beamY_RNITSR8_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_1_4_2.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_1_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_1_4_2.LUT_INIT=16'b1100100111000011;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_1_4_2 (
            .in0(N__14661),
            .in1(N__14891),
            .in2(N__10124),
            .in3(N__11247),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_0_9_LC_1_4_6.C_ON=1'b0;
    defparam beamY_RNISI4A_0_9_LC_1_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_0_9_LC_1_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNISI4A_0_9_LC_1_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18225),
            .lcout(beamY_RNISI4A_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIE925_6_LC_1_5_0.C_ON=1'b0;
    defparam beamY_RNIE925_6_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIE925_6_LC_1_5_0.LUT_INIT=16'b1010101010101001;
    LogicCell40 beamY_RNIE925_6_LC_1_5_0 (
            .in0(N__14782),
            .in1(N__12972),
            .in2(N__14658),
            .in3(N__12881),
            .lcout(),
            .ltout(beamY_RNIE925Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0DB_6_LC_1_5_1.C_ON=1'b0;
    defparam beamY_RNIJ0DB_6_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0DB_6_LC_1_5_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 beamY_RNIJ0DB_6_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__10133),
            .in2(N__10136),
            .in3(N__11248),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKOP3_0_6_LC_1_5_2.C_ON=1'b0;
    defparam beamY_RNIKOP3_0_6_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIKOP3_0_6_LC_1_5_2.LUT_INIT=16'b1010101010011001;
    LogicCell40 beamY_RNIKOP3_0_6_LC_1_5_2 (
            .in0(N__14781),
            .in1(N__12971),
            .in2(_gnd_net_),
            .in3(N__12880),
            .lcout(beamY_RNIKOP3_0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_1_5_4.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_1_5_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_RNIHUG2_3_LC_1_5_4 (
            .in0(_gnd_net_),
            .in1(N__20751),
            .in2(_gnd_net_),
            .in3(N__14417),
            .lcout(un5_visibley_c2),
            .ltout(un5_visibley_c2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITSR8_8_LC_1_5_5.C_ON=1'b0;
    defparam beamY_RNITSR8_8_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNITSR8_8_LC_1_5_5.LUT_INIT=16'b1110101000010101;
    LogicCell40 beamY_RNITSR8_8_LC_1_5_5 (
            .in0(N__10123),
            .in1(N__14617),
            .in2(N__10127),
            .in3(N__14877),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKOP3_6_LC_1_5_6.C_ON=1'b0;
    defparam beamY_RNIKOP3_6_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIKOP3_6_LC_1_5_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamY_RNIKOP3_6_LC_1_5_6 (
            .in0(N__14780),
            .in1(N__12970),
            .in2(_gnd_net_),
            .in3(N__12879),
            .lcout(un5_visibley_c6_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_3_LC_1_5_7.C_ON=1'b0;
    defparam beamY_RNIBFP3_3_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_3_LC_1_5_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 beamY_RNIBFP3_3_LC_1_5_7 (
            .in0(N__20752),
            .in1(N__14621),
            .in2(_gnd_net_),
            .in3(N__14421),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_1_c_LC_1_6_0.C_ON=1'b1;
    defparam un20_beamy_cry_1_c_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_1_c_LC_1_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un20_beamy_cry_1_c_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(N__23301),
            .in2(N__24859),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(un20_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_1_6_1.C_ON=1'b1;
    defparam beamY_2_LC_1_6_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_1_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_2_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(N__20789),
            .in2(_gnd_net_),
            .in3(N__10172),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(un20_beamy_cry_1),
            .carryout(un20_beamy_cry_2),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_3_LC_1_6_2.C_ON=1'b1;
    defparam beamY_3_LC_1_6_2.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_1_6_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_3_LC_1_6_2 (
            .in0(N__14146),
            .in1(N__14440),
            .in2(_gnd_net_),
            .in3(N__10169),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(un20_beamy_cry_2),
            .carryout(un20_beamy_cry_3),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_4_LC_1_6_3.C_ON=1'b1;
    defparam beamY_4_LC_1_6_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_1_6_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_4_LC_1_6_3 (
            .in0(N__14145),
            .in1(N__14657),
            .in2(_gnd_net_),
            .in3(N__10166),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un20_beamy_cry_3),
            .carryout(un20_beamy_cry_4),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_5_LC_1_6_4.C_ON=1'b1;
    defparam beamY_5_LC_1_6_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_1_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_1_6_4 (
            .in0(_gnd_net_),
            .in1(N__12898),
            .in2(_gnd_net_),
            .in3(N__10163),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un20_beamy_cry_4),
            .carryout(un20_beamy_cry_5),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_6_LC_1_6_5.C_ON=1'b1;
    defparam beamY_6_LC_1_6_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_1_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(N__12988),
            .in2(_gnd_net_),
            .in3(N__10160),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un20_beamy_cry_5),
            .carryout(un20_beamy_cry_6),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_7_LC_1_6_6.C_ON=1'b1;
    defparam beamY_7_LC_1_6_6.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_1_6_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_7_LC_1_6_6 (
            .in0(N__14147),
            .in1(N__14809),
            .in2(_gnd_net_),
            .in3(N__10157),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(un20_beamy_cry_6),
            .carryout(un20_beamy_cry_7),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_8_LC_1_6_7.C_ON=1'b1;
    defparam beamY_8_LC_1_6_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_1_6_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_1_6_7 (
            .in0(_gnd_net_),
            .in1(N__14889),
            .in2(_gnd_net_),
            .in3(N__10154),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un20_beamy_cry_7),
            .carryout(un20_beamy_cry_8),
            .clk(N__21053),
            .ce(N__17541),
            .sr(_gnd_net_));
    defparam beamY_9_LC_1_7_0.C_ON=1'b0;
    defparam beamY_9_LC_1_7_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_1_7_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_1_7_0 (
            .in0(N__14972),
            .in1(N__14144),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21052),
            .ce(N__17546),
            .sr(_gnd_net_));
    defparam beamY_RNICE3U5_5_LC_1_8_0.C_ON=1'b0;
    defparam beamY_RNICE3U5_5_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam beamY_RNICE3U5_5_LC_1_8_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 beamY_RNICE3U5_5_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(N__10604),
            .in2(_gnd_net_),
            .in3(N__10573),
            .lcout(r_N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x1_LC_1_8_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x1_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x1_LC_1_8_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x1_LC_1_8_1 (
            .in0(N__12292),
            .in1(N__14519),
            .in2(N__12457),
            .in3(N__11530),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc5_0_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x0_LC_1_8_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x0_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x0_LC_1_8_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x0_LC_1_8_3 (
            .in0(N__12293),
            .in1(N__14520),
            .in2(N__12458),
            .in3(N__11529),
            .lcout(),
            .ltout(if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_ns_LC_1_8_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_ns_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_ns_LC_1_8_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_ns_LC_1_8_4 (
            .in0(_gnd_net_),
            .in1(N__10190),
            .in2(N__10184),
            .in3(N__11560),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0_LC_1_8_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0_LC_1_8_5.LUT_INIT=16'b0000101011101000;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0_LC_1_8_5 (
            .in0(N__10603),
            .in1(N__13211),
            .in2(N__12456),
            .in3(N__14517),
            .lcout(if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_1_8_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_1_8_6.LUT_INIT=16'b1111111110001000;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_c4_LC_1_8_6 (
            .in0(N__14518),
            .in1(N__12415),
            .in2(_gnd_net_),
            .in3(N__10526),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x0_LC_1_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x0_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x0_LC_1_8_7.LUT_INIT=16'b1110000100011110;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_x0_LC_1_8_7 (
            .in0(N__10605),
            .in1(N__10574),
            .in2(N__10181),
            .in3(N__11528),
            .lcout(if_generate_plus_mult1_un68_sum_axbxc5_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_0_cry_0_0_c_LC_1_9_0.C_ON=1'b1;
    defparam un1_voltage_0_cry_0_0_c_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam un1_voltage_0_cry_0_0_c_LC_1_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_voltage_0_cry_0_0_c_LC_1_9_0 (
            .in0(_gnd_net_),
            .in1(N__18478),
            .in2(N__10295),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(un1_voltage_0_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_0_1_LC_1_9_1.C_ON=1'b1;
    defparam voltage_0_RNO_0_1_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_0_1_LC_1_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_0_RNO_0_1_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(N__19052),
            .in2(N__10250),
            .in3(N__10178),
            .lcout(voltage_0_RNO_0Z0Z_1),
            .ltout(),
            .carryin(un1_voltage_0_cry_0),
            .carryout(un1_voltage_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_0_2_LC_1_9_2.C_ON=1'b1;
    defparam voltage_0_RNO_0_2_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_0_2_LC_1_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_0_RNO_0_2_LC_1_9_2 (
            .in0(_gnd_net_),
            .in1(N__10196),
            .in2(N__16554),
            .in3(N__10175),
            .lcout(voltage_0_RNO_0Z0Z_2),
            .ltout(),
            .carryin(un1_voltage_0_cry_1),
            .carryout(un1_voltage_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_3_LC_1_9_3.C_ON=1'b0;
    defparam voltage_0_3_LC_1_9_3.SEQ_MODE=4'b1000;
    defparam voltage_0_3_LC_1_9_3.LUT_INIT=16'b0101011101011101;
    LogicCell40 voltage_0_3_LC_1_9_3 (
            .in0(N__10634),
            .in1(N__19412),
            .in2(N__17983),
            .in3(N__10202),
            .lcout(voltage_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19953),
            .ce(),
            .sr(N__18541));
    defparam ScreenBuffer_1_0_e_0_0_LC_1_10_0.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_0_LC_1_10_0.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_0_e_0_0_LC_1_10_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 ScreenBuffer_1_0_e_0_0_LC_1_10_0 (
            .in0(N__19182),
            .in1(N__18505),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(ScreenBuffer_1_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19954),
            .ce(N__18997),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_2_LC_1_10_1.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_2_LC_1_10_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_0_e_0_2_LC_1_10_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 ScreenBuffer_1_0_e_0_2_LC_1_10_1 (
            .in0(N__16584),
            .in1(N__19183),
            .in2(_gnd_net_),
            .in3(N__16544),
            .lcout(ScreenBuffer_1_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19954),
            .ce(N__18997),
            .sr(_gnd_net_));
    defparam voltage_0_RNITQ2M_0_LC_1_10_2.C_ON=1'b0;
    defparam voltage_0_RNITQ2M_0_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam voltage_0_RNITQ2M_0_LC_1_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 voltage_0_RNITQ2M_0_LC_1_10_2 (
            .in0(N__15391),
            .in1(N__18480),
            .in2(_gnd_net_),
            .in3(N__15720),
            .lcout(),
            .ltout(N_1503_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI49LH1_0_0_LC_1_10_3.C_ON=1'b0;
    defparam counter_RNI49LH1_0_0_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam counter_RNI49LH1_0_0_LC_1_10_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 counter_RNI49LH1_0_0_LC_1_10_3 (
            .in0(_gnd_net_),
            .in1(N__16277),
            .in2(N__10199),
            .in3(N__10225),
            .lcout(counter_RNI49LH1_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNITQ2M_0_0_LC_1_10_4.C_ON=1'b0;
    defparam voltage_0_RNITQ2M_0_0_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam voltage_0_RNITQ2M_0_0_LC_1_10_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 voltage_0_RNITQ2M_0_0_LC_1_10_4 (
            .in0(N__15390),
            .in1(N__18479),
            .in2(_gnd_net_),
            .in3(N__15718),
            .lcout(N_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNI1V2M_0_2_LC_1_10_5.C_ON=1'b0;
    defparam voltage_0_RNI1V2M_0_2_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam voltage_0_RNI1V2M_0_2_LC_1_10_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 voltage_0_RNI1V2M_0_2_LC_1_10_5 (
            .in0(N__15719),
            .in1(N__15301),
            .in2(_gnd_net_),
            .in3(N__16543),
            .lcout(N_1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_0_0_LC_1_10_6.C_ON=1'b0;
    defparam voltage_0_RNO_0_0_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_0_0_LC_1_10_6.LUT_INIT=16'b0111011110001000;
    LogicCell40 voltage_0_RNO_0_0_LC_1_10_6 (
            .in0(N__10447),
            .in1(N__10313),
            .in2(_gnd_net_),
            .in3(N__18481),
            .lcout(un1_voltage_0_axb_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATA1_ibuf_RNILOUG2_LC_1_10_7.C_ON=1'b0;
    defparam SDATA1_ibuf_RNILOUG2_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam SDATA1_ibuf_RNILOUG2_LC_1_10_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 SDATA1_ibuf_RNILOUG2_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(N__10397),
            .in2(_gnd_net_),
            .in3(N__10446),
            .lcout(SDATA1_ibuf_RNILOUGZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI2ACM1_0_0_LC_1_11_0.C_ON=1'b0;
    defparam counter_RNI2ACM1_0_0_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam counter_RNI2ACM1_0_0_LC_1_11_0.LUT_INIT=16'b0001000000000000;
    LogicCell40 counter_RNI2ACM1_0_0_LC_1_11_0 (
            .in0(N__19180),
            .in1(N__16251),
            .in2(N__13349),
            .in3(N__15739),
            .lcout(voltage_3_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_0_0_LC_1_11_1.C_ON=1'b0;
    defparam voltage_1_RNO_0_0_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_0_0_LC_1_11_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 voltage_1_RNO_0_0_LC_1_11_1 (
            .in0(N__10460),
            .in1(N__15329),
            .in2(_gnd_net_),
            .in3(N__10448),
            .lcout(),
            .ltout(un1_voltage_1_1_axb_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_0_LC_1_11_2.C_ON=1'b0;
    defparam voltage_1_0_LC_1_11_2.SEQ_MODE=4'b1000;
    defparam voltage_1_0_LC_1_11_2.LUT_INIT=16'b1111010111010101;
    LogicCell40 voltage_1_0_LC_1_11_2 (
            .in0(N__10733),
            .in1(N__11862),
            .in2(N__10235),
            .in3(N__15740),
            .lcout(voltage_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19956),
            .ce(),
            .sr(N__18543));
    defparam counter_RNI2ACM1_0_LC_1_11_3.C_ON=1'b0;
    defparam counter_RNI2ACM1_0_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam counter_RNI2ACM1_0_LC_1_11_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 counter_RNI2ACM1_0_LC_1_11_3 (
            .in0(N__16250),
            .in1(N__19179),
            .in2(N__15811),
            .in3(N__13343),
            .lcout(voltage_0_1_sqmuxa_1),
            .ltout(voltage_0_1_sqmuxa_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_1_0_LC_1_11_4.C_ON=1'b0;
    defparam voltage_3_RNO_1_0_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_1_0_LC_1_11_4.LUT_INIT=16'b0101111100010011;
    LogicCell40 voltage_3_RNO_1_0_LC_1_11_4 (
            .in0(N__10226),
            .in1(N__11921),
            .in2(N__10232),
            .in3(N__12038),
            .lcout(),
            .ltout(voltage_3_9_iv_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_0_LC_1_11_5.C_ON=1'b0;
    defparam voltage_3_0_LC_1_11_5.SEQ_MODE=4'b1000;
    defparam voltage_3_0_LC_1_11_5.LUT_INIT=16'b1000111111001111;
    LogicCell40 voltage_3_0_LC_1_11_5 (
            .in0(N__11861),
            .in1(N__10211),
            .in2(N__10229),
            .in3(N__15814),
            .lcout(voltage_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19956),
            .ce(),
            .sr(N__18543));
    defparam voltage_1_RNIV09O_0_LC_1_11_6.C_ON=1'b0;
    defparam voltage_1_RNIV09O_0_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam voltage_1_RNIV09O_0_LC_1_11_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 voltage_1_RNIV09O_0_LC_1_11_6 (
            .in0(N__15328),
            .in1(N__18503),
            .in2(_gnd_net_),
            .in3(N__15735),
            .lcout(N_1507),
            .ltout(N_1507_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI49LH1_0_LC_1_11_7.C_ON=1'b0;
    defparam counter_RNI49LH1_0_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam counter_RNI49LH1_0_LC_1_11_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 counter_RNI49LH1_0_LC_1_11_7 (
            .in0(N__16249),
            .in1(_gnd_net_),
            .in2(N__10214),
            .in3(N__10627),
            .lcout(un74_voltage_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_0_0_LC_1_12_0.C_ON=1'b1;
    defparam voltage_3_RNO_0_0_LC_1_12_0.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_0_0_LC_1_12_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 voltage_3_RNO_0_0_LC_1_12_0 (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__10268),
            .in3(N__10267),
            .lcout(voltage_3_RNO_0Z0Z_0),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(un1_voltage_3_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_0_1_LC_1_12_1.C_ON=1'b1;
    defparam voltage_3_RNO_0_1_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_0_1_LC_1_12_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 voltage_3_RNO_0_1_LC_1_12_1 (
            .in0(_gnd_net_),
            .in1(N__19369),
            .in2(_gnd_net_),
            .in3(N__10205),
            .lcout(voltage_3_RNO_0Z0Z_1),
            .ltout(),
            .carryin(un1_voltage_3_1_cry_0),
            .carryout(un1_voltage_3_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_0_2_LC_1_12_2.C_ON=1'b1;
    defparam voltage_3_RNO_0_2_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_0_2_LC_1_12_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 voltage_3_RNO_0_2_LC_1_12_2 (
            .in0(_gnd_net_),
            .in1(N__16585),
            .in2(_gnd_net_),
            .in3(N__10274),
            .lcout(voltage_3_RNO_0Z0Z_2),
            .ltout(),
            .carryin(un1_voltage_3_1_cry_1),
            .carryout(un1_voltage_3_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_0_3_LC_1_12_3.C_ON=1'b0;
    defparam voltage_3_RNO_0_3_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_0_3_LC_1_12_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 voltage_3_RNO_0_3_LC_1_12_3 (
            .in0(_gnd_net_),
            .in1(N__19450),
            .in2(_gnd_net_),
            .in3(N__10271),
            .lcout(voltage_3_RNO_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI4CSO_3_LC_1_12_4.C_ON=1'b0;
    defparam counter_RNI4CSO_3_LC_1_12_4.SEQ_MODE=4'b0000;
    defparam counter_RNI4CSO_3_LC_1_12_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 counter_RNI4CSO_3_LC_1_12_4 (
            .in0(N__16244),
            .in1(N__16407),
            .in2(N__15755),
            .in3(N__15467),
            .lcout(ScreenBuffer_0_0_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIAV5D_4_LC_1_13_1.C_ON=1'b0;
    defparam counter_RNIAV5D_4_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam counter_RNIAV5D_4_LC_1_13_1.LUT_INIT=16'b1000100010101010;
    LogicCell40 counter_RNIAV5D_4_LC_1_13_1 (
            .in0(N__13864),
            .in1(N__16361),
            .in2(_gnd_net_),
            .in3(N__13506),
            .lcout(un3_slaveselectlt9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_voltage_2_0__N_13_mux_i_LC_1_13_3.C_ON=1'b0;
    defparam un4_voltage_2_0__N_13_mux_i_LC_1_13_3.SEQ_MODE=4'b0000;
    defparam un4_voltage_2_0__N_13_mux_i_LC_1_13_3.LUT_INIT=16'b1011011110000100;
    LogicCell40 un4_voltage_2_0__N_13_mux_i_LC_1_13_3 (
            .in0(N__15976),
            .in1(N__10948),
            .in2(N__15754),
            .in3(N__16362),
            .lcout(),
            .ltout(un4_voltage_2_0__N_13_mux_iZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATA1_ibuf_RNI098K2_LC_1_13_4.C_ON=1'b0;
    defparam SDATA1_ibuf_RNI098K2_LC_1_13_4.SEQ_MODE=4'b0000;
    defparam SDATA1_ibuf_RNI098K2_LC_1_13_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 SDATA1_ibuf_RNI098K2_LC_1_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10253),
            .in3(N__10436),
            .lcout(SDATA1_ibuf_RNI098KZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1_LC_1_13_5.C_ON=1'b0;
    defparam counter_1_LC_1_13_5.SEQ_MODE=4'b1000;
    defparam counter_1_LC_1_13_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 counter_1_LC_1_13_5 (
            .in0(N__16269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15688),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19960),
            .ce(),
            .sr(N__12110));
    defparam counter_RNIE8FG_2_LC_1_13_6.C_ON=1'b0;
    defparam counter_RNIE8FG_2_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam counter_RNIE8FG_2_LC_1_13_6.LUT_INIT=16'b0000101000111010;
    LogicCell40 counter_RNIE8FG_2_LC_1_13_6 (
            .in0(N__10949),
            .in1(N__16268),
            .in2(N__15756),
            .in3(N__15977),
            .lcout(),
            .ltout(N_35_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIT58K2_2_LC_1_13_7.C_ON=1'b0;
    defparam counter_RNIT58K2_2_LC_1_13_7.SEQ_MODE=4'b0000;
    defparam counter_RNIT58K2_2_LC_1_13_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 counter_RNIT58K2_2_LC_1_13_7 (
            .in0(N__10437),
            .in1(_gnd_net_),
            .in2(N__10238),
            .in3(_gnd_net_),
            .lcout(counter_RNIT58K2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_voltage_2_0__N_5_i_LC_1_14_0.C_ON=1'b0;
    defparam un4_voltage_2_0__N_5_i_LC_1_14_0.SEQ_MODE=4'b0000;
    defparam un4_voltage_2_0__N_5_i_LC_1_14_0.LUT_INIT=16'b1011101010111110;
    LogicCell40 un4_voltage_2_0__N_5_i_LC_1_14_0 (
            .in0(N__13868),
            .in1(N__16212),
            .in2(N__15997),
            .in3(N__15664),
            .lcout(un4_voltage_2_0__N_5_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_0_3_LC_1_14_1.C_ON=1'b0;
    defparam voltage_2_RNO_0_3_LC_1_14_1.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_0_3_LC_1_14_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 voltage_2_RNO_0_3_LC_1_14_1 (
            .in0(N__10403),
            .in1(N__15205),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(un1_voltage_2_1_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNILOUG2_3_LC_1_14_2.C_ON=1'b0;
    defparam counter_RNILOUG2_3_LC_1_14_2.SEQ_MODE=4'b0000;
    defparam counter_RNILOUG2_3_LC_1_14_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 counter_RNILOUG2_3_LC_1_14_2 (
            .in0(_gnd_net_),
            .in1(N__10280),
            .in2(_gnd_net_),
            .in3(N__10433),
            .lcout(counter_RNILOUG2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI2RBA2_3_LC_1_14_3.C_ON=1'b0;
    defparam counter_RNI2RBA2_3_LC_1_14_3.SEQ_MODE=4'b0000;
    defparam counter_RNI2RBA2_3_LC_1_14_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 counter_RNI2RBA2_3_LC_1_14_3 (
            .in0(N__10435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10947),
            .lcout(counter_RNI2RBA2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_voltage_10_9__m3_LC_1_14_4.C_ON=1'b0;
    defparam un4_voltage_10_9__m3_LC_1_14_4.SEQ_MODE=4'b0000;
    defparam un4_voltage_10_9__m3_LC_1_14_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 un4_voltage_10_9__m3_LC_1_14_4 (
            .in0(N__10946),
            .in1(N__16406),
            .in2(N__15998),
            .in3(N__16273),
            .lcout(),
            .ltout(un4_voltage_10_9__N_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNIKG123_1_LC_1_14_5.C_ON=1'b0;
    defparam voltage_2_RNIKG123_1_LC_1_14_5.SEQ_MODE=4'b0000;
    defparam voltage_2_RNIKG123_1_LC_1_14_5.LUT_INIT=16'b0010000000100000;
    LogicCell40 voltage_2_RNIKG123_1_LC_1_14_5 (
            .in0(N__10434),
            .in1(N__15684),
            .in2(N__10316),
            .in3(N__15146),
            .lcout(voltage_2_RNIKG123Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATA1_ibuf_RNIFTO32_LC_1_14_6.C_ON=1'b0;
    defparam SDATA1_ibuf_RNIFTO32_LC_1_14_6.SEQ_MODE=4'b0000;
    defparam SDATA1_ibuf_RNIFTO32_LC_1_14_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 SDATA1_ibuf_RNIFTO32_LC_1_14_6 (
            .in0(N__19178),
            .in1(N__20217),
            .in2(_gnd_net_),
            .in3(N__16466),
            .lcout(voltage_0_1_sqmuxa),
            .ltout(voltage_0_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_0_cry_0_0_c_RNO_LC_1_14_7.C_ON=1'b0;
    defparam un1_voltage_0_cry_0_0_c_RNO_LC_1_14_7.SEQ_MODE=4'b0000;
    defparam un1_voltage_0_cry_0_0_c_RNO_LC_1_14_7.LUT_INIT=16'b1100000011000000;
    LogicCell40 un1_voltage_0_cry_0_0_c_RNO_LC_1_14_7 (
            .in0(_gnd_net_),
            .in1(N__10309),
            .in2(N__10298),
            .in3(_gnd_net_),
            .lcout(un1_voltage_0_cry_0_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_1_3_LC_1_15_0.C_ON=1'b0;
    defparam counter_RNI6R5D_1_3_LC_1_15_0.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_1_3_LC_1_15_0.LUT_INIT=16'b0011000101000100;
    LogicCell40 counter_RNI6R5D_1_3_LC_1_15_0 (
            .in0(N__16400),
            .in1(N__15989),
            .in2(N__15813),
            .in3(N__16261),
            .lcout(N_34_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNICVT22_LC_1_15_2.C_ON=1'b0;
    defparam slaveselect_RNICVT22_LC_1_15_2.SEQ_MODE=4'b0000;
    defparam slaveselect_RNICVT22_LC_1_15_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 slaveselect_RNICVT22_LC_1_15_2 (
            .in0(_gnd_net_),
            .in1(N__19181),
            .in2(_gnd_net_),
            .in3(N__16482),
            .lcout(un1_sclk17_9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_0_3_LC_1_15_4.C_ON=1'b0;
    defparam counter_RNI6R5D_0_3_LC_1_15_4.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_0_3_LC_1_15_4.LUT_INIT=16'b0101010100111100;
    LogicCell40 counter_RNI6R5D_0_3_LC_1_15_4 (
            .in0(N__16401),
            .in1(N__15988),
            .in2(N__15812),
            .in3(N__16260),
            .lcout(N_41_i),
            .ltout(N_41_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_1_1_cry_0_0_c_RNO_LC_1_15_5.C_ON=1'b0;
    defparam un1_voltage_1_1_cry_0_0_c_RNO_LC_1_15_5.SEQ_MODE=4'b0000;
    defparam un1_voltage_1_1_cry_0_0_c_RNO_LC_1_15_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 un1_voltage_1_1_cry_0_0_c_RNO_LC_1_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10451),
            .in3(N__10432),
            .lcout(un1_voltage_1_1_cry_0_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_2_3_LC_1_15_6.C_ON=1'b0;
    defparam voltage_2_RNO_2_3_LC_1_15_6.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_2_3_LC_1_15_6.LUT_INIT=16'b0000001000000000;
    LogicCell40 voltage_2_RNO_2_3_LC_1_15_6 (
            .in0(N__20195),
            .in1(N__16265),
            .in2(N__16423),
            .in3(N__15750),
            .lcout(ScreenBuffer_0_1_1_sqmuxa_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_voltage_2_0__m11_LC_1_15_7.C_ON=1'b0;
    defparam un4_voltage_2_0__m11_LC_1_15_7.SEQ_MODE=4'b0000;
    defparam un4_voltage_2_0__m11_LC_1_15_7.LUT_INIT=16'b0110000100011000;
    LogicCell40 un4_voltage_2_0__m11_LC_1_15_7 (
            .in0(N__15990),
            .in1(N__15749),
            .in2(N__16284),
            .in3(N__16402),
            .lcout(un4_voltage_2_0__i2_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_1_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_1_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_1_0 (
            .in0(_gnd_net_),
            .in1(N__12472),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_1_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCI1_LC_2_1_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCI1_LC_2_1_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCI1_LC_2_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCI1_LC_2_1_1 (
            .in0(_gnd_net_),
            .in1(N__10368),
            .in2(N__10478),
            .in3(N__10385),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSH2_LC_2_1_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSH2_LC_2_1_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSH2_LC_2_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSH2_LC_2_1_2 (
            .in0(_gnd_net_),
            .in1(N__10382),
            .in2(N__10373),
            .in3(N__10376),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI96513_LC_2_1_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI96513_LC_2_1_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI96513_LC_2_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI96513_LC_2_1_3 (
            .in0(_gnd_net_),
            .in1(N__10372),
            .in2(N__10352),
            .in3(N__10343),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIVCO88_LC_2_1_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIVCO88_LC_2_1_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIVCO88_LC_2_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIVCO88_LC_2_1_4 (
            .in0(N__11032),
            .in1(N__10340),
            .in2(N__10334),
            .in3(N__10319),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_LC_2_1_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_LC_2_1_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_LC_2_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_LC_2_1_5 (
            .in0(_gnd_net_),
            .in1(N__10487),
            .in2(_gnd_net_),
            .in3(N__10481),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_2_1_6.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_2_1_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_2_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_2_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12473),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_2_0.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_2_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12689),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un1_beamylto9_0_LC_2_4_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un1_beamylto9_0_LC_2_4_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un1_beamylto9_0_LC_2_4_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 un113_pixel_4_0_15__un1_beamylto9_0_LC_2_4_4 (
            .in0(N__14469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14824),
            .lcout(),
            .ltout(un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un1_beamylto9_3_0_LC_2_4_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un1_beamylto9_3_0_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un1_beamylto9_3_0_LC_2_4_5.LUT_INIT=16'b0001000000110000;
    LogicCell40 un113_pixel_4_0_15__un1_beamylto9_3_0_LC_2_4_5 (
            .in0(N__23284),
            .in1(N__14687),
            .in2(N__10469),
            .in3(N__20825),
            .lcout(un113_pixel_4_0_15__un1_beamylto9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIID25_8_LC_2_5_1.C_ON=1'b0;
    defparam beamY_RNIID25_8_LC_2_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIID25_8_LC_2_5_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamY_RNIID25_8_LC_2_5_1 (
            .in0(N__14783),
            .in1(N__12973),
            .in2(N__14890),
            .in3(N__12882),
            .lcout(),
            .ltout(un5_visibley_axbxc7_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_9_LC_2_5_2.C_ON=1'b0;
    defparam beamY_RNISI4A_9_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_9_LC_2_5_2.LUT_INIT=16'b1001101001011010;
    LogicCell40 beamY_RNISI4A_9_LC_2_5_2 (
            .in0(N__14973),
            .in1(N__14622),
            .in2(N__10466),
            .in3(N__11245),
            .lcout(chary_if_generate_plus_mult1_un33_sum_axb3),
            .ltout(chary_if_generate_plus_mult1_un33_sum_axb3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_1_tz_LC_2_5_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_1_tz_LC_2_5_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_1_tz_LC_2_5_3.LUT_INIT=16'b0000000100000100;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_1_tz_LC_2_5_3 (
            .in0(N__12477),
            .in1(N__12636),
            .in2(N__10463),
            .in3(N__18107),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_6_LC_2_5_4.C_ON=1'b0;
    defparam beamY_RNI2KA6_6_LC_2_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_6_LC_2_5_4.LUT_INIT=16'b0110000010100000;
    LogicCell40 beamY_RNI2KA6_6_LC_2_5_4 (
            .in0(N__12883),
            .in1(N__14623),
            .in2(N__12989),
            .in3(N__11246),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFS4T_0_7_LC_2_5_6.C_ON=1'b0;
    defparam beamY_RNIFS4T_0_7_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIFS4T_0_7_LC_2_5_6.LUT_INIT=16'b0000000010000010;
    LogicCell40 beamY_RNIFS4T_0_7_LC_2_5_6 (
            .in0(N__18108),
            .in1(N__14784),
            .in2(N__12768),
            .in3(N__18226),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_sx_LC_2_5_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_sx_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_sx_LC_2_5_7.LUT_INIT=16'b1010000011101100;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_sx_LC_2_5_7 (
            .in0(N__11404),
            .in1(N__10505),
            .in2(N__10499),
            .in3(N__13996),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9425_0_6_LC_2_6_1.C_ON=1'b0;
    defparam beamY_RNI9425_0_6_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI9425_0_6_LC_2_6_1.LUT_INIT=16'b1010100110011001;
    LogicCell40 beamY_RNI9425_0_6_LC_2_6_1 (
            .in0(N__12977),
            .in1(N__12884),
            .in2(N__14659),
            .in3(N__20753),
            .lcout(),
            .ltout(beamY_RNI9425_0Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPOR8_0_6_LC_2_6_2.C_ON=1'b0;
    defparam beamY_RNIPOR8_0_6_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIPOR8_0_6_LC_2_6_2.LUT_INIT=16'b1110001011010001;
    LogicCell40 beamY_RNIPOR8_0_6_LC_2_6_2 (
            .in0(N__12885),
            .in1(N__14418),
            .in2(N__10496),
            .in3(N__12978),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIL62O_0_7_LC_2_6_3.C_ON=1'b0;
    defparam beamY_RNIL62O_0_7_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIL62O_0_7_LC_2_6_3.LUT_INIT=16'b0000010000000001;
    LogicCell40 beamY_RNIL62O_0_7_LC_2_6_3 (
            .in0(N__12453),
            .in1(N__12749),
            .in2(N__10493),
            .in3(N__14789),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_d_0_LC_2_6_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_d_0_LC_2_6_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_d_0_LC_2_6_4.LUT_INIT=16'b0111001110110111;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_c4_d_0_LC_2_6_4 (
            .in0(N__18222),
            .in1(N__12626),
            .in2(N__18139),
            .in3(N__13965),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_c4_d),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_8_LC_2_6_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_8_LC_2_6_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_8_LC_2_6_5.LUT_INIT=16'b0010000000001000;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_8_LC_2_6_5 (
            .in0(N__12625),
            .in1(N__18102),
            .in2(N__13997),
            .in3(N__18223),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIL62O_7_LC_2_6_6.C_ON=1'b0;
    defparam beamY_RNIL62O_7_LC_2_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIL62O_7_LC_2_6_6.LUT_INIT=16'b0001001000000000;
    LogicCell40 beamY_RNIL62O_7_LC_2_6_6 (
            .in0(N__14790),
            .in1(N__12454),
            .in2(N__12761),
            .in3(N__12627),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_0_LC_2_6_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_0_LC_2_6_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_0_LC_2_6_7.LUT_INIT=16'b1110001000000000;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_0_LC_2_6_7 (
            .in0(N__11263),
            .in1(N__18106),
            .in2(N__10490),
            .in3(N__18224),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x0_LC_2_7_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x0_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x0_LC_2_7_1.LUT_INIT=16'b0000111000000111;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_x0_LC_2_7_1 (
            .in0(N__18135),
            .in1(N__14785),
            .in2(N__12663),
            .in3(N__18254),
            .lcout(if_generate_plus_mult1_un61_sum_ac0_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9425_6_LC_2_7_2.C_ON=1'b0;
    defparam beamY_RNI9425_6_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI9425_6_LC_2_7_2.LUT_INIT=16'b1111111011101110;
    LogicCell40 beamY_RNI9425_6_LC_2_7_2 (
            .in0(N__12979),
            .in1(N__12886),
            .in2(N__14660),
            .in3(N__20755),
            .lcout(),
            .ltout(beamY_RNI9425Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPOR8_6_LC_2_7_3.C_ON=1'b0;
    defparam beamY_RNIPOR8_6_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIPOR8_6_LC_2_7_3.LUT_INIT=16'b1111001111100010;
    LogicCell40 beamY_RNIPOR8_6_LC_2_7_3 (
            .in0(N__12890),
            .in1(N__14420),
            .in2(N__10541),
            .in3(N__12980),
            .lcout(un5_visibley_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x1_LC_2_7_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x1_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_x1_LC_2_7_4.LUT_INIT=16'b0000000011011011;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_x1_LC_2_7_4 (
            .in0(N__18253),
            .in1(N__18136),
            .in2(N__14810),
            .in3(N__12631),
            .lcout(if_generate_plus_mult1_un61_sum_ac0_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_5_LC_2_7_5.C_ON=1'b0;
    defparam beamY_RNI6125_5_LC_2_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_5_LC_2_7_5.LUT_INIT=16'b1000011100001111;
    LogicCell40 beamY_RNI6125_5_LC_2_7_5 (
            .in0(N__20754),
            .in1(N__14419),
            .in2(N__12899),
            .in3(N__14630),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_7_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_7_6.LUT_INIT=16'b0001011010000001;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_7_6 (
            .in0(N__18255),
            .in1(N__12632),
            .in2(N__14028),
            .in3(N__18138),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_7_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_7_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_7_7.LUT_INIT=16'b0010010010010010;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_7_7 (
            .in0(N__18137),
            .in1(N__18256),
            .in2(N__12664),
            .in3(N__14001),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_ns_LC_2_8_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_ns_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_ns_LC_2_8_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_ns_LC_2_8_0 (
            .in0(N__12745),
            .in1(N__10538),
            .in2(_gnd_net_),
            .in3(N__10532),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0_6),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI75QM4_5_LC_2_8_1.C_ON=1'b0;
    defparam beamY_RNI75QM4_5_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI75QM4_5_LC_2_8_1.LUT_INIT=16'b0000000011001000;
    LogicCell40 beamY_RNI75QM4_5_LC_2_8_1 (
            .in0(N__12407),
            .in1(N__10520),
            .in2(N__10511),
            .in3(N__11526),
            .lcout(beamY_RNI75QM4Z0Z_5),
            .ltout(beamY_RNI75QM4Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x1_LC_2_8_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x1_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_x1_LC_2_8_2.LUT_INIT=16'b0110011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_x1_LC_2_8_2 (
            .in0(N__11527),
            .in1(N__12286),
            .in2(N__10508),
            .in3(N__10606),
            .lcout(),
            .ltout(if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_ns_LC_2_8_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_ns_LC_2_8_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_ns_LC_2_8_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_ns_LC_2_8_3 (
            .in0(_gnd_net_),
            .in1(N__10616),
            .in2(N__10610),
            .in3(N__11556),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_LC_2_8_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_LC_2_8_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_LC_2_8_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_LC_2_8_4 (
            .in0(N__11358),
            .in1(N__11336),
            .in2(_gnd_net_),
            .in3(N__11377),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_c4_LC_2_8_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_c4_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_c4_LC_2_8_5.LUT_INIT=16'b0000110001001101;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_c4_LC_2_8_5 (
            .in0(N__10607),
            .in1(N__13230),
            .in2(N__12455),
            .in3(N__10572),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_cZ0Z4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_LC_2_8_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_LC_2_8_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_LC_2_8_6.LUT_INIT=16'b0011001111101110;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_LC_2_8_6 (
            .in0(N__13229),
            .in1(N__12408),
            .in2(_gnd_net_),
            .in3(N__14521),
            .lcout(),
            .ltout(if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_ns_LC_2_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_ns_LC_2_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_ns_LC_2_8_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_ns_LC_2_8_7 (
            .in0(_gnd_net_),
            .in1(N__10583),
            .in2(N__10577),
            .in3(N__10571),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_1_2_LC_2_9_0.C_ON=1'b0;
    defparam voltage_0_RNO_1_2_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_1_2_LC_2_9_0.LUT_INIT=16'b0010001110101111;
    LogicCell40 voltage_0_RNO_1_2_LC_2_9_0 (
            .in0(N__11697),
            .in1(N__11980),
            .in2(N__10702),
            .in3(N__11678),
            .lcout(),
            .ltout(voltage_0_10_iv_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_2_LC_2_9_1.C_ON=1'b0;
    defparam voltage_0_2_LC_2_9_1.SEQ_MODE=4'b1000;
    defparam voltage_0_2_LC_2_9_1.LUT_INIT=16'b0011111100001111;
    LogicCell40 voltage_0_2_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__17976),
            .in2(N__10553),
            .in3(N__10550),
            .lcout(voltage_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19955),
            .ce(),
            .sr(N__18542));
    defparam voltage_1_RNO_1_2_LC_2_9_2.C_ON=1'b0;
    defparam voltage_1_RNO_1_2_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_1_2_LC_2_9_2.LUT_INIT=16'b0000101110111011;
    LogicCell40 voltage_1_RNO_1_2_LC_2_9_2 (
            .in0(N__11698),
            .in1(N__11656),
            .in2(N__10703),
            .in3(N__11679),
            .lcout(),
            .ltout(voltage_1_9_iv_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_2_LC_2_9_3.C_ON=1'b0;
    defparam voltage_1_2_LC_2_9_3.SEQ_MODE=4'b1000;
    defparam voltage_1_2_LC_2_9_3.LUT_INIT=16'b1110111100001111;
    LogicCell40 voltage_1_2_LC_2_9_3 (
            .in0(N__11859),
            .in1(N__15766),
            .in2(N__10544),
            .in3(N__10889),
            .lcout(voltage_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19955),
            .ce(),
            .sr(N__18542));
    defparam counter_RNIVSBN2_0_LC_2_9_4.C_ON=1'b0;
    defparam counter_RNIVSBN2_0_LC_2_9_4.SEQ_MODE=4'b0000;
    defparam counter_RNIVSBN2_0_LC_2_9_4.LUT_INIT=16'b0000000010011001;
    LogicCell40 counter_RNIVSBN2_0_LC_2_9_4 (
            .in0(N__15764),
            .in1(N__16285),
            .in2(_gnd_net_),
            .in3(N__11858),
            .lcout(un1_voltage_012_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_1_2_LC_2_9_5.C_ON=1'b0;
    defparam voltage_3_RNO_1_2_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_1_2_LC_2_9_5.LUT_INIT=16'b0100010111001111;
    LogicCell40 voltage_3_RNO_1_2_LC_2_9_5 (
            .in0(N__11680),
            .in1(N__11699),
            .in2(N__11981),
            .in3(N__11933),
            .lcout(),
            .ltout(voltage_3_9_iv_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_2_LC_2_9_6.C_ON=1'b0;
    defparam voltage_3_2_LC_2_9_6.SEQ_MODE=4'b1000;
    defparam voltage_3_2_LC_2_9_6.LUT_INIT=16'b1100111101001111;
    LogicCell40 voltage_3_2_LC_2_9_6 (
            .in0(N__15765),
            .in1(N__10652),
            .in2(N__10643),
            .in3(N__11860),
            .lcout(voltage_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19955),
            .ce(),
            .sr(N__18542));
    defparam voltage_1_RNI359O_2_LC_2_9_7.C_ON=1'b0;
    defparam voltage_1_RNI359O_2_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam voltage_1_RNI359O_2_LC_2_9_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 voltage_1_RNI359O_2_LC_2_9_7 (
            .in0(N__16577),
            .in1(N__15245),
            .in2(_gnd_net_),
            .in3(N__15763),
            .lcout(N_1509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_1_0_LC_2_10_0.C_ON=1'b0;
    defparam voltage_2_RNO_1_0_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_1_0_LC_2_10_0.LUT_INIT=16'b0101000111110011;
    LogicCell40 voltage_2_RNO_1_0_LC_2_10_0 (
            .in0(N__11914),
            .in1(N__11645),
            .in2(N__12043),
            .in3(N__10746),
            .lcout(voltage_2_9_iv_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIO70L4_0_LC_2_10_1.C_ON=1'b0;
    defparam counter_RNIO70L4_0_LC_2_10_1.SEQ_MODE=4'b0000;
    defparam counter_RNIO70L4_0_LC_2_10_1.LUT_INIT=16'b1010110000000000;
    LogicCell40 counter_RNIO70L4_0_LC_2_10_1 (
            .in0(N__10756),
            .in1(N__15512),
            .in2(N__16286),
            .in3(N__10727),
            .lcout(),
            .ltout(CO2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI8TL66_0_LC_2_10_2.C_ON=1'b0;
    defparam counter_RNI8TL66_0_LC_2_10_2.SEQ_MODE=4'b0000;
    defparam counter_RNI8TL66_0_LC_2_10_2.LUT_INIT=16'b0101101000111100;
    LogicCell40 counter_RNI8TL66_0_LC_2_10_2 (
            .in0(N__10778),
            .in1(N__10820),
            .in2(N__10640),
            .in3(N__16282),
            .lcout(N_1155),
            .ltout(N_1155_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_0_3_LC_2_10_3.C_ON=1'b0;
    defparam voltage_0_RNO_0_3_LC_2_10_3.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_0_3_LC_2_10_3.LUT_INIT=16'b0000101110111011;
    LogicCell40 voltage_0_RNO_0_3_LC_2_10_3 (
            .in0(N__10799),
            .in1(N__10684),
            .in2(N__10637),
            .in3(N__11963),
            .lcout(voltage_0_10_iv_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_1_1_LC_2_10_4.C_ON=1'b0;
    defparam voltage_2_RNO_1_1_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_1_1_LC_2_10_4.LUT_INIT=16'b0000110111011101;
    LogicCell40 voltage_2_RNO_1_1_LC_2_10_4 (
            .in0(N__11915),
            .in1(N__11774),
            .in2(N__11657),
            .in3(N__12003),
            .lcout(voltage_2_9_iv_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_1_0_LC_2_10_5.C_ON=1'b0;
    defparam voltage_0_RNO_1_0_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_1_0_LC_2_10_5.LUT_INIT=16'b0101111100010011;
    LogicCell40 voltage_0_RNO_1_0_LC_2_10_5 (
            .in0(N__10747),
            .in1(N__11961),
            .in2(N__10694),
            .in3(N__10628),
            .lcout(voltage_0_10_iv_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIO70L4_0_0_LC_2_10_6.C_ON=1'b0;
    defparam counter_RNIO70L4_0_0_LC_2_10_6.SEQ_MODE=4'b0000;
    defparam counter_RNIO70L4_0_0_LC_2_10_6.LUT_INIT=16'b0110011001011010;
    LogicCell40 counter_RNIO70L4_0_0_LC_2_10_6 (
            .in0(N__10726),
            .in1(N__10757),
            .in2(N__15519),
            .in3(N__16278),
            .lcout(N_1154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNO_1_1_LC_2_10_7.C_ON=1'b0;
    defparam voltage_0_RNO_1_1_LC_2_10_7.SEQ_MODE=4'b0000;
    defparam voltage_0_RNO_1_1_LC_2_10_7.LUT_INIT=16'b0000101110111011;
    LogicCell40 voltage_0_RNO_1_1_LC_2_10_7 (
            .in0(N__11773),
            .in1(N__10683),
            .in2(N__12005),
            .in3(N__11962),
            .lcout(voltage_0_10_iv_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_1_3_LC_2_11_0.C_ON=1'b0;
    defparam voltage_1_RNO_1_3_LC_2_11_0.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_1_3_LC_2_11_0.LUT_INIT=16'b0101111100010011;
    LogicCell40 voltage_1_RNO_1_3_LC_2_11_0 (
            .in0(N__10714),
            .in1(N__11643),
            .in2(N__10695),
            .in3(N__10794),
            .lcout(voltage_1_9_iv_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_1_3_LC_2_11_1.C_ON=1'b0;
    defparam voltage_3_RNO_1_3_LC_2_11_1.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_1_3_LC_2_11_1.LUT_INIT=16'b0010001110101111;
    LogicCell40 voltage_3_RNO_1_3_LC_2_11_1 (
            .in0(N__10795),
            .in1(N__11913),
            .in2(N__11975),
            .in3(N__10715),
            .lcout(voltage_3_9_iv_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_1_0_LC_2_11_2.C_ON=1'b0;
    defparam voltage_1_RNO_1_0_LC_2_11_2.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_1_0_LC_2_11_2.LUT_INIT=16'b0101000111110011;
    LogicCell40 voltage_1_RNO_1_0_LC_2_11_2 (
            .in0(N__10748),
            .in1(N__10685),
            .in2(N__12042),
            .in3(N__11644),
            .lcout(voltage_1_9_iv_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNICMA33_0_LC_2_11_3.C_ON=1'b0;
    defparam counter_RNICMA33_0_LC_2_11_3.SEQ_MODE=4'b0000;
    defparam counter_RNICMA33_0_LC_2_11_3.LUT_INIT=16'b1000110010000000;
    LogicCell40 counter_RNICMA33_0_LC_2_11_3 (
            .in0(N__13118),
            .in1(N__12031),
            .in2(N__16283),
            .in3(N__11726),
            .lcout(CO1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI2ACM1_1_0_LC_2_11_4.C_ON=1'b0;
    defparam counter_RNI2ACM1_1_0_LC_2_11_4.SEQ_MODE=4'b0000;
    defparam counter_RNI2ACM1_1_0_LC_2_11_4.LUT_INIT=16'b0001000000000000;
    LogicCell40 counter_RNI2ACM1_1_0_LC_2_11_4 (
            .in0(N__19309),
            .in1(N__15742),
            .in2(N__13348),
            .in3(N__16256),
            .lcout(voltage_2_1_sqmuxa),
            .ltout(voltage_2_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_1_3_LC_2_11_5.C_ON=1'b0;
    defparam voltage_2_RNO_1_3_LC_2_11_5.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_1_3_LC_2_11_5.LUT_INIT=16'b0000101110111011;
    LogicCell40 voltage_2_RNO_1_3_LC_2_11_5 (
            .in0(N__10793),
            .in1(N__11912),
            .in2(N__10718),
            .in3(N__10713),
            .lcout(voltage_2_9_iv_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI2ACM1_2_0_LC_2_11_6.C_ON=1'b0;
    defparam counter_RNI2ACM1_2_0_LC_2_11_6.SEQ_MODE=4'b0000;
    defparam counter_RNI2ACM1_2_0_LC_2_11_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNI2ACM1_2_0_LC_2_11_6 (
            .in0(N__19308),
            .in1(N__15741),
            .in2(N__13347),
            .in3(N__16255),
            .lcout(voltage_1_1_sqmuxa),
            .ltout(voltage_1_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_1_1_LC_2_11_7.C_ON=1'b0;
    defparam voltage_1_RNO_1_1_LC_2_11_7.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_1_1_LC_2_11_7.LUT_INIT=16'b0011111100010101;
    LogicCell40 voltage_1_RNO_1_1_LC_2_11_7 (
            .in0(N__11642),
            .in1(N__12004),
            .in2(N__10841),
            .in3(N__11771),
            .lcout(voltage_1_9_iv_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_3_LC_2_12_0.C_ON=1'b0;
    defparam voltage_1_3_LC_2_12_0.SEQ_MODE=4'b1000;
    defparam voltage_1_3_LC_2_12_0.LUT_INIT=16'b1111110101010101;
    LogicCell40 voltage_1_3_LC_2_12_0 (
            .in0(N__10838),
            .in1(N__11863),
            .in2(N__15733),
            .in3(N__10874),
            .lcout(voltage_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19961),
            .ce(),
            .sr(N__18544));
    defparam voltage_1_RNI579O_3_LC_2_12_1.C_ON=1'b0;
    defparam voltage_1_RNI579O_3_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam voltage_1_RNI579O_3_LC_2_12_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 voltage_1_RNI579O_3_LC_2_12_1 (
            .in0(N__19449),
            .in1(N__15162),
            .in2(_gnd_net_),
            .in3(N__15641),
            .lcout(N_1510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_3_LC_2_12_2.C_ON=1'b0;
    defparam voltage_3_3_LC_2_12_2.SEQ_MODE=4'b1000;
    defparam voltage_3_3_LC_2_12_2.LUT_INIT=16'b1011101100111011;
    LogicCell40 voltage_3_3_LC_2_12_2 (
            .in0(N__10832),
            .in1(N__10826),
            .in2(N__15734),
            .in3(N__11864),
            .lcout(voltage_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19961),
            .ce(),
            .sr(N__18544));
    defparam voltage_0_RNI313M_3_LC_2_12_4.C_ON=1'b0;
    defparam voltage_0_RNI313M_3_LC_2_12_4.SEQ_MODE=4'b0000;
    defparam voltage_0_RNI313M_3_LC_2_12_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 voltage_0_RNI313M_3_LC_2_12_4 (
            .in0(N__15642),
            .in1(N__15209),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(),
            .ltout(N_1506_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIGLLH1_0_LC_2_12_5.C_ON=1'b0;
    defparam counter_RNIGLLH1_0_LC_2_12_5.SEQ_MODE=4'b0000;
    defparam counter_RNIGLLH1_0_LC_2_12_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 counter_RNIGLLH1_0_LC_2_12_5 (
            .in0(_gnd_net_),
            .in1(N__10816),
            .in2(N__10805),
            .in3(N__16243),
            .lcout(counter_RNIGLLH1Z0Z_0),
            .ltout(counter_RNIGLLH1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI4K0L4_0_LC_2_12_6.C_ON=1'b0;
    defparam counter_RNI4K0L4_0_LC_2_12_6.SEQ_MODE=4'b0000;
    defparam counter_RNI4K0L4_0_LC_2_12_6.LUT_INIT=16'b1111000010100101;
    LogicCell40 counter_RNI4K0L4_0_LC_2_12_6 (
            .in0(N__11591),
            .in1(_gnd_net_),
            .in2(N__10802),
            .in3(N__11772),
            .lcout(N_2063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_RNI313M_0_3_LC_2_12_7.C_ON=1'b0;
    defparam voltage_0_RNI313M_0_3_LC_2_12_7.SEQ_MODE=4'b0000;
    defparam voltage_0_RNI313M_0_3_LC_2_12_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 voltage_0_RNI313M_0_3_LC_2_12_7 (
            .in0(N__19419),
            .in1(_gnd_net_),
            .in2(N__15219),
            .in3(N__15643),
            .lcout(N_1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_1_1_cry_0_0_c_LC_2_13_0.C_ON=1'b1;
    defparam un1_voltage_1_1_cry_0_0_c_LC_2_13_0.SEQ_MODE=4'b0000;
    defparam un1_voltage_1_1_cry_0_0_c_LC_2_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_voltage_1_1_cry_0_0_c_LC_2_13_0 (
            .in0(_gnd_net_),
            .in1(N__15339),
            .in2(N__10769),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(un1_voltage_1_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_0_1_LC_2_13_1.C_ON=1'b1;
    defparam voltage_1_RNO_0_1_LC_2_13_1.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_0_1_LC_2_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_1_RNO_0_1_LC_2_13_1 (
            .in0(_gnd_net_),
            .in1(N__15104),
            .in2(N__10907),
            .in3(N__10898),
            .lcout(voltage_1_RNO_0Z0Z_1),
            .ltout(),
            .carryin(un1_voltage_1_1_cry_0),
            .carryout(un1_voltage_1_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_0_2_LC_2_13_2.C_ON=1'b1;
    defparam voltage_1_RNO_0_2_LC_2_13_2.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_0_2_LC_2_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_1_RNO_0_2_LC_2_13_2 (
            .in0(_gnd_net_),
            .in1(N__10895),
            .in2(N__15262),
            .in3(N__10880),
            .lcout(voltage_1_RNO_0Z0Z_2),
            .ltout(),
            .carryin(un1_voltage_1_1_cry_1),
            .carryout(un1_voltage_1_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNO_0_3_LC_2_13_3.C_ON=1'b0;
    defparam voltage_1_RNO_0_3_LC_2_13_3.SEQ_MODE=4'b0000;
    defparam voltage_1_RNO_0_3_LC_2_13_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 voltage_1_RNO_0_3_LC_2_13_3 (
            .in0(N__15163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10877),
            .lcout(voltage_1_RNO_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIJTI6_2_LC_2_13_4.C_ON=1'b0;
    defparam counter_RNIJTI6_2_LC_2_13_4.SEQ_MODE=4'b0000;
    defparam counter_RNIJTI6_2_LC_2_13_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 counter_RNIJTI6_2_LC_2_13_4 (
            .in0(N__15936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15721),
            .lcout(Z_decfrac4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI1SFG_5_LC_2_13_5.C_ON=1'b0;
    defparam counter_RNI1SFG_5_LC_2_13_5.SEQ_MODE=4'b0000;
    defparam counter_RNI1SFG_5_LC_2_13_5.LUT_INIT=16'b0000000100000000;
    LogicCell40 counter_RNI1SFG_5_LC_2_13_5 (
            .in0(N__13863),
            .in1(N__13771),
            .in2(N__16399),
            .in3(N__13643),
            .lcout(),
            .ltout(un6_slaveselectlto9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIS6CQ_2_LC_2_13_6.C_ON=1'b0;
    defparam counter_RNIS6CQ_2_LC_2_13_6.SEQ_MODE=4'b0000;
    defparam counter_RNIS6CQ_2_LC_2_13_6.LUT_INIT=16'b0101000001110000;
    LogicCell40 counter_RNIS6CQ_2_LC_2_13_6 (
            .in0(N__15937),
            .in1(N__16267),
            .in2(N__10868),
            .in3(N__15722),
            .lcout(),
            .ltout(un6_slaveselect_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIHC2O1_2_LC_2_13_7.C_ON=1'b0;
    defparam counter_RNIHC2O1_2_LC_2_13_7.SEQ_MODE=4'b0000;
    defparam counter_RNIHC2O1_2_LC_2_13_7.LUT_INIT=16'b0000000000001010;
    LogicCell40 counter_RNIHC2O1_2_LC_2_13_7 (
            .in0(N__13625),
            .in1(_gnd_net_),
            .in2(N__10865),
            .in3(N__10862),
            .lcout(un5_slaveselect),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_2_1_cry_0_c_LC_2_14_0.C_ON=1'b1;
    defparam un1_voltage_2_1_cry_0_c_LC_2_14_0.SEQ_MODE=4'b0000;
    defparam un1_voltage_2_1_cry_0_c_LC_2_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_voltage_2_1_cry_0_c_LC_2_14_0 (
            .in0(_gnd_net_),
            .in1(N__15395),
            .in2(N__13100),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(un1_voltage_2_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_0_1_LC_2_14_1.C_ON=1'b1;
    defparam voltage_2_RNO_0_1_LC_2_14_1.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_0_1_LC_2_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_2_RNO_0_1_LC_2_14_1 (
            .in0(_gnd_net_),
            .in1(N__15142),
            .in2(N__10856),
            .in3(N__10844),
            .lcout(voltage_2_RNO_0Z0Z_1),
            .ltout(),
            .carryin(un1_voltage_2_1_cry_0),
            .carryout(un1_voltage_2_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_0_2_LC_2_14_2.C_ON=1'b1;
    defparam voltage_2_RNO_0_2_LC_2_14_2.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_0_2_LC_2_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 voltage_2_RNO_0_2_LC_2_14_2 (
            .in0(_gnd_net_),
            .in1(N__10979),
            .in2(N__15305),
            .in3(N__10973),
            .lcout(voltage_2_RNO_0Z0Z_2),
            .ltout(),
            .carryin(un1_voltage_2_1_cry_1),
            .carryout(un1_voltage_2_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_3_LC_2_14_3.C_ON=1'b0;
    defparam voltage_2_3_LC_2_14_3.SEQ_MODE=4'b1000;
    defparam voltage_2_3_LC_2_14_3.LUT_INIT=16'b0001111100101111;
    LogicCell40 voltage_2_3_LC_2_14_3 (
            .in0(N__10970),
            .in1(N__13421),
            .in2(N__10964),
            .in3(N__10952),
            .lcout(voltage_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19966),
            .ce(),
            .sr(N__18547));
    defparam counter_RNIJTI6_3_LC_2_15_0.C_ON=1'b0;
    defparam counter_RNIJTI6_3_LC_2_15_0.SEQ_MODE=4'b0000;
    defparam counter_RNIJTI6_3_LC_2_15_0.LUT_INIT=16'b0000000010101010;
    LogicCell40 counter_RNIJTI6_3_LC_2_15_0 (
            .in0(N__16257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16408),
            .lcout(N_46_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_3_RNO_0_0_LC_2_15_1.C_ON=1'b0;
    defparam ScreenBuffer_0_3_RNO_0_0_LC_2_15_1.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_3_RNO_0_0_LC_2_15_1.LUT_INIT=16'b0000000000000010;
    LogicCell40 ScreenBuffer_0_3_RNO_0_0_LC_2_15_1 (
            .in0(N__16410),
            .in1(N__15992),
            .in2(N__15816),
            .in3(N__16259),
            .lcout(),
            .ltout(un1_sclk17_2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_3_0_LC_2_15_2.C_ON=1'b0;
    defparam ScreenBuffer_0_3_0_LC_2_15_2.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_3_0_LC_2_15_2.LUT_INIT=16'b1011111110000000;
    LogicCell40 ScreenBuffer_0_3_0_LC_2_15_2 (
            .in0(N__20194),
            .in1(N__20062),
            .in2(N__10928),
            .in3(N__23647),
            .lcout(ScreenBuffer_0_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19969),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_10_RNO_0_0_LC_2_15_3.C_ON=1'b0;
    defparam ScreenBuffer_0_10_RNO_0_0_LC_2_15_3.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_10_RNO_0_0_LC_2_15_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 ScreenBuffer_0_10_RNO_0_0_LC_2_15_3 (
            .in0(N__16409),
            .in1(N__15991),
            .in2(N__15815),
            .in3(N__16258),
            .lcout(),
            .ltout(un1_sclk17_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_10_0_LC_2_15_4.C_ON=1'b0;
    defparam ScreenBuffer_0_10_0_LC_2_15_4.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_10_0_LC_2_15_4.LUT_INIT=16'b1011111110000000;
    LogicCell40 ScreenBuffer_0_10_0_LC_2_15_4 (
            .in0(N__20193),
            .in1(N__20061),
            .in2(N__10925),
            .in3(N__23707),
            .lcout(ScreenBuffer_0_10Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19969),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_1_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_1_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_1_0 (
            .in0(_gnd_net_),
            .in1(N__13276),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_1_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3Q404_LC_4_1_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3Q404_LC_4_1_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3Q404_LC_4_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3Q404_LC_4_1_1 (
            .in0(_gnd_net_),
            .in1(N__11034),
            .in2(N__10922),
            .in3(N__10910),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40I45_LC_4_1_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40I45_LC_4_1_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40I45_LC_4_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40I45_LC_4_1_2 (
            .in0(_gnd_net_),
            .in1(N__11036),
            .in2(N__11093),
            .in3(N__11081),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3S246_LC_4_1_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3S246_LC_4_1_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3S246_LC_4_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3S246_LC_4_1_3 (
            .in0(_gnd_net_),
            .in1(N__11035),
            .in2(N__11078),
            .in3(N__11066),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIRSJ6F_LC_4_1_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIRSJ6F_LC_4_1_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIRSJ6F_LC_4_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIRSJ6F_LC_4_1_4 (
            .in0(N__11188),
            .in1(N__11009),
            .in2(N__11063),
            .in3(N__11051),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_LC_4_1_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_LC_4_1_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_LC_4_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_LC_4_1_5 (
            .in0(_gnd_net_),
            .in1(N__11048),
            .in2(_gnd_net_),
            .in3(N__11039),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_0_LC_4_1_7.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_0_LC_4_1_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_0_LC_4_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_0_LC_4_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11033),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_4_2_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_4_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_4_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_4_2_0 (
            .in0(_gnd_net_),
            .in1(N__12555),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_2_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIV79_LC_4_2_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIV79_LC_4_2_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIV79_LC_4_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIV79_LC_4_2_1 (
            .in0(_gnd_net_),
            .in1(N__11183),
            .in2(N__11282),
            .in3(N__11003),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80D_LC_4_2_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80D_LC_4_2_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80D_LC_4_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80D_LC_4_2_2 (
            .in0(_gnd_net_),
            .in1(N__11000),
            .in2(N__11189),
            .in3(N__10994),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4E_LC_4_2_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4E_LC_4_2_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4E_LC_4_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4E_LC_4_2_3 (
            .in0(_gnd_net_),
            .in1(N__11187),
            .in2(N__10991),
            .in3(N__10982),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIK4SNU_LC_4_2_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIK4SNU_LC_4_2_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIK4SNU_LC_4_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIK4SNU_LC_4_2_4 (
            .in0(N__11121),
            .in1(N__11165),
            .in2(N__11210),
            .in3(N__11201),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJF_LC_4_2_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJF_LC_4_2_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJF_LC_4_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJF_LC_4_2_5 (
            .in0(_gnd_net_),
            .in1(N__11198),
            .in2(_gnd_net_),
            .in3(N__11192),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_0_LC_4_2_7.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_0_LC_4_2_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_0_LC_4_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_0_LC_4_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11182),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_3_0.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(N__12172),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_LC_4_3_1.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_LC_4_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_LC_4_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_LC_4_3_1 (
            .in0(_gnd_net_),
            .in1(N__11122),
            .in2(N__11291),
            .in3(N__11159),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUO_LC_4_3_2.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUO_LC_4_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUO_LC_4_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUO_LC_4_3_2 (
            .in0(_gnd_net_),
            .in1(N__11120),
            .in2(N__11156),
            .in3(N__11147),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NS_LC_4_3_3.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NS_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NS_LC_4_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NS_LC_4_3_3 (
            .in0(_gnd_net_),
            .in1(N__11123),
            .in2(N__11144),
            .in3(N__11135),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_4_3_4.C_ON=1'b1;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_4_3_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_4_3_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_4_3_4 (
            .in0(_gnd_net_),
            .in1(N__11099),
            .in2(N__11132),
            .in3(N__11119),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RU_LC_4_3_5.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RU_LC_4_3_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RU_LC_4_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RU_LC_4_3_5 (
            .in0(_gnd_net_),
            .in1(N__11300),
            .in2(_gnd_net_),
            .in3(N__11294),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_4_3_6.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_4_3_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_4_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_4_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12556),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_0.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13262),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEDF31_6_LC_4_4_3.C_ON=1'b0;
    defparam beamY_RNIEDF31_6_LC_4_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIEDF31_6_LC_4_4_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamY_RNIEDF31_6_LC_4_4_3 (
            .in0(N__14037),
            .in1(N__12690),
            .in2(N__12485),
            .in3(N__18291),
            .lcout(beamY_RNIEDF31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_4_4_7.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_4_4_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_4_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_4_4_7 (
            .in0(N__12176),
            .in1(N__21871),
            .in2(_gnd_net_),
            .in3(N__20832),
            .lcout(beamY_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6EUJ1_7_LC_4_5_0.C_ON=1'b0;
    defparam beamY_RNI6EUJ1_7_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI6EUJ1_7_LC_4_5_0.LUT_INIT=16'b0111011101010111;
    LogicCell40 beamY_RNI6EUJ1_7_LC_4_5_0 (
            .in0(N__18261),
            .in1(N__11270),
            .in2(N__11414),
            .in3(N__14020),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c4_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m1_5_LC_4_5_1.C_ON=1'b0;
    defparam row_1_if_m1_5_LC_4_5_1.SEQ_MODE=4'b0000;
    defparam row_1_if_m1_5_LC_4_5_1.LUT_INIT=16'b1001011001100101;
    LogicCell40 row_1_if_m1_5_LC_4_5_1 (
            .in0(N__12687),
            .in1(N__18140),
            .in2(N__14036),
            .in3(N__18260),
            .lcout(if_m1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_0_6_LC_4_5_2.C_ON=1'b0;
    defparam beamY_RNI2KA6_0_6_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_0_6_LC_4_5_2.LUT_INIT=16'b0001010001000100;
    LogicCell40 beamY_RNI2KA6_0_6_LC_4_5_2 (
            .in0(N__13001),
            .in1(N__12911),
            .in2(N__14701),
            .in3(N__11252),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4QBV1_6_LC_4_5_3.C_ON=1'b0;
    defparam beamY_RNI4QBV1_6_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI4QBV1_6_LC_4_5_3.LUT_INIT=16'b1101110011001100;
    LogicCell40 beamY_RNI4QBV1_6_LC_4_5_3 (
            .in0(N__14021),
            .in1(N__12323),
            .in2(N__11222),
            .in3(N__18141),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILILV4_8_LC_4_5_4.C_ON=1'b0;
    defparam beamY_RNILILV4_8_LC_4_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNILILV4_8_LC_4_5_4.LUT_INIT=16'b1111110011111101;
    LogicCell40 beamY_RNILILV4_8_LC_4_5_4 (
            .in0(N__18142),
            .in1(N__11219),
            .in2(N__11213),
            .in3(N__11423),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEG4HI_3_LC_4_5_5.C_ON=1'b0;
    defparam beamY_RNIEG4HI_3_LC_4_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIEG4HI_3_LC_4_5_5.LUT_INIT=16'b1111111011111010;
    LogicCell40 beamY_RNIEG4HI_3_LC_4_5_5 (
            .in0(N__11393),
            .in1(N__13310),
            .in2(N__11417),
            .in3(N__13231),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIER061_6_LC_4_5_7.C_ON=1'b0;
    defparam beamY_RNIER061_6_LC_4_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIER061_6_LC_4_5_7.LUT_INIT=16'b1000001000000000;
    LogicCell40 beamY_RNIER061_6_LC_4_5_7 (
            .in0(N__12719),
            .in1(N__18262),
            .in2(N__18169),
            .in3(N__11413),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIED3U1_0_7_LC_4_6_0.C_ON=1'b0;
    defparam beamY_RNIED3U1_0_7_LC_4_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIED3U1_0_7_LC_4_6_0.LUT_INIT=16'b0100101100101101;
    LogicCell40 beamY_RNIED3U1_0_7_LC_4_6_0 (
            .in0(N__12677),
            .in1(N__12721),
            .in2(N__11315),
            .in3(N__14035),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_4_6_1.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_4_6_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_0_3_LC_4_6_1 (
            .in0(_gnd_net_),
            .in1(N__14441),
            .in2(_gnd_net_),
            .in3(N__20790),
            .lcout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x0_LC_4_6_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x0_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x0_LC_4_6_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_ac0_5_x0_LC_4_6_2 (
            .in0(N__11334),
            .in1(N__11359),
            .in2(N__11387),
            .in3(N__11383),
            .lcout(if_generate_plus_mult1_un75_sum_ac0_5_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x1_LC_4_6_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x1_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_x1_LC_4_6_3.LUT_INIT=16'b1100110011001000;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_ac0_5_x1_LC_4_6_3 (
            .in0(N__11384),
            .in1(N__12544),
            .in2(N__11363),
            .in3(N__11335),
            .lcout(if_generate_plus_mult1_un75_sum_ac0_5_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFS4T_7_LC_4_6_4.C_ON=1'b0;
    defparam beamY_RNIFS4T_7_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIFS4T_7_LC_4_6_4.LUT_INIT=16'b1100001101101001;
    LogicCell40 beamY_RNIFS4T_7_LC_4_6_4 (
            .in0(N__18163),
            .in1(N__14812),
            .in2(N__12776),
            .in3(N__18285),
            .lcout(beamY_RNIFS4TZ0Z_7),
            .ltout(beamY_RNIFS4TZ0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIED3U1_7_LC_4_6_5.C_ON=1'b0;
    defparam beamY_RNIED3U1_7_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIED3U1_7_LC_4_6_5.LUT_INIT=16'b0101101111011010;
    LogicCell40 beamY_RNIED3U1_7_LC_4_6_5 (
            .in0(N__12720),
            .in1(N__14033),
            .in2(N__11306),
            .in3(N__12676),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQTGS2_8_LC_4_6_6.C_ON=1'b0;
    defparam beamY_RNIQTGS2_8_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIQTGS2_8_LC_4_6_6.LUT_INIT=16'b1010010101111000;
    LogicCell40 beamY_RNIQTGS2_8_LC_4_6_6 (
            .in0(N__18164),
            .in1(N__14034),
            .in2(N__11303),
            .in3(N__18286),
            .lcout(beamY_RNIQTGS2Z0Z_8),
            .ltout(beamY_RNIQTGS2Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPNEA3_6_LC_4_6_7.C_ON=1'b0;
    defparam beamY_RNIPNEA3_6_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIPNEA3_6_LC_4_6_7.LUT_INIT=16'b1100000011111100;
    LogicCell40 beamY_RNIPNEA3_6_LC_4_6_7 (
            .in0(_gnd_net_),
            .in1(N__12481),
            .in2(N__11474),
            .in3(N__12678),
            .lcout(chary_if_generate_plus_mult1_un54_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIO8DB4_6_LC_4_7_0.C_ON=1'b0;
    defparam beamY_RNIO8DB4_6_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIO8DB4_6_LC_4_7_0.LUT_INIT=16'b0100101100101101;
    LogicCell40 beamY_RNIO8DB4_6_LC_4_7_0 (
            .in0(N__12471),
            .in1(N__11455),
            .in2(N__12575),
            .in3(N__12692),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIECMV4_5_LC_4_7_1.C_ON=1'b0;
    defparam beamY_RNIECMV4_5_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIECMV4_5_LC_4_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNIECMV4_5_LC_4_7_1 (
            .in0(N__11449),
            .in1(N__11464),
            .in2(_gnd_net_),
            .in3(N__12469),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0JK7C_5_LC_4_7_2.C_ON=1'b0;
    defparam beamY_RNI0JK7C_5_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI0JK7C_5_LC_4_7_2.LUT_INIT=16'b0100101111010010;
    LogicCell40 beamY_RNI0JK7C_5_LC_4_7_2 (
            .in0(N__12567),
            .in1(N__11450),
            .in2(N__11471),
            .in3(N__11434),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb3),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axb3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIS0VDC_3_LC_4_7_3.C_ON=1'b0;
    defparam beamY_RNIS0VDC_3_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIS0VDC_3_LC_4_7_3.LUT_INIT=16'b0101000010100000;
    LogicCell40 beamY_RNIS0VDC_3_LC_4_7_3 (
            .in0(N__13270),
            .in1(_gnd_net_),
            .in2(N__11468),
            .in3(N__12545),
            .lcout(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_1_0_LC_4_7_4.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_1_0_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_1_0_LC_4_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un113_pixel_3_0_11__g0_1_0_LC_4_7_4 (
            .in0(_gnd_net_),
            .in1(N__14476),
            .in2(_gnd_net_),
            .in3(N__20831),
            .lcout(un5_visibley_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPNEA3_0_6_LC_4_7_5.C_ON=1'b0;
    defparam beamY_RNIPNEA3_0_6_LC_4_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIPNEA3_0_6_LC_4_7_5.LUT_INIT=16'b0101101010100101;
    LogicCell40 beamY_RNIPNEA3_0_6_LC_4_7_5 (
            .in0(N__12691),
            .in1(_gnd_net_),
            .in2(N__11456),
            .in3(N__12470),
            .lcout(beamY_RNIPNEA3_0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0K169_6_LC_4_7_6.C_ON=1'b0;
    defparam beamY_RNI0K169_6_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI0K169_6_LC_4_7_6.LUT_INIT=16'b0110101010101001;
    LogicCell40 beamY_RNI0K169_6_LC_4_7_6 (
            .in0(N__11465),
            .in1(N__11454),
            .in2(N__12574),
            .in3(N__11435),
            .lcout(beamY_RNI0K169Z0Z_6),
            .ltout(beamY_RNI0K169Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV42D31_0_6_LC_4_7_7.C_ON=1'b0;
    defparam beamY_RNIV42D31_0_6_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIV42D31_0_6_LC_4_7_7.LUT_INIT=16'b0110101010101001;
    LogicCell40 beamY_RNIV42D31_0_6_LC_4_7_7 (
            .in0(N__12520),
            .in1(N__13070),
            .in2(N__11426),
            .in3(N__13046),
            .lcout(beamY_RNIV42D31_0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g1_0_0_LC_4_8_0.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g1_0_0_LC_4_8_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g1_0_0_LC_4_8_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un113_pixel_3_0_11__g1_0_0_LC_4_8_0 (
            .in0(_gnd_net_),
            .in1(N__20841),
            .in2(_gnd_net_),
            .in3(N__14479),
            .lcout(un113_pixel_3_0_11__g1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_5_LC_4_8_1.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_5_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_5_LC_4_8_1.LUT_INIT=16'b0101101100011010;
    LogicCell40 un113_pixel_3_0_11__g0_5_LC_4_8_1 (
            .in0(N__13309),
            .in1(N__12818),
            .in2(N__13277),
            .in3(N__11573),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_3_LC_4_8_2.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_3_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_3_LC_4_8_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 un113_pixel_3_0_11__g0_3_LC_4_8_2 (
            .in0(N__12819),
            .in1(N__13159),
            .in2(N__11567),
            .in3(N__14481),
            .lcout(un113_pixel_3_0_11__N_4_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m1_x1_LC_4_8_3.C_ON=1'b0;
    defparam row_1_if_m1_x1_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam row_1_if_m1_x1_LC_4_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_m1_x1_LC_4_8_3 (
            .in0(N__12298),
            .in1(N__11540),
            .in2(N__14298),
            .in3(N__14689),
            .lcout(),
            .ltout(if_m1_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m1_ns_LC_4_8_4.C_ON=1'b0;
    defparam row_1_if_m1_ns_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam row_1_if_m1_ns_LC_4_8_4.LUT_INIT=16'b1111000010101010;
    LogicCell40 row_1_if_m1_ns_LC_4_8_4 (
            .in0(N__11504),
            .in1(_gnd_net_),
            .in2(N__11564),
            .in3(N__11561),
            .lcout(if_m1_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m1_x0_LC_4_8_5.C_ON=1'b0;
    defparam row_1_if_m1_x0_LC_4_8_5.SEQ_MODE=4'b0000;
    defparam row_1_if_m1_x0_LC_4_8_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 row_1_if_m1_x0_LC_4_8_5 (
            .in0(N__12297),
            .in1(N__11539),
            .in2(N__14297),
            .in3(N__14688),
            .lcout(if_m1_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_7_LC_4_8_6.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_7_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_7_LC_4_8_6.LUT_INIT=16'b1111111110011001;
    LogicCell40 un113_pixel_3_0_11__g0_7_LC_4_8_6 (
            .in0(N__13158),
            .in1(N__13308),
            .in2(_gnd_net_),
            .in3(N__14480),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_2_0_LC_4_8_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_2_0_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_2_0_LC_4_8_7.LUT_INIT=16'b1011100011100010;
    LogicCell40 un113_pixel_3_0_11__g0_2_0_LC_4_8_7 (
            .in0(N__11498),
            .in1(N__12820),
            .in2(N__11492),
            .in3(N__14690),
            .lcout(g1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_4_9_1.C_ON=1'b0;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_4_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19993),
            .lcout(GB_BUFFER_Clock12MHz_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIKUA33_0_LC_4_9_2.C_ON=1'b0;
    defparam counter_RNIKUA33_0_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam counter_RNIKUA33_0_LC_4_9_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNIKUA33_0_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(N__11587),
            .in2(_gnd_net_),
            .in3(N__11765),
            .lcout(N_1159_i),
            .ltout(N_1159_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_1_2_LC_4_9_3.C_ON=1'b0;
    defparam voltage_2_RNO_1_2_LC_4_9_3.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_1_2_LC_4_9_3.LUT_INIT=16'b0101000111110011;
    LogicCell40 voltage_2_RNO_1_2_LC_4_9_3 (
            .in0(N__11684),
            .in1(N__11932),
            .in2(N__11660),
            .in3(N__11655),
            .lcout(voltage_2_9_iv_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNIO5RB1_LC_4_9_5.C_ON=1'b0;
    defparam slaveselect_RNIO5RB1_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam slaveselect_RNIO5RB1_LC_4_9_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 slaveselect_RNIO5RB1_LC_4_9_5 (
            .in0(_gnd_net_),
            .in1(N__19292),
            .in2(_gnd_net_),
            .in3(N__13562),
            .lcout(voltage_0_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_4_LC_4_9_7.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_4_LC_4_9_7.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_4_LC_4_9_7.LUT_INIT=16'b0011001100110011;
    LogicCell40 slaveselect_RNILOQC2_4_LC_4_9_7 (
            .in0(_gnd_net_),
            .in1(N__11600),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_1_LC_4_10_0.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_1_LC_4_10_0.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_1_LC_4_10_0.LUT_INIT=16'b1000100010111011;
    LogicCell40 slaveselect_RNILOQC2_1_LC_4_10_0 (
            .in0(N__13556),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__17185),
            .lcout(slaveselect_RNILOQC2Z0Z_1),
            .ltout(slaveselect_RNILOQC2Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_4_LC_4_10_1.C_ON=1'b0;
    defparam ScreenBuffer_1_1_4_LC_4_10_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_1_4_LC_4_10_1.LUT_INIT=16'b1111001100000011;
    LogicCell40 ScreenBuffer_1_1_4_LC_4_10_1 (
            .in0(_gnd_net_),
            .in1(N__19288),
            .in2(N__11594),
            .in3(N__17149),
            .lcout(ScreenBuffer_1_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19962),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNICHLH1_0_LC_4_10_2.C_ON=1'b0;
    defparam counter_RNICHLH1_0_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam counter_RNICHLH1_0_LC_4_10_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 counter_RNICHLH1_0_LC_4_10_2 (
            .in0(N__16213),
            .in1(N__15521),
            .in2(_gnd_net_),
            .in3(N__15533),
            .lcout(counter_RNICHLH1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNIQDU22_LC_4_10_4.C_ON=1'b0;
    defparam slaveselect_RNIQDU22_LC_4_10_4.SEQ_MODE=4'b0000;
    defparam slaveselect_RNIQDU22_LC_4_10_4.LUT_INIT=16'b0101110001011100;
    LogicCell40 slaveselect_RNIQDU22_LC_4_10_4 (
            .in0(N__13557),
            .in1(N__18568),
            .in2(N__19328),
            .in3(_gnd_net_),
            .lcout(un1_counter_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNIE1PG2_LC_4_10_5.C_ON=1'b0;
    defparam slaveselect_RNIE1PG2_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam slaveselect_RNIE1PG2_LC_4_10_5.LUT_INIT=16'b1100110001010101;
    LogicCell40 slaveselect_RNIE1PG2_LC_4_10_5 (
            .in0(N__13336),
            .in1(N__13555),
            .in2(_gnd_net_),
            .in3(N__19284),
            .lcout(un1_voltage_012_0),
            .ltout(un1_voltage_012_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIVSBN2_0_0_LC_4_10_6.C_ON=1'b0;
    defparam counter_RNIVSBN2_0_0_LC_4_10_6.SEQ_MODE=4'b0000;
    defparam counter_RNIVSBN2_0_0_LC_4_10_6.LUT_INIT=16'b0000010100001010;
    LogicCell40 counter_RNIVSBN2_0_0_LC_4_10_6 (
            .in0(N__16214),
            .in1(_gnd_net_),
            .in2(N__12047),
            .in3(N__15862),
            .lcout(un1_voltage_012_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNICMA33_0_0_LC_4_11_0.C_ON=1'b0;
    defparam counter_RNICMA33_0_0_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam counter_RNICMA33_0_0_LC_4_11_0.LUT_INIT=16'b0010011111011000;
    LogicCell40 counter_RNICMA33_0_0_LC_4_11_0 (
            .in0(N__16248),
            .in1(N__13117),
            .in2(N__11725),
            .in3(N__12044),
            .lcout(N_1153),
            .ltout(N_1153_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_RNO_1_1_LC_4_11_1.C_ON=1'b0;
    defparam voltage_3_RNO_1_1_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam voltage_3_RNO_1_1_LC_4_11_1.LUT_INIT=16'b0000110111011101;
    LogicCell40 voltage_3_RNO_1_1_LC_4_11_1 (
            .in0(N__11976),
            .in1(N__11761),
            .in2(N__11936),
            .in3(N__11931),
            .lcout(),
            .ltout(voltage_3_9_iv_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_3_1_LC_4_11_2.C_ON=1'b0;
    defparam voltage_3_1_LC_4_11_2.SEQ_MODE=4'b1000;
    defparam voltage_3_1_LC_4_11_2.LUT_INIT=16'b1100111101001111;
    LogicCell40 voltage_3_1_LC_4_11_2 (
            .in0(N__15821),
            .in1(N__11882),
            .in2(N__11867),
            .in3(N__11840),
            .lcout(voltage_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19964),
            .ce(),
            .sr(N__18545));
    defparam voltage_1_1_LC_4_11_3.C_ON=1'b0;
    defparam voltage_1_1_LC_4_11_3.SEQ_MODE=4'b1000;
    defparam voltage_1_1_LC_4_11_3.LUT_INIT=16'b1111001110110011;
    LogicCell40 voltage_1_1_LC_4_11_3 (
            .in0(N__11839),
            .in1(N__11807),
            .in2(N__11798),
            .in3(N__15822),
            .lcout(voltage_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19964),
            .ce(),
            .sr(N__18545));
    defparam voltage_0_RNIVS2M_1_LC_4_11_4.C_ON=1'b0;
    defparam voltage_0_RNIVS2M_1_LC_4_11_4.SEQ_MODE=4'b0000;
    defparam voltage_0_RNIVS2M_1_LC_4_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 voltage_0_RNIVS2M_1_LC_4_11_4 (
            .in0(N__15820),
            .in1(N__15127),
            .in2(_gnd_net_),
            .in3(N__19051),
            .lcout(N_1504),
            .ltout(N_1504_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_1_c_RNO_LC_4_11_5.C_ON=1'b0;
    defparam un42_cry_1_c_RNO_LC_4_11_5.SEQ_MODE=4'b0000;
    defparam un42_cry_1_c_RNO_LC_4_11_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 un42_cry_1_c_RNO_LC_4_11_5 (
            .in0(_gnd_net_),
            .in1(N__16246),
            .in2(N__11783),
            .in3(N__11714),
            .lcout(un42_cry_1_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI8DLH1_0_LC_4_11_6.C_ON=1'b0;
    defparam counter_RNI8DLH1_0_LC_4_11_6.SEQ_MODE=4'b0000;
    defparam counter_RNI8DLH1_0_LC_4_11_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 counter_RNI8DLH1_0_LC_4_11_6 (
            .in0(N__16247),
            .in1(_gnd_net_),
            .in2(N__11724),
            .in3(N__11780),
            .lcout(counter_RNI8DLH1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_1_RNI139O_1_LC_4_11_7.C_ON=1'b0;
    defparam voltage_1_RNI139O_1_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam voltage_1_RNI139O_1_LC_4_11_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 voltage_1_RNI139O_1_LC_4_11_7 (
            .in0(N__19352),
            .in1(N__15086),
            .in2(_gnd_net_),
            .in3(N__15819),
            .lcout(N_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_3_LC_4_12_0.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_3_LC_4_12_0.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_3_LC_4_12_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 slaveselect_RNILOQC2_3_LC_4_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12064),
            .lcout(un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_4_LC_4_12_2.C_ON=1'b0;
    defparam ScreenBuffer_1_0_4_LC_4_12_2.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_0_4_LC_4_12_2.LUT_INIT=16'b1101110100010001;
    LogicCell40 ScreenBuffer_1_0_4_LC_4_12_2 (
            .in0(N__19291),
            .in1(N__12065),
            .in2(_gnd_net_),
            .in3(N__16954),
            .lcout(ScreenBuffer_1_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19967),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_3_LC_4_12_3.C_ON=1'b0;
    defparam counter_RNI6R5D_3_LC_4_12_3.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_3_LC_4_12_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 counter_RNI6R5D_3_LC_4_12_3 (
            .in0(N__16181),
            .in1(N__16347),
            .in2(_gnd_net_),
            .in3(N__13517),
            .lcout(Z_decfrac4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIE36D_0_5_LC_4_12_5.C_ON=1'b0;
    defparam counter_RNIE36D_0_5_LC_4_12_5.SEQ_MODE=4'b0000;
    defparam counter_RNIE36D_0_5_LC_4_12_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNIE36D_0_5_LC_4_12_5 (
            .in0(N__13855),
            .in1(N__16346),
            .in2(N__15974),
            .in3(N__13764),
            .lcout(voltage_011_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_2_LC_4_12_7.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_2_LC_4_12_7.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_2_LC_4_12_7.LUT_INIT=16'b1101110100010001;
    LogicCell40 slaveselect_RNILOQC2_2_LC_4_12_7 (
            .in0(N__13478),
            .in1(N__19290),
            .in2(_gnd_net_),
            .in3(N__13553),
            .lcout(slaveselect_RNILOQC2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_cry_1_c_LC_4_13_0.C_ON=1'b1;
    defparam counter_cry_1_c_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam counter_cry_1_c_LC_4_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 counter_cry_1_c_LC_4_13_0 (
            .in0(_gnd_net_),
            .in1(N__15810),
            .in2(N__16242),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_4_13_1.C_ON=1'b1;
    defparam counter_2_LC_4_13_1.SEQ_MODE=4'b1000;
    defparam counter_2_LC_4_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_4_13_1 (
            .in0(_gnd_net_),
            .in1(N__15935),
            .in2(_gnd_net_),
            .in3(N__12056),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(counter_cry_1),
            .carryout(counter_cry_2),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_3_LC_4_13_2.C_ON=1'b1;
    defparam counter_3_LC_4_13_2.SEQ_MODE=4'b1000;
    defparam counter_3_LC_4_13_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_4_13_2 (
            .in0(_gnd_net_),
            .in1(N__16393),
            .in2(_gnd_net_),
            .in3(N__12053),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(counter_cry_2),
            .carryout(counter_cry_3),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_4_LC_4_13_3.C_ON=1'b1;
    defparam counter_4_LC_4_13_3.SEQ_MODE=4'b1000;
    defparam counter_4_LC_4_13_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_4_13_3 (
            .in0(_gnd_net_),
            .in1(N__13862),
            .in2(_gnd_net_),
            .in3(N__12050),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(counter_cry_3),
            .carryout(counter_cry_4),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_5_LC_4_13_4.C_ON=1'b1;
    defparam counter_5_LC_4_13_4.SEQ_MODE=4'b1000;
    defparam counter_5_LC_4_13_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_5_LC_4_13_4 (
            .in0(_gnd_net_),
            .in1(N__13767),
            .in2(_gnd_net_),
            .in3(N__12125),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(counter_cry_4),
            .carryout(counter_cry_5),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_6_LC_4_13_5.C_ON=1'b1;
    defparam counter_6_LC_4_13_5.SEQ_MODE=4'b1000;
    defparam counter_6_LC_4_13_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_4_13_5 (
            .in0(_gnd_net_),
            .in1(N__13795),
            .in2(_gnd_net_),
            .in3(N__12122),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(counter_cry_5),
            .carryout(counter_cry_6),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_7_LC_4_13_6.C_ON=1'b1;
    defparam counter_7_LC_4_13_6.SEQ_MODE=4'b1000;
    defparam counter_7_LC_4_13_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_7_LC_4_13_6 (
            .in0(_gnd_net_),
            .in1(N__13898),
            .in2(_gnd_net_),
            .in3(N__12119),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(counter_cry_6),
            .carryout(counter_cry_7),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_8_LC_4_13_7.C_ON=1'b1;
    defparam counter_8_LC_4_13_7.SEQ_MODE=4'b1000;
    defparam counter_8_LC_4_13_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_8_LC_4_13_7 (
            .in0(_gnd_net_),
            .in1(N__13720),
            .in2(_gnd_net_),
            .in3(N__12116),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(counter_cry_7),
            .carryout(counter_cry_8),
            .clk(N__19970),
            .ce(),
            .sr(N__12102));
    defparam counter_9_LC_4_14_0.C_ON=1'b0;
    defparam counter_9_LC_4_14_0.SEQ_MODE=4'b1000;
    defparam counter_9_LC_4_14_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_9_LC_4_14_0 (
            .in0(_gnd_net_),
            .in1(N__13924),
            .in2(_gnd_net_),
            .in3(N__12113),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19973),
            .ce(),
            .sr(N__12109));
    defparam counter_0_LC_4_14_2.C_ON=1'b0;
    defparam counter_0_LC_4_14_2.SEQ_MODE=4'b1000;
    defparam counter_0_LC_4_14_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 counter_0_LC_4_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16150),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19973),
            .ce(),
            .sr(N__12109));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_3_0.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_3_0 (
            .in0(_gnd_net_),
            .in1(N__22611),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2579_LC_5_3_1.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2579_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2579_LC_5_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2579_LC_5_3_1 (
            .in0(_gnd_net_),
            .in1(N__12073),
            .in2(N__14048),
            .in3(N__12080),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTAS4_LC_5_3_2.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTAS4_LC_5_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTAS4_LC_5_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTAS4_LC_5_3_2 (
            .in0(_gnd_net_),
            .in1(N__14071),
            .in2(N__13658),
            .in3(N__12077),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_3_3.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_3_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_3_3 (
            .in0(N__14070),
            .in1(N__12074),
            .in2(N__14096),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKP36_LC_5_3_4.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKP36_LC_5_3_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKP36_LC_5_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKP36_LC_5_3_4 (
            .in0(_gnd_net_),
            .in1(N__14084),
            .in2(_gnd_net_),
            .in3(N__12245),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un173_pixellto5_LC_5_3_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un173_pixellto5_LC_5_3_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un173_pixellto5_LC_5_3_6.LUT_INIT=16'b1110010100001000;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un173_pixellto5_LC_5_3_6 (
            .in0(N__12227),
            .in1(N__23088),
            .in2(N__22622),
            .in3(N__12242),
            .lcout(chessboardpixel_un173_pixellt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un151_pixel_if_generate_plus_mult1_remainder_0_6_LC_5_3_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un151_pixel_if_generate_plus_mult1_remainder_0_6_LC_5_3_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un151_pixel_if_generate_plus_mult1_remainder_0_6_LC_5_3_7.LUT_INIT=16'b0011100111001100;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un151_pixel_if_generate_plus_mult1_remainder_0_6_LC_5_3_7 (
            .in0(N__12241),
            .in1(N__12233),
            .in2(N__22621),
            .in3(N__12226),
            .lcout(chessboardpixel_un151_pixel_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_0_LC_5_4_0.C_ON=1'b0;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_0_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_0_LC_5_4_0.LUT_INIT=16'b1111111101010101;
    LogicCell40 chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_0_LC_5_4_0 (
            .in0(N__12175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12193),
            .lcout(),
            .ltout(chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un177_pixel_if_generate_plus_mult1_remainder_0_5_LC_5_4_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un177_pixel_if_generate_plus_mult1_remainder_0_5_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un177_pixel_if_generate_plus_mult1_remainder_0_5_LC_5_4_1.LUT_INIT=16'b1010100110101010;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un177_pixel_if_generate_plus_mult1_remainder_0_5_LC_5_4_1 (
            .in0(N__12218),
            .in1(N__12185),
            .in2(N__12212),
            .in3(N__12151),
            .lcout(),
            .ltout(chessboardpixel_un177_pixel_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un174_pixel_LC_5_4_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un174_pixel_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un174_pixel_LC_5_4_2.LUT_INIT=16'b0001000100011110;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un174_pixel_LC_5_4_2 (
            .in0(N__12209),
            .in1(N__12203),
            .in2(N__12197),
            .in3(N__12131),
            .lcout(chessboardpixel_un174_pixel),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_1_LC_5_4_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_1_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_1_LC_5_4_5.LUT_INIT=16'b0010101001000000;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_1_LC_5_4_5 (
            .in0(N__12194),
            .in1(N__12173),
            .in2(N__12152),
            .in3(N__12184),
            .lcout(),
            .ltout(un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_LC_5_4_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_LC_5_4_6.LUT_INIT=16'b1001000000000000;
    LogicCell40 un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_LC_5_4_6 (
            .in0(N__12174),
            .in1(N__12150),
            .in2(N__12134),
            .in3(N__23231),
            .lcout(chessboardpixel_un199_pixellt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSyncZ0_LC_5_4_7.C_ON=1'b0;
    defparam VSyncZ0_LC_5_4_7.SEQ_MODE=4'b1000;
    defparam VSyncZ0_LC_5_4_7.LUT_INIT=16'b1111110111111111;
    LogicCell40 VSyncZ0_LC_5_4_7 (
            .in0(N__14207),
            .in1(N__14991),
            .in2(N__14930),
            .in3(N__12347),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21057),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_a3_0_3_LC_5_5_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_a3_0_3_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_a3_0_3_LC_5_5_2.LUT_INIT=16'b0001000100110011;
    LogicCell40 un113_pixel_4_0_15__g0_i_a3_0_3_LC_5_5_2 (
            .in0(N__23264),
            .in1(N__14838),
            .in2(_gnd_net_),
            .in3(N__20840),
            .lcout(),
            .ltout(un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_a3_0_LC_5_5_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_a3_0_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_a3_0_LC_5_5_3.LUT_INIT=16'b0000000001000000;
    LogicCell40 un113_pixel_4_0_15__g0_i_a3_0_LC_5_5_3 (
            .in0(N__14495),
            .in1(N__12314),
            .in2(N__12326),
            .in3(N__13013),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII8O41_9_LC_5_5_4.C_ON=1'b0;
    defparam beamY_RNII8O41_9_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNII8O41_9_LC_5_5_4.LUT_INIT=16'b0000000000000100;
    LogicCell40 beamY_RNII8O41_9_LC_5_5_4 (
            .in0(N__12478),
            .in1(N__18158),
            .in2(N__12722),
            .in3(N__18287),
            .lcout(beamY_RNII8O41Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_a3_0_4_LC_5_5_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_a3_0_4_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_a3_0_4_LC_5_5_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 un113_pixel_4_0_15__g0_i_a3_0_4_LC_5_5_5 (
            .in0(N__14696),
            .in1(N__14925),
            .in2(N__12929),
            .in3(N__14990),
            .lcout(un113_pixel_4_0_15__g0_i_a3_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_5_5_6.C_ON=1'b0;
    defparam beamY_1_LC_5_5_6.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_5_5_6.LUT_INIT=16'b0001001010101010;
    LogicCell40 beamY_1_LC_5_5_6 (
            .in0(N__23265),
            .in1(N__14125),
            .in2(N__24639),
            .in3(N__17519),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21055),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_5_6_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_5_6_0.LUT_INIT=16'b0100110111010011;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_5_6_0 (
            .in0(N__12668),
            .in1(N__18162),
            .in2(N__14039),
            .in3(N__18284),
            .lcout(if_generate_plus_mult1_un54_sum_axbxc5),
            .ltout(if_generate_plus_mult1_un54_sum_axbxc5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m4_0_LC_5_6_1.C_ON=1'b0;
    defparam row_1_if_m4_0_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam row_1_if_m4_0_LC_5_6_1.LUT_INIT=16'b0101011010010101;
    LogicCell40 row_1_if_m4_0_LC_5_6_1 (
            .in0(N__13263),
            .in1(N__12308),
            .in2(N__12302),
            .in3(N__12299),
            .lcout(),
            .ltout(row_1_if_i2_mux_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_ns_LC_5_6_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_ns_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_5_ns_LC_5_6_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_ac0_5_ns_LC_5_6_2 (
            .in0(_gnd_net_),
            .in1(N__12260),
            .in2(N__12254),
            .in3(N__12251),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_ac0_5),
            .ltout(row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x0_LC_5_6_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x0_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x0_LC_5_6_3.LUT_INIT=16'b1001000101100100;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_c5_x0_LC_5_6_3 (
            .in0(N__13264),
            .in1(N__14299),
            .in2(N__12779),
            .in3(N__12479),
            .lcout(if_generate_plus_mult1_un75_sum_c5_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x1_LC_5_6_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x1_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x1_LC_5_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x1_LC_5_6_4 (
            .in0(N__12480),
            .in1(N__13265),
            .in2(N__14310),
            .in3(N__12501),
            .lcout(if_generate_plus_mult1_un82_sum_axbxc5_0_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un5_beamx_4_LC_5_6_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un5_beamx_4_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un5_beamx_4_LC_5_6_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 un113_pixel_4_0_15__un5_beamx_4_LC_5_6_5 (
            .in0(_gnd_net_),
            .in1(N__13011),
            .in2(_gnd_net_),
            .in3(N__12921),
            .lcout(un1_beamy_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJNLC_9_LC_5_6_6.C_ON=1'b0;
    defparam beamY_RNIJNLC_9_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIJNLC_9_LC_5_6_6.LUT_INIT=16'b1001110111010101;
    LogicCell40 beamY_RNIJNLC_9_LC_5_6_6 (
            .in0(N__14989),
            .in1(N__14892),
            .in2(N__12775),
            .in3(N__14811),
            .lcout(beamY_RNIJNLCZ0Z_9),
            .ltout(beamY_RNIJNLCZ0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVGU01_9_LC_5_6_7.C_ON=1'b0;
    defparam beamY_RNIVGU01_9_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIVGU01_9_LC_5_6_7.LUT_INIT=16'b0011110011000011;
    LogicCell40 beamY_RNIVGU01_9_LC_5_6_7 (
            .in0(_gnd_net_),
            .in1(N__14032),
            .in2(N__12695),
            .in3(N__12669),
            .lcout(beamY_RNIVGU01Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIR51RF1_3_LC_5_7_0.C_ON=1'b0;
    defparam beamY_RNIR51RF1_3_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIR51RF1_3_LC_5_7_0.LUT_INIT=16'b0101000110111010;
    LogicCell40 beamY_RNIR51RF1_3_LC_5_7_0 (
            .in0(N__13307),
            .in1(N__12817),
            .in2(N__12557),
            .in3(N__13269),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV42D31_6_LC_5_7_1.C_ON=1'b0;
    defparam beamY_RNIV42D31_6_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIV42D31_6_LC_5_7_1.LUT_INIT=16'b1000011100011110;
    LogicCell40 beamY_RNIV42D31_6_LC_5_7_1 (
            .in0(N__13069),
            .in1(N__13055),
            .in2(N__12521),
            .in3(N__13045),
            .lcout(beamY_RNIV42D31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x0_LC_5_7_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x0_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x0_LC_5_7_2.LUT_INIT=16'b0110100110011001;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x0_LC_5_7_2 (
            .in0(N__12467),
            .in1(N__14303),
            .in2(N__12506),
            .in3(N__13266),
            .lcout(if_generate_plus_mult1_un82_sum_axbxc5_0_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x1_LC_5_7_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x1_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_x1_LC_5_7_3.LUT_INIT=16'b1110110111011110;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_c5_x1_LC_5_7_3 (
            .in0(N__13267),
            .in1(N__12505),
            .in2(N__14311),
            .in3(N__12468),
            .lcout(),
            .ltout(if_generate_plus_mult1_un75_sum_c5_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_ns_LC_5_7_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_ns_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_ns_LC_5_7_4.LUT_INIT=16'b1110001011100010;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_c5_ns_LC_5_7_4 (
            .in0(N__13082),
            .in1(N__14186),
            .in2(N__13073),
            .in3(_gnd_net_),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7SK1V_3_LC_5_7_5.C_ON=1'b0;
    defparam beamY_RNI7SK1V_3_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI7SK1V_3_LC_5_7_5.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI7SK1V_3_LC_5_7_5 (
            .in0(N__13068),
            .in1(N__13054),
            .in2(_gnd_net_),
            .in3(N__13044),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axbxc5_0),
            .ltout(chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDHF0F2_3_LC_5_7_6.C_ON=1'b0;
    defparam beamY_RNIDHF0F2_3_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIDHF0F2_3_LC_5_7_6.LUT_INIT=16'b0001111010110100;
    LogicCell40 beamY_RNIDHF0F2_3_LC_5_7_6 (
            .in0(N__13025),
            .in1(N__13174),
            .in2(N__13016),
            .in3(N__13268),
            .lcout(chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_beamylto6_LC_5_7_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_beamylto6_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_beamylto6_LC_5_7_7.LUT_INIT=16'b0000000010000000;
    LogicCell40 un113_pixel_4_0_15__un4_beamylto6_LC_5_7_7 (
            .in0(N__14695),
            .in1(N__13012),
            .in2(N__12928),
            .in3(N__14371),
            .lcout(un4_beamylt8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0VHAB1_3_LC_5_8_0.C_ON=1'b0;
    defparam beamY_RNI0VHAB1_3_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI0VHAB1_3_LC_5_8_0.LUT_INIT=16'b1110111010111011;
    LogicCell40 beamY_RNI0VHAB1_3_LC_5_8_0 (
            .in0(N__14471),
            .in1(N__13156),
            .in2(_gnd_net_),
            .in3(N__13305),
            .lcout(chary_if_generate_plus_mult1_un75_sum_c5_N_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPLAE31_4_LC_5_8_1.C_ON=1'b0;
    defparam beamY_RNIPLAE31_4_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIPLAE31_4_LC_5_8_1.LUT_INIT=16'b1010101001010101;
    LogicCell40 beamY_RNIPLAE31_4_LC_5_8_1 (
            .in0(N__12813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14694),
            .lcout(),
            .ltout(beamY_RNIPLAE31Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4TRT4_3_LC_5_8_2.C_ON=1'b0;
    defparam beamY_RNIN4TRT4_3_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4TRT4_3_LC_5_8_2.LUT_INIT=16'b0101001110101100;
    LogicCell40 beamY_RNIN4TRT4_3_LC_5_8_2 (
            .in0(N__14372),
            .in1(N__12836),
            .in2(N__12830),
            .in3(N__12827),
            .lcout(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVGVF22_3_LC_5_8_3.C_ON=1'b0;
    defparam beamY_RNIVGVF22_3_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIVGVF22_3_LC_5_8_3.LUT_INIT=16'b0101101010100101;
    LogicCell40 beamY_RNIVGVF22_3_LC_5_8_3 (
            .in0(N__13157),
            .in1(_gnd_net_),
            .in2(N__12821),
            .in3(N__14472),
            .lcout(chary_if_generate_plus_mult1_un1_sum_axbxc3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_1_LC_5_8_4.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_1_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_1_LC_5_8_4.LUT_INIT=16'b0010010000011000;
    LogicCell40 un113_pixel_3_0_11__g0_1_LC_5_8_4 (
            .in0(N__13133),
            .in1(N__12791),
            .in2(N__20858),
            .in3(N__12785),
            .lcout(un113_pixel_3_0_11__g1_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_1_3_LC_5_8_5.C_ON=1'b0;
    defparam beamY_RNIHUG2_1_3_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_1_3_LC_5_8_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIHUG2_1_3_LC_5_8_5 (
            .in0(_gnd_net_),
            .in1(N__14470),
            .in2(_gnd_net_),
            .in3(N__20826),
            .lcout(un4_beamylt6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_2_LC_5_8_6.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_2_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_2_LC_5_8_6.LUT_INIT=16'b1001011000000000;
    LogicCell40 un113_pixel_3_0_11__g0_2_LC_5_8_6 (
            .in0(N__20827),
            .in1(N__13271),
            .in2(N__14487),
            .in3(N__13306),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_0_x2_0_0_LC_5_8_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_0_x2_0_0_LC_5_8_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_0_x2_0_0_LC_5_8_7.LUT_INIT=16'b0101001110101100;
    LogicCell40 un113_pixel_3_0_11__g0_0_x2_0_0_LC_5_8_7 (
            .in0(N__13272),
            .in1(N__13175),
            .in2(N__13163),
            .in3(N__13160),
            .lcout(un113_pixel_3_0_11__g0_0_x2_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_0_LC_5_9_0.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_0_LC_5_9_0.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_1_e_0_0_LC_5_9_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 ScreenBuffer_1_1_e_0_0_LC_5_9_0 (
            .in0(N__15344),
            .in1(N__15379),
            .in2(_gnd_net_),
            .in3(N__19305),
            .lcout(ScreenBuffer_1_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19963),
            .ce(N__13127),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_2_LC_5_9_1.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_2_LC_5_9_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_1_e_0_2_LC_5_9_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_1_e_0_2_LC_5_9_1 (
            .in0(N__19303),
            .in1(N__15261),
            .in2(_gnd_net_),
            .in3(N__15294),
            .lcout(ScreenBuffer_1_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19963),
            .ce(N__13127),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_3_LC_5_9_2.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_3_LC_5_9_2.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_1_e_0_3_LC_5_9_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 ScreenBuffer_1_1_e_0_3_LC_5_9_2 (
            .in0(N__15224),
            .in1(N__19304),
            .in2(_gnd_net_),
            .in3(N__15176),
            .lcout(ScreenBuffer_1_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19963),
            .ce(N__13127),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_1_LC_5_9_3.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_1_LC_5_9_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_1_e_0_1_LC_5_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 ScreenBuffer_1_1_e_0_1_LC_5_9_3 (
            .in0(N__19302),
            .in1(N__15129),
            .in2(_gnd_net_),
            .in3(N__15100),
            .lcout(ScreenBuffer_1_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19963),
            .ce(N__13127),
            .sr(_gnd_net_));
    defparam voltage_0_RNIVS2M_0_1_LC_5_9_4.C_ON=1'b0;
    defparam voltage_0_RNIVS2M_0_1_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam voltage_0_RNIVS2M_0_1_LC_5_9_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 voltage_0_RNIVS2M_0_1_LC_5_9_4 (
            .in0(N__15128),
            .in1(N__19047),
            .in2(_gnd_net_),
            .in3(N__15836),
            .lcout(N_1520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_voltage_2_1_cry_0_c_RNO_LC_5_10_1.C_ON=1'b0;
    defparam un1_voltage_2_1_cry_0_c_RNO_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam un1_voltage_2_1_cry_0_c_RNO_LC_5_10_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 un1_voltage_2_1_cry_0_c_RNO_LC_5_10_1 (
            .in0(N__20218),
            .in1(N__19280),
            .in2(N__15389),
            .in3(N__13468),
            .lcout(un1_voltage_2_1_cry_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_RNO_0_0_LC_5_10_2.C_ON=1'b0;
    defparam voltage_2_RNO_0_0_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam voltage_2_RNO_0_0_LC_5_10_2.LUT_INIT=16'b0111111110000000;
    LogicCell40 voltage_2_RNO_0_0_LC_5_10_2 (
            .in0(N__13469),
            .in1(N__20219),
            .in2(N__19327),
            .in3(N__15375),
            .lcout(),
            .ltout(un1_voltage_2_1_axb_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_2_0_LC_5_10_3.C_ON=1'b0;
    defparam voltage_2_0_LC_5_10_3.SEQ_MODE=4'b1000;
    defparam voltage_2_0_LC_5_10_3.LUT_INIT=16'b0011001111110011;
    LogicCell40 voltage_2_0_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(N__13451),
            .in2(N__13442),
            .in3(N__13412),
            .lcout(voltage_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19965),
            .ce(),
            .sr(N__18546));
    defparam voltage_2_2_LC_5_10_4.C_ON=1'b0;
    defparam voltage_2_2_LC_5_10_4.SEQ_MODE=4'b1000;
    defparam voltage_2_2_LC_5_10_4.LUT_INIT=16'b0111011100110011;
    LogicCell40 voltage_2_2_LC_5_10_4 (
            .in0(N__13414),
            .in1(N__13439),
            .in2(_gnd_net_),
            .in3(N__13433),
            .lcout(voltage_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19965),
            .ce(),
            .sr(N__18546));
    defparam voltage_2_1_LC_5_10_6.C_ON=1'b0;
    defparam voltage_2_1_LC_5_10_6.SEQ_MODE=4'b1000;
    defparam voltage_2_1_LC_5_10_6.LUT_INIT=16'b0111011100110011;
    LogicCell40 voltage_2_1_LC_5_10_6 (
            .in0(N__13413),
            .in1(N__13397),
            .in2(_gnd_net_),
            .in3(N__13388),
            .lcout(voltage_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19965),
            .ce(),
            .sr(N__18546));
    defparam voltage_0_RNI1V2M_2_LC_5_10_7.C_ON=1'b0;
    defparam voltage_0_RNI1V2M_2_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam voltage_0_RNI1V2M_2_LC_5_10_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 voltage_0_RNI1V2M_2_LC_5_10_7 (
            .in0(N__15286),
            .in1(N__16555),
            .in2(_gnd_net_),
            .in3(N__15817),
            .lcout(N_1505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_1_c_LC_5_11_0.C_ON=1'b1;
    defparam un42_cry_1_c_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam un42_cry_1_c_LC_5_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un42_cry_1_c_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(N__13376),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(un42_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_2_c_LC_5_11_1.C_ON=1'b1;
    defparam un42_cry_2_c_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam un42_cry_2_c_LC_5_11_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un42_cry_2_c_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(N__21912),
            .in2(N__15485),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un42_cry_1),
            .carryout(un42_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_3_c_LC_5_11_2.C_ON=1'b1;
    defparam un42_cry_3_c_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam un42_cry_3_c_LC_5_11_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un42_cry_3_c_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(N__13370),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un42_cry_2),
            .carryout(un42_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_3_c_RNIMRT41_LC_5_11_3.C_ON=1'b0;
    defparam un42_cry_3_c_RNIMRT41_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam un42_cry_3_c_RNIMRT41_LC_5_11_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 un42_cry_3_c_RNIMRT41_LC_5_11_3 (
            .in0(N__13358),
            .in1(N__13598),
            .in2(_gnd_net_),
            .in3(N__13352),
            .lcout(voltage_011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_4_LC_5_11_4.C_ON=1'b0;
    defparam ScreenBuffer_1_3_4_LC_5_11_4.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_3_4_LC_5_11_4.LUT_INIT=16'b1101110100010001;
    LogicCell40 ScreenBuffer_1_3_4_LC_5_11_4 (
            .in0(N__19306),
            .in1(N__15458),
            .in2(_gnd_net_),
            .in3(N__17332),
            .lcout(ScreenBuffer_1_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19968),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_2_0_LC_5_11_5.C_ON=1'b0;
    defparam ScreenBuffer_0_2_0_LC_5_11_5.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_2_0_LC_5_11_5.LUT_INIT=16'b1011100011110000;
    LogicCell40 ScreenBuffer_0_2_0_LC_5_11_5 (
            .in0(N__20205),
            .in1(N__13487),
            .in2(N__17210),
            .in3(N__19307),
            .lcout(ScreenBuffer_0_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19968),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_LC_5_11_7.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_LC_5_11_7.LUT_INIT=16'b1011101100010001;
    LogicCell40 slaveselect_RNILOQC2_LC_5_11_7 (
            .in0(N__19289),
            .in1(N__13486),
            .in2(_gnd_net_),
            .in3(N__13561),
            .lcout(slaveselect_RNILOQCZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIE36D_5_LC_5_12_0.C_ON=1'b0;
    defparam counter_RNIE36D_5_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam counter_RNIE36D_5_LC_5_12_0.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIE36D_5_LC_5_12_0 (
            .in0(N__13859),
            .in1(N__16360),
            .in2(N__15975),
            .in3(N__13765),
            .lcout(ScreenBuffer_1_122_1),
            .ltout(ScreenBuffer_1_122_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNITIV01_0_LC_5_12_1.C_ON=1'b0;
    defparam counter_RNITIV01_0_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam counter_RNITIV01_0_LC_5_12_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 counter_RNITIV01_0_LC_5_12_1 (
            .in0(N__13594),
            .in1(N__16216),
            .in2(N__13490),
            .in3(N__15832),
            .lcout(ScreenBuffer_1_3_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNITIV01_2_0_LC_5_12_2.C_ON=1'b0;
    defparam counter_RNITIV01_2_0_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam counter_RNITIV01_2_0_LC_5_12_2.LUT_INIT=16'b0000010000000000;
    LogicCell40 counter_RNITIV01_2_0_LC_5_12_2 (
            .in0(N__16215),
            .in1(N__13612),
            .in2(N__15854),
            .in3(N__13596),
            .lcout(ScreenBuffer_1_0_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_1_0_LC_5_12_3.C_ON=1'b0;
    defparam ScreenBuffer_0_1_0_LC_5_12_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_1_0_LC_5_12_3.LUT_INIT=16'b1111100001110000;
    LogicCell40 ScreenBuffer_0_1_0_LC_5_12_3 (
            .in0(N__19301),
            .in1(N__13571),
            .in2(N__16979),
            .in3(N__20203),
            .lcout(ScreenBuffer_0_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19971),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNITIV01_1_0_LC_5_12_4.C_ON=1'b0;
    defparam counter_RNITIV01_1_0_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam counter_RNITIV01_1_0_LC_5_12_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 counter_RNITIV01_1_0_LC_5_12_4 (
            .in0(N__16217),
            .in1(N__13611),
            .in2(N__15855),
            .in3(N__13595),
            .lcout(ScreenBuffer_1_1_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_4_RNO_0_0_LC_5_12_6.C_ON=1'b0;
    defparam ScreenBuffer_0_4_RNO_0_0_LC_5_12_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_4_RNO_0_0_LC_5_12_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 ScreenBuffer_0_4_RNO_0_0_LC_5_12_6 (
            .in0(_gnd_net_),
            .in1(N__19300),
            .in2(_gnd_net_),
            .in3(N__13467),
            .lcout(),
            .ltout(un1_sclk17_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_4_0_LC_5_12_7.C_ON=1'b0;
    defparam ScreenBuffer_0_4_0_LC_5_12_7.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_4_0_LC_5_12_7.LUT_INIT=16'b1110101000101010;
    LogicCell40 ScreenBuffer_0_4_0_LC_5_12_7 (
            .in0(N__18958),
            .in1(N__16498),
            .in2(N__13646),
            .in3(N__20204),
            .lcout(ScreenBuffer_0_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19971),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIUJ6D_9_LC_5_13_0.C_ON=1'b0;
    defparam counter_RNIUJ6D_9_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam counter_RNIUJ6D_9_LC_5_13_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 counter_RNIUJ6D_9_LC_5_13_0 (
            .in0(N__13922),
            .in1(N__13718),
            .in2(_gnd_net_),
            .in3(N__13642),
            .lcout(un39_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIT7J6_6_LC_5_13_1.C_ON=1'b0;
    defparam counter_RNIT7J6_6_LC_5_13_1.SEQ_MODE=4'b0000;
    defparam counter_RNIT7J6_6_LC_5_13_1.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_RNIT7J6_6_LC_5_13_1 (
            .in0(_gnd_net_),
            .in1(N__13895),
            .in2(_gnd_net_),
            .in3(N__13793),
            .lcout(un39_0_3),
            .ltout(un39_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIB6GG_9_LC_5_13_2.C_ON=1'b0;
    defparam counter_RNIB6GG_9_LC_5_13_2.SEQ_MODE=4'b0000;
    defparam counter_RNIB6GG_9_LC_5_13_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNIB6GG_9_LC_5_13_2 (
            .in0(N__13921),
            .in1(N__13717),
            .in2(N__13628),
            .in3(N__13763),
            .lcout(un5_slaveselect_1),
            .ltout(un5_slaveselect_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNITIV01_4_LC_5_13_3.C_ON=1'b0;
    defparam counter_RNITIV01_4_LC_5_13_3.SEQ_MODE=4'b0000;
    defparam counter_RNITIV01_4_LC_5_13_3.LUT_INIT=16'b1010000011110000;
    LogicCell40 counter_RNITIV01_4_LC_5_13_3 (
            .in0(N__13874),
            .in1(_gnd_net_),
            .in2(N__13616),
            .in3(N__13860),
            .lcout(un10_slaveselect),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNITIV01_0_0_LC_5_13_4.C_ON=1'b0;
    defparam counter_RNITIV01_0_0_LC_5_13_4.SEQ_MODE=4'b0000;
    defparam counter_RNITIV01_0_0_LC_5_13_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 counter_RNITIV01_0_0_LC_5_13_4 (
            .in0(N__13613),
            .in1(N__13597),
            .in2(N__16241),
            .in3(N__15818),
            .lcout(ScreenBuffer_1_2_1_sqmuxa),
            .ltout(ScreenBuffer_1_2_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_0_LC_5_13_5.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_0_LC_5_13_5.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_0_LC_5_13_5.LUT_INIT=16'b1100111100000011;
    LogicCell40 slaveselect_RNILOQC2_0_LC_5_13_5 (
            .in0(_gnd_net_),
            .in1(N__19329),
            .in2(N__13565),
            .in3(N__13554),
            .lcout(slaveselect_RNILOQC2Z0Z_0),
            .ltout(slaveselect_RNILOQC2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_5_LC_5_13_6.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_5_LC_5_13_6.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_5_LC_5_13_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 slaveselect_RNILOQC2_5_LC_5_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13520),
            .in3(_gnd_net_),
            .lcout(un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIAAPJ_7_LC_5_13_7.C_ON=1'b0;
    defparam counter_RNIAAPJ_7_LC_5_13_7.SEQ_MODE=4'b0000;
    defparam counter_RNIAAPJ_7_LC_5_13_7.LUT_INIT=16'b0000000000001000;
    LogicCell40 counter_RNIAAPJ_7_LC_5_13_7 (
            .in0(N__13516),
            .in1(N__13811),
            .in2(N__13928),
            .in3(N__13896),
            .lcout(slaveselect_1lto9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIEUS9_6_LC_5_14_1.C_ON=1'b0;
    defparam counter_RNIEUS9_6_LC_5_14_1.SEQ_MODE=4'b0000;
    defparam counter_RNIEUS9_6_LC_5_14_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 counter_RNIEUS9_6_LC_5_14_1 (
            .in0(N__13923),
            .in1(N__13897),
            .in2(_gnd_net_),
            .in3(N__13794),
            .lcout(),
            .ltout(un1_counter_1lto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI283N_8_LC_5_14_2.C_ON=1'b0;
    defparam counter_RNI283N_8_LC_5_14_2.SEQ_MODE=4'b0000;
    defparam counter_RNI283N_8_LC_5_14_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 counter_RNI283N_8_LC_5_14_2 (
            .in0(N__13810),
            .in1(N__13719),
            .in2(N__13877),
            .in3(N__13766),
            .lcout(un1_counter_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_6_0_LC_5_14_4.C_ON=1'b0;
    defparam ScreenBuffer_0_6_0_LC_5_14_4.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_6_0_LC_5_14_4.LUT_INIT=16'b1111100001110000;
    LogicCell40 ScreenBuffer_0_6_0_LC_5_14_4 (
            .in0(N__16520),
            .in1(N__16507),
            .in2(N__18940),
            .in3(N__20199),
            .lcout(ScreenBuffer_0_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19977),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_2_3_LC_5_14_6.C_ON=1'b0;
    defparam counter_RNI6R5D_2_3_LC_5_14_6.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_2_3_LC_5_14_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNI6R5D_2_3_LC_5_14_6 (
            .in0(N__16344),
            .in1(N__15923),
            .in2(N__15861),
            .in3(N__16109),
            .lcout(un10_slaveselectlt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIN1J6_4_LC_5_14_7.C_ON=1'b0;
    defparam counter_RNIN1J6_4_LC_5_14_7.SEQ_MODE=4'b0000;
    defparam counter_RNIN1J6_4_LC_5_14_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_RNIN1J6_4_LC_5_14_7 (
            .in0(_gnd_net_),
            .in1(N__13861),
            .in2(_gnd_net_),
            .in3(N__16345),
            .lcout(un1_counter_1lt9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIBRS9_6_LC_5_15_6.C_ON=1'b0;
    defparam counter_RNIBRS9_6_LC_5_15_6.SEQ_MODE=4'b0000;
    defparam counter_RNIBRS9_6_LC_5_15_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 counter_RNIBRS9_6_LC_5_15_6 (
            .in0(N__13799),
            .in1(N__13772),
            .in2(_gnd_net_),
            .in3(N__13724),
            .lcout(slaveselect_1lto9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNIIRSC1_LC_5_16_5.C_ON=1'b0;
    defparam slaveselect_RNIIRSC1_LC_5_16_5.SEQ_MODE=4'b0000;
    defparam slaveselect_RNIIRSC1_LC_5_16_5.LUT_INIT=16'b1111100011111111;
    LogicCell40 slaveselect_RNIIRSC1_LC_5_16_5 (
            .in0(N__13694),
            .in1(N__13685),
            .in2(N__19997),
            .in3(N__19330),
            .lcout(SCLK1_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0 (
            .in0(_gnd_net_),
            .in1(N__22462),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJE1_LC_6_2_1.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJE1_LC_6_2_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJE1_LC_6_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJE1_LC_6_2_1 (
            .in0(_gnd_net_),
            .in1(N__14056),
            .in2(N__16610),
            .in3(N__13649),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LB2_LC_6_2_2.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LB2_LC_6_2_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LB2_LC_6_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LB2_LC_6_2_2 (
            .in0(_gnd_net_),
            .in1(N__16630),
            .in2(N__16667),
            .in3(N__14087),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGAHS5_LC_6_2_3.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGAHS5_LC_6_2_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGAHS5_LC_6_2_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGAHS5_LC_6_2_3 (
            .in0(N__14072),
            .in1(N__14057),
            .in2(N__16655),
            .in3(N__14078),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3H63_LC_6_2_4.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3H63_LC_6_2_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3H63_LC_6_2_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3H63_LC_6_2_4 (
            .in0(_gnd_net_),
            .in1(N__16643),
            .in2(_gnd_net_),
            .in3(N__14075),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_0_LC_6_2_6.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_0_LC_6_2_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_0_LC_6_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_0_LC_6_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16629),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_6_3_2.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_6_3_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22459),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_6_3_5.C_ON=1'b0;
    defparam beamX_0_LC_6_3_5.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_6_3_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_0_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(N__17529),
            .in2(_gnd_net_),
            .in3(N__18698),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21059),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_3_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_3_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un5_beamx_2_0_LC_6_4_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un5_beamx_2_0_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un5_beamx_2_0_LC_6_4_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 un113_pixel_4_0_15__un5_beamx_2_0_LC_6_4_3 (
            .in0(N__23232),
            .in1(N__15002),
            .in2(_gnd_net_),
            .in3(N__14837),
            .lcout(un113_pixel_4_0_15__un5_beamx_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_row_2_LC_6_5_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_row_2_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_row_2_LC_6_5_0.LUT_INIT=16'b1100000001110000;
    LogicCell40 un113_pixel_4_0_15__un4_row_2_LC_6_5_0 (
            .in0(N__14038),
            .in1(N__18168),
            .in2(N__18041),
            .in3(N__18292),
            .lcout(un113_pixel_4_0_15__un4_rowZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un5_beamx_4_0_LC_6_5_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un5_beamx_4_0_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un5_beamx_4_0_LC_6_5_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 un113_pixel_4_0_15__un5_beamx_4_0_LC_6_5_2 (
            .in0(N__14700),
            .in1(N__14494),
            .in2(N__14929),
            .in3(N__20883),
            .lcout(),
            .ltout(un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un5_beamx_LC_6_5_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un5_beamx_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un5_beamx_LC_6_5_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 un113_pixel_4_0_15__un5_beamx_LC_6_5_3 (
            .in0(N__14156),
            .in1(N__24593),
            .in2(N__14150),
            .in3(N__14203),
            .lcout(un5_beamx_0),
            .ltout(un5_beamx_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_6_5_4.C_ON=1'b0;
    defparam beamY_0_LC_6_5_4.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_6_5_4.LUT_INIT=16'b0000010110101010;
    LogicCell40 beamY_0_LC_6_5_4 (
            .in0(N__24594),
            .in1(_gnd_net_),
            .in2(N__14111),
            .in3(N__17533),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21058),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un3_beamx_5_LC_6_5_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un3_beamx_5_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un3_beamx_5_LC_6_5_5.LUT_INIT=16'b0001000000000000;
    LogicCell40 un113_pixel_4_0_15__un3_beamx_5_LC_6_5_5 (
            .in0(N__17867),
            .in1(N__17902),
            .in2(N__17790),
            .in3(N__17466),
            .lcout(),
            .ltout(un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un3_beamx_7_LC_6_5_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un3_beamx_7_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un3_beamx_7_LC_6_5_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 un113_pixel_4_0_15__un3_beamx_7_LC_6_5_6 (
            .in0(N__17830),
            .in1(N__18704),
            .in2(N__14108),
            .in3(N__17686),
            .lcout(un113_pixel_4_0_15__un3_beamxZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un13_beamylto3_LC_6_5_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un13_beamylto3_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un13_beamylto3_LC_6_5_7.LUT_INIT=16'b0000000001111111;
    LogicCell40 un113_pixel_4_0_15__un13_beamylto3_LC_6_5_7 (
            .in0(N__17866),
            .in1(N__17901),
            .in2(N__18720),
            .in3(N__17829),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un13_beamylto10_LC_6_6_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un13_beamylto10_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un13_beamylto10_LC_6_6_0.LUT_INIT=16'b0011011100000000;
    LogicCell40 un113_pixel_4_0_15__un13_beamylto10_LC_6_6_0 (
            .in0(N__14105),
            .in1(N__17614),
            .in2(N__17687),
            .in3(N__16805),
            .lcout(un13_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un13_beamylto5_LC_6_6_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un13_beamylto5_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un13_beamylto5_LC_6_6_1.LUT_INIT=16'b0100010000000000;
    LogicCell40 un113_pixel_4_0_15__un13_beamylto5_LC_6_6_1 (
            .in0(N__14335),
            .in1(N__17726),
            .in2(_gnd_net_),
            .in3(N__17783),
            .lcout(un13_beamylt6_0),
            .ltout(un13_beamylt6_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_6_LC_6_6_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_6_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_6_LC_6_6_2.LUT_INIT=16'b0011011100000000;
    LogicCell40 un113_pixel_4_0_15__g0_6_LC_6_6_2 (
            .in0(N__17684),
            .in1(N__17615),
            .in2(N__14099),
            .in3(N__16806),
            .lcout(un13_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un18_beamylto9_LC_6_6_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un18_beamylto9_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un18_beamylto9_LC_6_6_3.LUT_INIT=16'b1101110000000000;
    LogicCell40 un113_pixel_4_0_15__un18_beamylto9_LC_6_6_3 (
            .in0(N__14336),
            .in1(N__17727),
            .in2(N__17792),
            .in3(N__16841),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_row_5_LC_6_6_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_row_5_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_row_5_LC_6_6_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 un113_pixel_4_0_15__un4_row_5_LC_6_6_4 (
            .in0(N__14327),
            .in1(N__14321),
            .in2(N__14315),
            .in3(N__20576),
            .lcout(un113_pixel_4_0_15__un4_rowZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un3_beamx_LC_6_6_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un3_beamx_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un3_beamx_LC_6_6_5.LUT_INIT=16'b0000000000001000;
    LogicCell40 un113_pixel_4_0_15__un3_beamx_LC_6_6_5 (
            .in0(N__16807),
            .in1(N__14249),
            .in2(N__17621),
            .in3(N__17728),
            .lcout(un3_beamx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un1_beamxlto6_LC_6_6_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un1_beamxlto6_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un1_beamxlto6_LC_6_6_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 un113_pixel_4_0_15__un1_beamxlto6_LC_6_6_6 (
            .in0(N__17729),
            .in1(N__17685),
            .in2(N__17791),
            .in3(N__17834),
            .lcout(),
            .ltout(un1_beamxlt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSyncZ0_LC_6_6_7.C_ON=1'b0;
    defparam HSyncZ0_LC_6_6_7.SEQ_MODE=4'b1000;
    defparam HSyncZ0_LC_6_6_7.LUT_INIT=16'b1111111111111101;
    LogicCell40 HSyncZ0_LC_6_6_7 (
            .in0(N__16808),
            .in1(N__17619),
            .in2(N__14243),
            .in3(N__17467),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21056),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un15_beamy_2_LC_6_7_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un15_beamy_2_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un15_beamy_2_LC_6_7_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 un113_pixel_4_0_15__un15_beamy_2_LC_6_7_1 (
            .in0(N__14714),
            .in1(N__17468),
            .in2(N__14552),
            .in3(N__14225),
            .lcout(un113_pixel_4_0_15__un15_beamyZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_ns_LC_6_7_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_ns_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_ns_LC_6_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_ns_LC_6_7_4 (
            .in0(N__14184),
            .in1(N__14219),
            .in2(_gnd_net_),
            .in3(N__14213),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un8_beamylto9_1_LC_6_7_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un8_beamylto9_1_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un8_beamylto9_1_LC_6_7_5.LUT_INIT=16'b0000000100000000;
    LogicCell40 un113_pixel_4_0_15__un8_beamylto9_1_LC_6_7_5 (
            .in0(N__14983),
            .in1(N__14920),
            .in2(N__14845),
            .in3(N__14202),
            .lcout(un113_pixel_4_0_15__un8_beamylto9Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_row_LC_6_7_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_row_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_row_LC_6_7_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 un113_pixel_4_0_15__un4_row_LC_6_7_6 (
            .in0(N__14185),
            .in1(N__23615),
            .in2(N__14165),
            .in3(N__23108),
            .lcout(un4_row),
            .ltout(un4_row_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_5_LC_6_7_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_5_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_5_LC_6_7_7.LUT_INIT=16'b0000010000000000;
    LogicCell40 un113_pixel_4_0_15__g0_5_LC_6_7_7 (
            .in0(N__15023),
            .in1(N__15014),
            .in2(N__15005),
            .in3(N__16937),
            .lcout(Pixel_3_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_beamylto9_LC_6_8_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_beamylto9_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_beamylto9_LC_6_8_0.LUT_INIT=16'b1010101010101000;
    LogicCell40 un113_pixel_4_0_15__un4_beamylto9_LC_6_8_0 (
            .in0(N__14998),
            .in1(N__14921),
            .in2(N__14846),
            .in3(N__14720),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un8_beamylto9_LC_6_8_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un8_beamylto9_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un8_beamylto9_LC_6_8_2.LUT_INIT=16'b0010101010101010;
    LogicCell40 un113_pixel_4_0_15__un8_beamylto9_LC_6_8_2 (
            .in0(N__14708),
            .in1(N__20886),
            .in2(N__14702),
            .in3(N__14478),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_a9_LC_6_8_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_a9_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_a9_LC_6_8_3.LUT_INIT=16'b0000001100100001;
    LogicCell40 un113_pixel_4_0_15__g0_i_a9_LC_6_8_3 (
            .in0(N__20888),
            .in1(N__23244),
            .in2(N__14540),
            .in3(N__20677),
            .lcout(N_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_x4_0_LC_6_8_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_x4_0_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_x4_0_LC_6_8_4.LUT_INIT=16'b0101010110101010;
    LogicCell40 un113_pixel_4_0_15__g0_i_x4_0_LC_6_8_4 (
            .in0(N__20924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20966),
            .lcout(N_6_i),
            .ltout(N_6_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_a9_0_LC_6_8_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_a9_0_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_a9_0_LC_6_8_5.LUT_INIT=16'b1000000001000000;
    LogicCell40 un113_pixel_4_0_15__g0_i_a9_0_LC_6_8_5 (
            .in0(N__20887),
            .in1(N__23243),
            .in2(N__14531),
            .in3(N__20676),
            .lcout(N_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m2_2_LC_6_8_6.C_ON=1'b0;
    defparam row_1_if_m2_2_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam row_1_if_m2_2_LC_6_8_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 row_1_if_m2_2_LC_6_8_6 (
            .in0(N__17251),
            .in1(N__14528),
            .in2(_gnd_net_),
            .in3(N__14477),
            .lcout(),
            .ltout(if_m2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_6_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_6_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_6_8_7.LUT_INIT=16'b0111010010001011;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_6_8_7 (
            .in0(N__14370),
            .in1(N__14354),
            .in2(N__14345),
            .in3(N__14342),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_6_9_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_6_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__16876),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PA3_LC_6_9_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PA3_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PA3_LC_6_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PA3_LC_6_9_1 (
            .in0(_gnd_net_),
            .in1(N__16793),
            .in2(_gnd_net_),
            .in3(N__15056),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PA3_LC_6_9_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PA3_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PA3_LC_6_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PA3_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__16904),
            .in2(N__21888),
            .in3(N__15053),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_6_9_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_6_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_6_9_3 (
            .in0(_gnd_net_),
            .in1(N__16888),
            .in2(_gnd_net_),
            .in3(N__15050),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_6_9_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_6_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15047),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_0_LC_6_9_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_0_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_0_LC_6_9_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_0_LC_6_9_7 (
            .in0(N__16877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_6_10_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_6_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17077),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBS1_LC_6_10_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBS1_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBS1_LC_6_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBS1_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(N__15419),
            .in2(N__15044),
            .in3(N__15035),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5B3_LC_6_10_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5B3_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5B3_LC_6_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5B3_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(N__15032),
            .in2(N__15410),
            .in3(N__15026),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_6_10_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_6_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_6_10_3 (
            .in0(_gnd_net_),
            .in1(N__15434),
            .in2(N__15443),
            .in3(N__15405),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5B3_LC_6_10_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5B3_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5B3_LC_6_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5B3_LC_6_10_4 (
            .in0(N__15409),
            .in1(N__15428),
            .in2(N__16898),
            .in3(N__15422),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_6_10_5.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_6_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15418),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_5_1_LC_6_10_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_5_1_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_5_1_LC_6_10_6.LUT_INIT=16'b1111111011111101;
    LogicCell40 un113_pixel_4_0_15__g0_5_1_LC_6_10_6 (
            .in0(N__17073),
            .in1(N__20996),
            .in2(N__18736),
            .in3(N__17117),
            .lcout(un113_pixel_4_0_15__g0_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_e_0_0_LC_6_11_0.C_ON=1'b0;
    defparam ScreenBuffer_1_2_e_0_0_LC_6_11_0.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_2_e_0_0_LC_6_11_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_2_e_0_0_LC_6_11_0 (
            .in0(N__19319),
            .in1(N__15380),
            .in2(_gnd_net_),
            .in3(N__15343),
            .lcout(ScreenBuffer_1_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19972),
            .ce(N__15068),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_e_0_2_LC_6_11_1.C_ON=1'b0;
    defparam ScreenBuffer_1_2_e_0_2_LC_6_11_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_2_e_0_2_LC_6_11_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 ScreenBuffer_1_2_e_0_2_LC_6_11_1 (
            .in0(N__15293),
            .in1(N__19322),
            .in2(_gnd_net_),
            .in3(N__15263),
            .lcout(ScreenBuffer_1_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19972),
            .ce(N__15068),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_e_0_3_LC_6_11_2.C_ON=1'b0;
    defparam ScreenBuffer_1_2_e_0_3_LC_6_11_2.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_2_e_0_3_LC_6_11_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_2_e_0_3_LC_6_11_2 (
            .in0(N__19320),
            .in1(N__15223),
            .in2(_gnd_net_),
            .in3(N__15175),
            .lcout(ScreenBuffer_1_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19972),
            .ce(N__15068),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_e_0_1_LC_6_11_3.C_ON=1'b0;
    defparam ScreenBuffer_1_2_e_0_1_LC_6_11_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_2_e_0_1_LC_6_11_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 ScreenBuffer_1_2_e_0_1_LC_6_11_3 (
            .in0(N__15135),
            .in1(N__19321),
            .in2(_gnd_net_),
            .in3(N__15099),
            .lcout(ScreenBuffer_1_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19972),
            .ce(N__15068),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_15_LC_6_11_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_15_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_15_LC_6_11_4.LUT_INIT=16'b1001100111001100;
    LogicCell40 un113_pixel_4_0_15__g0_15_LC_6_11_4 (
            .in0(N__17078),
            .in1(N__21159),
            .in2(_gnd_net_),
            .in3(N__17118),
            .lcout(font_un3_pixel_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un42_cry_2_c_RNO_LC_6_11_5.C_ON=1'b0;
    defparam un42_cry_2_c_RNO_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam un42_cry_2_c_RNO_LC_6_11_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 un42_cry_2_c_RNO_LC_6_11_5 (
            .in0(N__15532),
            .in1(N__16245),
            .in2(_gnd_net_),
            .in3(N__15520),
            .lcout(un42_cry_2_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_11_RNO_0_0_LC_6_12_0.C_ON=1'b0;
    defparam ScreenBuffer_0_11_RNO_0_0_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_11_RNO_0_0_LC_6_12_0.LUT_INIT=16'b0000000100000000;
    LogicCell40 ScreenBuffer_0_11_RNO_0_0_LC_6_12_0 (
            .in0(N__16274),
            .in1(N__15980),
            .in2(N__16426),
            .in3(N__19249),
            .lcout(),
            .ltout(un1_sclk17_6_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_11_0_LC_6_12_1.C_ON=1'b0;
    defparam ScreenBuffer_0_11_0_LC_6_12_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_11_0_LC_6_12_1.LUT_INIT=16'b1101111110000000;
    LogicCell40 ScreenBuffer_0_11_0_LC_6_12_1 (
            .in0(N__16511),
            .in1(N__20207),
            .in2(N__15473),
            .in3(N__23686),
            .lcout(ScreenBuffer_0_11Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19974),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_12_RNO_0_0_LC_6_12_2.C_ON=1'b0;
    defparam ScreenBuffer_0_12_RNO_0_0_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_12_RNO_0_0_LC_6_12_2.LUT_INIT=16'b0000001000000000;
    LogicCell40 ScreenBuffer_0_12_RNO_0_0_LC_6_12_2 (
            .in0(N__16275),
            .in1(N__15981),
            .in2(N__16427),
            .in3(N__19250),
            .lcout(),
            .ltout(un1_sclk17_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_12_0_LC_6_12_3.C_ON=1'b0;
    defparam ScreenBuffer_0_12_0_LC_6_12_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_12_0_LC_6_12_3.LUT_INIT=16'b1101111110000000;
    LogicCell40 ScreenBuffer_0_12_0_LC_6_12_3 (
            .in0(N__16512),
            .in1(N__20208),
            .in2(N__15470),
            .in3(N__18973),
            .lcout(ScreenBuffer_0_12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19974),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATA1_ibuf_RNI800F_LC_6_12_4.C_ON=1'b0;
    defparam SDATA1_ibuf_RNI800F_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam SDATA1_ibuf_RNI800F_LC_6_12_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 SDATA1_ibuf_RNI800F_LC_6_12_4 (
            .in0(N__20206),
            .in1(N__19248),
            .in2(_gnd_net_),
            .in3(N__15978),
            .lcout(ScreenBuffer_0_0_1_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_RNILOQC2_6_LC_6_12_5.C_ON=1'b0;
    defparam slaveselect_RNILOQC2_6_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam slaveselect_RNILOQC2_6_LC_6_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 slaveselect_RNILOQC2_6_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15457),
            .lcout(un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_5_RNO_0_0_LC_6_12_6.C_ON=1'b0;
    defparam ScreenBuffer_0_5_RNO_0_0_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_5_RNO_0_0_LC_6_12_6.LUT_INIT=16'b0001000000000000;
    LogicCell40 ScreenBuffer_0_5_RNO_0_0_LC_6_12_6 (
            .in0(N__16276),
            .in1(N__15979),
            .in2(N__15863),
            .in3(N__19251),
            .lcout(),
            .ltout(un1_sclk17_8_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_5_0_LC_6_12_7.C_ON=1'b0;
    defparam ScreenBuffer_0_5_0_LC_6_12_7.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_5_0_LC_6_12_7.LUT_INIT=16'b1101111110000000;
    LogicCell40 ScreenBuffer_0_5_0_LC_6_12_7 (
            .in0(N__16513),
            .in1(N__20209),
            .in2(N__15446),
            .in3(N__19525),
            .lcout(ScreenBuffer_0_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19974),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_e_0_2_LC_6_13_5.C_ON=1'b0;
    defparam ScreenBuffer_1_3_e_0_2_LC_6_13_5.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_3_e_0_2_LC_6_13_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_3_e_0_2_LC_6_13_5 (
            .in0(N__19334),
            .in1(N__16592),
            .in2(_gnd_net_),
            .in3(N__16559),
            .lcout(ScreenBuffer_1_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19978),
            .ce(N__18430),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_6_RNO_0_0_LC_6_14_0.C_ON=1'b0;
    defparam ScreenBuffer_0_6_RNO_0_0_LC_6_14_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_6_RNO_0_0_LC_6_14_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 ScreenBuffer_0_6_RNO_0_0_LC_6_14_0 (
            .in0(N__16222),
            .in1(N__15994),
            .in2(N__15856),
            .in3(N__19331),
            .lcout(un1_sclk17_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_0_LC_6_14_3.C_ON=1'b0;
    defparam ScreenBuffer_0_7_0_LC_6_14_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_7_0_LC_6_14_3.LUT_INIT=16'b1111100001110000;
    LogicCell40 ScreenBuffer_0_7_0_LC_6_14_3 (
            .in0(N__16499),
            .in1(N__15539),
            .in2(N__19547),
            .in3(N__20162),
            .lcout(ScreenBuffer_0_7Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19981),
            .ce(),
            .sr(_gnd_net_));
    defparam SDATAZ0Z2_LC_6_14_4.C_ON=1'b0;
    defparam SDATAZ0Z2_LC_6_14_4.SEQ_MODE=4'b1000;
    defparam SDATAZ0Z2_LC_6_14_4.LUT_INIT=16'b1010000011001100;
    LogicCell40 SDATAZ0Z2_LC_6_14_4 (
            .in0(N__20161),
            .in1(N__16441),
            .in2(N__16514),
            .in3(N__19332),
            .lcout(SDATA2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19981),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_8_RNO_0_0_LC_6_14_5.C_ON=1'b0;
    defparam ScreenBuffer_0_8_RNO_0_0_LC_6_14_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_8_RNO_0_0_LC_6_14_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 ScreenBuffer_0_8_RNO_0_0_LC_6_14_5 (
            .in0(N__15995),
            .in1(N__15841),
            .in2(N__16425),
            .in3(N__16223),
            .lcout(),
            .ltout(un1_sclk17_9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_8_0_LC_6_14_6.C_ON=1'b0;
    defparam ScreenBuffer_0_8_0_LC_6_14_6.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_8_0_LC_6_14_6.LUT_INIT=16'b1011111110000000;
    LogicCell40 ScreenBuffer_0_8_0_LC_6_14_6 (
            .in0(N__20163),
            .in1(N__20074),
            .in2(N__16430),
            .in3(N__17020),
            .lcout(ScreenBuffer_0_8Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19981),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_9_RNO_0_0_LC_6_14_7.C_ON=1'b0;
    defparam ScreenBuffer_0_9_RNO_0_0_LC_6_14_7.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_9_RNO_0_0_LC_6_14_7.LUT_INIT=16'b0000000010000000;
    LogicCell40 ScreenBuffer_0_9_RNO_0_0_LC_6_14_7 (
            .in0(N__15993),
            .in1(N__15837),
            .in2(N__16424),
            .in3(N__16221),
            .lcout(un1_sclk17_5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNO_0_0_LC_6_15_4.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNO_0_0_LC_6_15_4.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNO_0_0_LC_6_15_4.LUT_INIT=16'b0000010000000000;
    LogicCell40 ScreenBuffer_0_7_RNO_0_0_LC_6_15_4 (
            .in0(N__16266),
            .in1(N__15996),
            .in2(N__15857),
            .in3(N__19333),
            .lcout(un1_sclk17_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_0_LC_7_1_5.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_0_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_0_LC_7_1_5.LUT_INIT=16'b0011001100110011;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_0_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(N__19715),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_7_2_0.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_7_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_7_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(N__22731),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3V_LC_7_2_1.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3V_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3V_LC_7_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3V_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(N__16673),
            .in2(N__16601),
            .in3(N__16658),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKID91_LC_7_2_2.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKID91_LC_7_2_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKID91_LC_7_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKID91_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(N__19718),
            .in2(N__19775),
            .in3(N__16646),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIU1G53_LC_7_2_3.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIU1G53_LC_7_2_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIU1G53_LC_7_2_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIU1G53_LC_7_2_3 (
            .in0(N__16631),
            .in1(N__16616),
            .in2(N__19757),
            .in3(N__16637),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_LC_7_2_4.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_LC_7_2_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_LC_7_2_4 (
            .in0(_gnd_net_),
            .in1(N__19736),
            .in2(_gnd_net_),
            .in3(N__16634),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30T_LC_7_2_5.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30T_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30T_LC_7_2_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30T_LC_7_2_5 (
            .in0(N__19756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19717),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_7_2_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_7_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22732),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_7_2_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_7_2_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_7_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_7_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22253),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_7_3_0.C_ON=1'b0;
    defparam beamX_1_LC_7_3_0.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_7_3_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__17900),
            .in2(_gnd_net_),
            .in3(N__18699),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21060),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_7_4_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__22305),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_7_4_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_7_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__18299),
            .in2(_gnd_net_),
            .in3(N__16694),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_7_4_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__16682),
            .in2(N__21851),
            .in3(N__16691),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_7_4_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_7_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__22004),
            .in2(_gnd_net_),
            .in3(N__16688),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_7_4_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_7_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16685),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_4_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_7_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_7_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22003),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__ANC4_0_i_LC_7_4_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__ANC4_0_i_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__ANC4_0_i_LC_7_4_6.LUT_INIT=16'b1111111101010101;
    LogicCell40 un113_pixel_4_0_15__ANC4_0_i_LC_7_4_6 (
            .in0(N__22005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22140),
            .lcout(N_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__N_32_i_LC_7_5_0.C_ON=1'b1;
    defparam un113_pixel_4_0_15__N_32_i_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__N_32_i_LC_7_5_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un113_pixel_4_0_15__N_32_i_LC_7_5_0 (
            .in0(_gnd_net_),
            .in1(N__22255),
            .in2(_gnd_net_),
            .in3(N__22309),
            .lcout(N_32_i),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_5_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(N__16748),
            .in2(N__19792),
            .in3(N__16676),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_5_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_5_2 (
            .in0(_gnd_net_),
            .in1(N__16738),
            .in2(N__16784),
            .in3(N__16775),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_7_5_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_7_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_7_5_3 (
            .in0(N__16834),
            .in1(N__16724),
            .in2(N__16772),
            .in3(N__16763),
            .lcout(charx_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_7_5_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_7_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_7_5_4 (
            .in0(N__16739),
            .in1(N__22020),
            .in2(N__16760),
            .in3(N__16751),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_7_5_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_7_5_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_7_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16747),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5),
            .ltout(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_5_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16727),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un26_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_5_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_5_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_5_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_7_5_7 (
            .in0(N__22256),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(N__22743),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_7_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_7_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__16816),
            .in2(N__16718),
            .in3(N__16709),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_7_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_7_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(N__16835),
            .in2(N__16706),
            .in3(N__16697),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_7_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_7_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_7_6_3 (
            .in0(N__22776),
            .in1(N__16817),
            .in2(N__16862),
            .in3(N__16853),
            .lcout(charx_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_7_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_7_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_7_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_7_6_4 (
            .in0(_gnd_net_),
            .in1(N__16850),
            .in2(_gnd_net_),
            .in3(N__16844),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un18_beamylto9_2_LC_7_6_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un18_beamylto9_2_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un18_beamylto9_2_LC_7_6_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 un113_pixel_4_0_15__un18_beamylto9_2_LC_7_6_6 (
            .in0(N__18367),
            .in1(N__17680),
            .in2(N__17620),
            .in3(N__18334),
            .lcout(un113_pixel_4_0_15__un18_beamylto9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_7_6_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_7_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_7_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16833),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_0_LC_7_7_1.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_0_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_0_LC_7_7_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_0_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__17069),
            .in2(_gnd_net_),
            .in3(N__17120),
            .lcout(g1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un3_beamx_2_LC_7_7_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un3_beamx_2_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un3_beamx_2_LC_7_7_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 un113_pixel_4_0_15__un3_beamx_2_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__18335),
            .in2(_gnd_net_),
            .in3(N__18368),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_LC_7_8_0.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_LC_7_8_0.LUT_INIT=16'b1000101001110101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_LC_7_8_0 (
            .in0(N__18614),
            .in1(N__24349),
            .in2(N__18406),
            .in3(N__18381),
            .lcout(charx_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI80GJR1_LC_7_8_1.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI80GJR1_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI80GJR1_LC_7_8_1.LUT_INIT=16'b1010101001010101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI80GJR1_LC_7_8_1 (
            .in0(N__24354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18617),
            .lcout(charx_if_generate_plus_mult1_un1_sum_axb1),
            .ltout(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_LC_7_8_2.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_LC_7_8_2.LUT_INIT=16'b1111000000001111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16787),
            .in3(N__17119),
            .lcout(font_un3_pixel_28),
            .ltout(font_un3_pixel_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un61_pixel_LC_7_8_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un61_pixel_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un61_pixel_LC_7_8_3.LUT_INIT=16'b0000000000000010;
    LogicCell40 un113_pixel_4_0_15__font_un61_pixel_LC_7_8_3 (
            .in0(N__18814),
            .in1(N__21623),
            .in2(N__16940),
            .in3(N__18724),
            .lcout(),
            .ltout(font_un61_pixel_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_1_LC_7_8_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_1_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_1_LC_7_8_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 un113_pixel_4_0_15__font_un125_pixel_m_6_1_LC_7_8_4 (
            .in0(N__16936),
            .in1(N__16925),
            .in2(N__16913),
            .in3(N__16910),
            .lcout(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_0_LC_7_8_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_0_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_0_LC_7_8_5.LUT_INIT=16'b1010011001010101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_0_LC_7_8_5 (
            .in0(N__18382),
            .in1(N__18402),
            .in2(N__24358),
            .in3(N__18615),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_1_LC_7_8_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_1_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_1_LC_7_8_6.LUT_INIT=16'b0111010110001010;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_1_LC_7_8_6 (
            .in0(N__18616),
            .in1(N__24353),
            .in2(N__18407),
            .in3(N__18383),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_LC_7_8_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_LC_7_8_7.LUT_INIT=16'b1001100111001100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_LC_7_8_7 (
            .in0(N__24348),
            .in1(N__18398),
            .in2(_gnd_net_),
            .in3(N__18613),
            .lcout(charx_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIKML437_LC_7_9_0.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIKML437_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIKML437_LC_7_9_0.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIKML437_LC_7_9_0 (
            .in0(N__17065),
            .in1(N__21157),
            .in2(_gnd_net_),
            .in3(N__17113),
            .lcout(font_un3_pixel_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNI5D2AEA_LC_7_9_1.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNI5D2AEA_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNI5D2AEA_LC_7_9_1.LUT_INIT=16'b0110011011000110;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNI5D2AEA_LC_7_9_1 (
            .in0(N__17114),
            .in1(N__16868),
            .in2(N__21163),
            .in3(N__17066),
            .lcout(font_un3_pixel_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9A68G8_0_2_LC_7_9_2.C_ON=1'b0;
    defparam beamY_RNI9A68G8_0_2_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI9A68G8_0_2_LC_7_9_2.LUT_INIT=16'b0010010000011000;
    LogicCell40 beamY_RNI9A68G8_0_2_LC_7_9_2 (
            .in0(N__20934),
            .in1(N__20678),
            .in2(N__20893),
            .in3(N__20981),
            .lcout(font_un28_pixel_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFBK6ED_1_LC_7_9_3.C_ON=1'b0;
    defparam beamY_RNIFBK6ED_1_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIFBK6ED_1_LC_7_9_3.LUT_INIT=16'b1000000000001000;
    LogicCell40 beamY_RNIFBK6ED_1_LC_7_9_3 (
            .in0(N__23285),
            .in1(N__18838),
            .in2(N__20690),
            .in3(N__20882),
            .lcout(font_un67_pixel_ac0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g2_LC_7_9_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g2_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g2_LC_7_9_4.LUT_INIT=16'b1010101001010101;
    LogicCell40 un113_pixel_4_0_15__g2_LC_7_9_4 (
            .in0(N__17068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17116),
            .lcout(un113_pixel_4_0_15__gZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_x2_LC_7_9_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_x2_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_x2_LC_7_9_5.LUT_INIT=16'b1010101001010101;
    LogicCell40 un113_pixel_4_0_15__g0_i_x2_LC_7_9_5 (
            .in0(N__17115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17067),
            .lcout(),
            .ltout(N_9_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_2_LC_7_9_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_2_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_2_LC_7_9_6.LUT_INIT=16'b1111111110111111;
    LogicCell40 un113_pixel_4_0_15__g0_i_2_LC_7_9_6 (
            .in0(N__18725),
            .in1(N__21158),
            .in2(N__17033),
            .in3(N__17030),
            .lcout(un113_pixel_4_0_15__g0_iZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_6_0_LC_7_9_7.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_6_0_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_6_0_LC_7_9_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 un113_pixel_7_1_7__g0_6_0_LC_7_9_7 (
            .in0(N__20982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20935),
            .lcout(un113_pixel_7_1_7__g0_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_8_RNIV2FB2F_0_LC_7_10_0.C_ON=1'b0;
    defparam ScreenBuffer_0_8_RNIV2FB2F_0_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_8_RNIV2FB2F_0_LC_7_10_0.LUT_INIT=16'b0101101001111011;
    LogicCell40 ScreenBuffer_0_8_RNIV2FB2F_0_LC_7_10_0 (
            .in0(N__23510),
            .in1(N__25958),
            .in2(N__23603),
            .in3(N__17024),
            .lcout(),
            .ltout(currentchar_1_9_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_RNIBIJQMK_0_LC_7_10_1.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_RNIBIJQMK_0_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_e_0_RNIBIJQMK_0_LC_7_10_1.LUT_INIT=16'b1000111110000101;
    LogicCell40 ScreenBuffer_1_0_e_0_RNIBIJQMK_0_LC_7_10_1 (
            .in0(N__25960),
            .in1(N__17006),
            .in2(N__16997),
            .in3(N__17164),
            .lcout(ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_9_RNI06IC2F_0_LC_7_10_2.C_ON=1'b0;
    defparam ScreenBuffer_0_9_RNI06IC2F_0_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_9_RNI06IC2F_0_LC_7_10_2.LUT_INIT=16'b0101101001111011;
    LogicCell40 ScreenBuffer_0_9_RNI06IC2F_0_LC_7_10_2 (
            .in0(N__23511),
            .in1(N__25959),
            .in2(N__23604),
            .in3(N__20018),
            .lcout(),
            .ltout(currentchar_1_6_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_RNIEVE0NK_0_LC_7_10_3.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_RNIEVE0NK_0_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_e_0_RNIEVE0NK_0_LC_7_10_3.LUT_INIT=16'b1000111110000101;
    LogicCell40 ScreenBuffer_1_1_e_0_RNIEVE0NK_0_LC_7_10_3 (
            .in0(N__25961),
            .in1(N__16994),
            .in2(N__16982),
            .in3(N__16978),
            .lcout(ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_RNISJ0D2F_4_LC_7_10_4.C_ON=1'b0;
    defparam ScreenBuffer_1_0_RNISJ0D2F_4_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_RNISJ0D2F_4_LC_7_10_4.LUT_INIT=16'b1110110110100101;
    LogicCell40 ScreenBuffer_1_0_RNISJ0D2F_4_LC_7_10_4 (
            .in0(N__23512),
            .in1(N__25962),
            .in2(N__23605),
            .in3(N__16958),
            .lcout(),
            .ltout(ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_RNIQ3KT7J1_4_LC_7_10_5.C_ON=1'b0;
    defparam ScreenBuffer_1_0_RNIQ3KT7J1_4_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_RNIQ3KT7J1_4_LC_7_10_5.LUT_INIT=16'b1101100101010001;
    LogicCell40 ScreenBuffer_1_0_RNIQ3KT7J1_4_LC_7_10_5 (
            .in0(N__17132),
            .in1(N__25539),
            .in2(N__17285),
            .in3(N__17126),
            .lcout(),
            .ltout(ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_RNIVUON9Q2_4_LC_7_10_6.C_ON=1'b0;
    defparam ScreenBuffer_1_0_RNIVUON9Q2_4_LC_7_10_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_RNIVUON9Q2_4_LC_7_10_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 ScreenBuffer_1_0_RNIVUON9Q2_4_LC_7_10_6 (
            .in0(_gnd_net_),
            .in1(N__22984),
            .in2(N__17282),
            .in3(N__25396),
            .lcout(currentchar_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_LC_7_11_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_LC_7_11_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_LC_7_11_0 (
            .in0(N__17237),
            .in1(N__17279),
            .in2(N__17264),
            .in3(N__23513),
            .lcout(un3_rowlto0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_7_11_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_7_11_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_7_11_1 (
            .in0(N__17278),
            .in1(N__17260),
            .in2(_gnd_net_),
            .in3(N__17236),
            .lcout(un3_rowlto1),
            .ltout(un3_rowlto1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_e_0_RNINV7VE9_0_LC_7_11_2.C_ON=1'b0;
    defparam ScreenBuffer_1_2_e_0_RNINV7VE9_0_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_2_e_0_RNINV7VE9_0_LC_7_11_2.LUT_INIT=16'b1110110101001000;
    LogicCell40 ScreenBuffer_1_2_e_0_RNINV7VE9_0_LC_7_11_2 (
            .in0(N__23502),
            .in1(N__17219),
            .in2(N__17213),
            .in3(N__17206),
            .lcout(ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_0_0_LC_7_11_3.C_ON=1'b0;
    defparam ScreenBuffer_0_0_0_LC_7_11_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_0_0_LC_7_11_3.LUT_INIT=16'b1111100001110000;
    LogicCell40 ScreenBuffer_0_0_0_LC_7_11_3 (
            .in0(N__19326),
            .in1(N__17189),
            .in2(N__17168),
            .in3(N__20210),
            .lcout(ScreenBuffer_0_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19975),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_RNITM3E2F_4_LC_7_11_4.C_ON=1'b0;
    defparam ScreenBuffer_1_1_RNITM3E2F_4_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_RNITM3E2F_4_LC_7_11_4.LUT_INIT=16'b1110110110100101;
    LogicCell40 ScreenBuffer_1_1_RNITM3E2F_4_LC_7_11_4 (
            .in0(N__23503),
            .in1(N__25985),
            .in2(N__23607),
            .in3(N__17153),
            .lcout(),
            .ltout(ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_RNI4PNO0E3_4_LC_7_11_5.C_ON=1'b0;
    defparam ScreenBuffer_1_1_RNI4PNO0E3_4_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_RNI4PNO0E3_4_LC_7_11_5.LUT_INIT=16'b0000010110111011;
    LogicCell40 ScreenBuffer_1_1_RNI4PNO0E3_4_LC_7_11_5 (
            .in0(N__25545),
            .in1(N__17315),
            .in2(N__17135),
            .in3(N__25740),
            .lcout(currentchar_1_11_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_RNIUP6F2F_4_LC_7_11_6.C_ON=1'b0;
    defparam ScreenBuffer_1_2_RNIUP6F2F_4_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_2_RNIUP6F2F_4_LC_7_11_6.LUT_INIT=16'b1110110110100101;
    LogicCell40 ScreenBuffer_1_2_RNIUP6F2F_4_LC_7_11_6 (
            .in0(N__23504),
            .in1(N__25986),
            .in2(N__23608),
            .in3(N__17390),
            .lcout(ScreenBuffer_1_2_RNIUP6F2FZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_0_1_LC_7_11_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_0_1_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_0_1_LC_7_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 un113_pixel_4_0_15__g0_0_1_LC_7_11_7 (
            .in0(N__24130),
            .in1(N__17300),
            .in2(_gnd_net_),
            .in3(N__17291),
            .lcout(N_4566_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_RNIVS9G2F_4_LC_7_12_0.C_ON=1'b0;
    defparam ScreenBuffer_1_3_RNIVS9G2F_4_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_3_RNIVS9G2F_4_LC_7_12_0.LUT_INIT=16'b1110110110100101;
    LogicCell40 ScreenBuffer_1_3_RNIVS9G2F_4_LC_7_12_0 (
            .in0(N__23527),
            .in1(N__25984),
            .in2(N__23606),
            .in3(N__17333),
            .lcout(ScreenBuffer_1_3_RNIVS9G2FZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam g1_1_LC_7_12_1.C_ON=1'b0;
    defparam g1_1_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam g1_1_LC_7_12_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 g1_1_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(N__23585),
            .in2(_gnd_net_),
            .in3(N__23528),
            .lcout(),
            .ltout(g1Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_22_LC_7_12_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_22_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_22_LC_7_12_2.LUT_INIT=16'b1110000000100000;
    LogicCell40 un113_pixel_4_0_15__g0_22_LC_7_12_2 (
            .in0(N__19385),
            .in1(N__25546),
            .in2(N__17309),
            .in3(N__19379),
            .lcout(),
            .ltout(N_1428_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g1_1_0_LC_7_12_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g1_1_0_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g1_1_0_LC_7_12_3.LUT_INIT=16'b0000000001001100;
    LogicCell40 un113_pixel_4_0_15__g1_1_0_LC_7_12_3 (
            .in0(N__25395),
            .in1(N__23870),
            .in2(N__17306),
            .in3(N__23972),
            .lcout(),
            .ltout(un113_pixel_4_0_15__g1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_21_LC_7_12_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_21_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_21_LC_7_12_4.LUT_INIT=16'b1010100011101100;
    LogicCell40 un113_pixel_4_0_15__g0_21_LC_7_12_4 (
            .in0(N__24514),
            .in1(N__24777),
            .in2(N__17303),
            .in3(N__17339),
            .lcout(N_1300_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_24_LC_7_12_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_24_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_24_LC_7_12_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 un113_pixel_4_0_15__g0_24_LC_7_12_5 (
            .in0(N__25136),
            .in1(N__25028),
            .in2(_gnd_net_),
            .in3(N__24513),
            .lcout(),
            .ltout(un112_pixel_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_1_2_LC_7_12_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_1_2_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_1_2_LC_7_12_6.LUT_INIT=16'b0001110100001100;
    LogicCell40 un113_pixel_4_0_15__g0_1_2_LC_7_12_6 (
            .in0(N__25029),
            .in1(N__24776),
            .in2(N__17294),
            .in3(N__25211),
            .lcout(N_1293_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m10_0_x1_LC_7_13_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m10_0_x1_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m10_0_x1_LC_7_13_0.LUT_INIT=16'b0000011100000000;
    LogicCell40 un113_pixel_4_0_15__m10_0_x1_LC_7_13_0 (
            .in0(N__25991),
            .in1(N__25405),
            .in2(N__23030),
            .in3(N__21526),
            .lcout(m10_0_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_2_4_LC_7_13_1.C_ON=1'b0;
    defparam ScreenBuffer_1_2_4_LC_7_13_1.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_2_4_LC_7_13_1.LUT_INIT=16'b1101110100010001;
    LogicCell40 ScreenBuffer_1_2_4_LC_7_13_1 (
            .in0(N__19318),
            .in1(N__17399),
            .in2(_gnd_net_),
            .in3(N__17389),
            .lcout(ScreenBuffer_1_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19982),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_1_2_2_LC_7_13_2.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_1_2_2_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_1_2_2_LC_7_13_2.LUT_INIT=16'b1111111001011110;
    LogicCell40 un113_pixel_3_0_11__currentchar_1_2_2_LC_7_13_2 (
            .in0(N__25738),
            .in1(N__17375),
            .in2(N__25538),
            .in3(N__17369),
            .lcout(),
            .ltout(un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_1_4_2_LC_7_13_3.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_1_4_2_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_1_4_2_LC_7_13_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 un113_pixel_3_0_11__currentchar_1_4_2_LC_7_13_3 (
            .in0(N__25403),
            .in1(N__25989),
            .in2(N__17354),
            .in3(N__22874),
            .lcout(un113_pixel_3_0_11__currentchar_1_4Z0Z_2),
            .ltout(un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un112_pixel_1_2_x1_LC_7_13_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un112_pixel_1_2_x1_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un112_pixel_1_2_x1_LC_7_13_4.LUT_INIT=16'b1100110111001111;
    LogicCell40 un113_pixel_4_0_15__un112_pixel_1_2_x1_LC_7_13_4 (
            .in0(N__25990),
            .in1(N__22994),
            .in2(N__17351),
            .in3(N__25404),
            .lcout(un112_pixel_1_2_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m10_0_ns_LC_7_13_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m10_0_ns_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m10_0_ns_LC_7_13_5.LUT_INIT=16'b1100110000001010;
    LogicCell40 un113_pixel_4_0_15__m10_0_ns_LC_7_13_5 (
            .in0(N__21527),
            .in1(N__17348),
            .in2(N__23018),
            .in3(N__19511),
            .lcout(un112_pixel_2_2),
            .ltout(un112_pixel_2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_LC_7_13_6.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_LC_7_13_6.LUT_INIT=16'b0010001010111000;
    LogicCell40 ScreenBuffer_0_7_RNIHMH43T2_0_LC_7_13_6 (
            .in0(N__23433),
            .in1(N__25007),
            .in2(N__17342),
            .in3(N__24504),
            .lcout(ScreenBuffer_0_7_RNIHMH43T2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_0_0_LC_7_13_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_0_0_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_0_0_LC_7_13_7.LUT_INIT=16'b1101001000000000;
    LogicCell40 un113_pixel_3_0_11__g0_0_0_LC_7_13_7 (
            .in0(N__21528),
            .in1(N__23015),
            .in2(N__25068),
            .in3(N__23886),
            .lcout(un113_pixel_3_0_11__g0_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_4_am_7_LC_7_14_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_4_am_7_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_4_am_7_LC_7_14_0.LUT_INIT=16'b0010001010001000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_4_am_7_LC_7_14_0 (
            .in0(N__23421),
            .in1(N__25017),
            .in2(_gnd_net_),
            .in3(N__24476),
            .lcout(un115_pixel_4_am_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDQUNU91_0_LC_7_14_1.C_ON=1'b0;
    defparam beamY_RNIDQUNU91_0_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIDQUNU91_0_LC_7_14_1.LUT_INIT=16'b0010111100001111;
    LogicCell40 beamY_RNIDQUNU91_0_LC_7_14_1 (
            .in0(N__24477),
            .in1(N__25026),
            .in2(N__24860),
            .in3(N__23424),
            .lcout(),
            .ltout(beamY_RNIDQUNU91Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7RM4IF_0_LC_7_14_2.C_ON=1'b0;
    defparam beamY_RNI7RM4IF_0_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI7RM4IF_0_LC_7_14_2.LUT_INIT=16'b1010101011110000;
    LogicCell40 beamY_RNI7RM4IF_0_LC_7_14_2 (
            .in0(N__17429),
            .in1(_gnd_net_),
            .in2(N__17423),
            .in3(N__24138),
            .lcout(beamY_RNI7RM4IFZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC0GLNQ_0_LC_7_14_3.C_ON=1'b0;
    defparam beamY_RNIC0GLNQ_0_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIC0GLNQ_0_LC_7_14_3.LUT_INIT=16'b1100101011000000;
    LogicCell40 beamY_RNIC0GLNQ_0_LC_7_14_3 (
            .in0(N__25016),
            .in1(N__23423),
            .in2(N__24861),
            .in3(N__25133),
            .lcout(),
            .ltout(un115_pixel_2_sn_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPQEDM42_0_LC_7_14_4.C_ON=1'b0;
    defparam beamY_RNIPQEDM42_0_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIPQEDM42_0_LC_7_14_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 beamY_RNIPQEDM42_0_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(N__17414),
            .in2(N__17420),
            .in3(N__24479),
            .lcout(beamY_RNIPQEDM42Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un112_pixel_7_LC_7_14_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un112_pixel_7_LC_7_14_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un112_pixel_7_LC_7_14_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 un113_pixel_4_0_15__un112_pixel_7_LC_7_14_5 (
            .in0(N__24478),
            .in1(N__25027),
            .in2(_gnd_net_),
            .in3(N__25134),
            .lcout(),
            .ltout(un112_pixel_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_1_4_LC_7_14_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_1_4_LC_7_14_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_1_4_LC_7_14_6.LUT_INIT=16'b0001101100001010;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_1_4_LC_7_14_6 (
            .in0(N__24760),
            .in1(N__25018),
            .in2(N__17417),
            .in3(N__25207),
            .lcout(N_1293),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIINK7J73_0_LC_7_14_7.C_ON=1'b0;
    defparam beamY_RNIINK7J73_0_LC_7_14_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIINK7J73_0_LC_7_14_7.LUT_INIT=16'b0001000111001100;
    LogicCell40 beamY_RNIINK7J73_0_LC_7_14_7 (
            .in0(N__25015),
            .in1(N__24759),
            .in2(_gnd_net_),
            .in3(N__23422),
            .lcout(beamY_RNIINK7J73Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_8_1_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_8_1_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_8_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_8_1_0 (
            .in0(_gnd_net_),
            .in1(N__17903),
            .in2(N__18742),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_8_1_1.C_ON=1'b1;
    defparam beamX_2_LC_8_1_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_8_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_8_1_1 (
            .in0(_gnd_net_),
            .in1(N__17859),
            .in2(_gnd_net_),
            .in3(N__17408),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_8_1_2.C_ON=1'b1;
    defparam beamX_3_LC_8_1_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_8_1_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_8_1_2 (
            .in0(_gnd_net_),
            .in1(N__17828),
            .in2(_gnd_net_),
            .in3(N__17405),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_8_1_3.C_ON=1'b1;
    defparam beamX_4_LC_8_1_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_8_1_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_8_1_3 (
            .in0(N__17545),
            .in1(N__17762),
            .in2(_gnd_net_),
            .in3(N__17402),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_8_1_4.C_ON=1'b1;
    defparam beamX_5_LC_8_1_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_8_1_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_8_1_4 (
            .in0(_gnd_net_),
            .in1(N__17712),
            .in2(_gnd_net_),
            .in3(N__17561),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_8_1_5.C_ON=1'b1;
    defparam beamX_6_LC_8_1_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_8_1_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_8_1_5 (
            .in0(_gnd_net_),
            .in1(N__17661),
            .in2(_gnd_net_),
            .in3(N__17558),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_8_1_6.C_ON=1'b1;
    defparam beamX_7_LC_8_1_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_8_1_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_8_1_6 (
            .in0(_gnd_net_),
            .in1(N__17596),
            .in2(_gnd_net_),
            .in3(N__17555),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_8_1_7.C_ON=1'b1;
    defparam beamX_8_LC_8_1_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_8_1_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_8_1_7 (
            .in0(_gnd_net_),
            .in1(N__18359),
            .in2(_gnd_net_),
            .in3(N__17552),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__21062),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_8_2_0.C_ON=1'b1;
    defparam beamX_9_LC_8_2_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_8_2_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_8_2_0 (
            .in0(_gnd_net_),
            .in1(N__18326),
            .in2(_gnd_net_),
            .in3(N__17549),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__21061),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_8_2_1.C_ON=1'b0;
    defparam beamX_10_LC_8_2_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_8_2_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_8_2_1 (
            .in0(N__17462),
            .in1(N__17540),
            .in2(_gnd_net_),
            .in3(N__17471),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21061),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_2_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_2_2.LUT_INIT=16'b0101010111111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_2_2 (
            .in0(N__22141),
            .in1(N__22254),
            .in2(_gnd_net_),
            .in3(N__22072),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_2_3.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_2_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_2_3 (
            .in0(N__22074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22143),
            .lcout(if_generate_plus_mult1_un47_sum_0_cry_3_ma),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__N_1184_0_i_LC_8_2_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__N_1184_0_i_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__N_1184_0_i_LC_8_2_4.LUT_INIT=16'b0011001111111111;
    LogicCell40 un113_pixel_4_0_15__N_1184_0_i_LC_8_2_4 (
            .in0(_gnd_net_),
            .in1(N__22147),
            .in2(_gnd_net_),
            .in3(N__22075),
            .lcout(N_1184_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_2_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_2_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_2_7.LUT_INIT=16'b1101011111011000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_2_7 (
            .in0(N__22073),
            .in1(N__22142),
            .in2(N__22157),
            .in3(N__22188),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_8_3_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__18700),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_8_3_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_8_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(N__17891),
            .in2(_gnd_net_),
            .in3(N__17870),
            .lcout(charx_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_8_3_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_8_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(N__17860),
            .in2(_gnd_net_),
            .in3(N__17837),
            .lcout(charx_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_8_3_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_8_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_8_3_3 (
            .in0(_gnd_net_),
            .in1(N__17819),
            .in2(N__21870),
            .in3(N__17795),
            .lcout(chessboardpixel_un151_pixel_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_3_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_8_3_4 (
            .in0(_gnd_net_),
            .in1(N__17763),
            .in2(_gnd_net_),
            .in3(N__17732),
            .lcout(charx_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_3_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(N__17713),
            .in2(_gnd_net_),
            .in3(N__17690),
            .lcout(charx_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_3_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_3_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(N__21844),
            .in2(N__17679),
            .in3(N__17624),
            .lcout(charx_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_3_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_8_3_7 (
            .in0(_gnd_net_),
            .in1(N__17597),
            .in2(_gnd_net_),
            .in3(N__17564),
            .lcout(charx_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_4_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_4_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__18360),
            .in2(N__21900),
            .in3(N__18338),
            .lcout(un5_visiblex_cry_7_c_RNIVZ0Z952),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_4_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_4_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__18327),
            .in2(_gnd_net_),
            .in3(N__18305),
            .lcout(CO3_0),
            .ltout(CO3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_4_2.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_4_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18302),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un26_sum_s_2_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un4_row_1_LC_8_4_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un4_row_1_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un4_row_1_LC_8_4_3.LUT_INIT=16'b0111000000000000;
    LogicCell40 un113_pixel_4_0_15__un4_row_1_LC_8_4_3 (
            .in0(N__18293),
            .in1(N__18170),
            .in2(N__18050),
            .in3(N__20348),
            .lcout(un113_pixel_4_0_15__un4_rowZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_4_4.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_4_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_8_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22310),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam voltage_0_0_LC_8_5_0.C_ON=1'b0;
    defparam voltage_0_0_LC_8_5_0.SEQ_MODE=4'b1000;
    defparam voltage_0_0_LC_8_5_0.LUT_INIT=16'b0011001110111011;
    LogicCell40 voltage_0_0_LC_8_5_0 (
            .in0(N__18026),
            .in1(N__18008),
            .in2(_gnd_net_),
            .in3(N__17990),
            .lcout(voltage_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19980),
            .ce(),
            .sr(N__18548));
    defparam voltage_0_1_LC_8_5_1.C_ON=1'b0;
    defparam voltage_0_1_LC_8_5_1.SEQ_MODE=4'b1000;
    defparam voltage_0_1_LC_8_5_1.LUT_INIT=16'b0111011100110011;
    LogicCell40 voltage_0_1_LC_8_5_1 (
            .in0(N__17989),
            .in1(N__17957),
            .in2(_gnd_net_),
            .in3(N__17945),
            .lcout(voltage_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19980),
            .ce(),
            .sr(N__18548));
    defparam nCS1_1_LC_8_5_2.C_ON=1'b0;
    defparam nCS1_1_LC_8_5_2.SEQ_MODE=4'b1001;
    defparam nCS1_1_LC_8_5_2.LUT_INIT=16'b1101110100010001;
    LogicCell40 nCS1_1_LC_8_5_2 (
            .in0(N__18578),
            .in1(N__19113),
            .in2(_gnd_net_),
            .in3(N__17914),
            .lcout(nCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19980),
            .ce(),
            .sr(N__18548));
    defparam slaveselect_LC_8_5_3.C_ON=1'b0;
    defparam slaveselect_LC_8_5_3.SEQ_MODE=4'b1000;
    defparam slaveselect_LC_8_5_3.LUT_INIT=16'b1110111011101110;
    LogicCell40 slaveselect_LC_8_5_3 (
            .in0(N__19114),
            .in1(N__18577),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(slaveselectZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19980),
            .ce(),
            .sr(N__18548));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_8_5_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_8_5_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_8_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22817),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_e_0_0_LC_8_6_0.C_ON=1'b0;
    defparam ScreenBuffer_1_3_e_0_0_LC_8_6_0.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_3_e_0_0_LC_8_6_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_3_e_0_0_LC_8_6_0 (
            .in0(N__19110),
            .in1(N__18518),
            .in2(_gnd_net_),
            .in3(N__18456),
            .lcout(ScreenBuffer_1_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19976),
            .ce(N__18434),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_e_0_3_LC_8_6_2.C_ON=1'b0;
    defparam ScreenBuffer_1_3_e_0_3_LC_8_6_2.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_3_e_0_3_LC_8_6_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_3_e_0_3_LC_8_6_2 (
            .in0(N__19111),
            .in1(N__19463),
            .in2(_gnd_net_),
            .in3(N__19433),
            .lcout(ScreenBuffer_1_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19976),
            .ce(N__18434),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_e_0_1_LC_8_6_3.C_ON=1'b0;
    defparam ScreenBuffer_1_3_e_0_1_LC_8_6_3.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_3_e_0_1_LC_8_6_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 ScreenBuffer_1_3_e_0_1_LC_8_6_3 (
            .in0(N__19030),
            .in1(N__19373),
            .in2(_gnd_net_),
            .in3(N__19112),
            .lcout(ScreenBuffer_1_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19976),
            .ce(N__18434),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_8_6_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_8_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22769),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_7_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_8_7_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_8_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(N__18628),
            .in2(N__18599),
            .in3(N__18386),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPME1_LC_8_7_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPME1_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPME1_LC_8_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPME1_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__20381),
            .in2(N__20441),
            .in3(N__18371),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_7_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(N__18629),
            .in2(N__20420),
            .in3(N__20379),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHR1_LC_8_7_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHR1_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHR1_LC_8_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHR1_LC_8_7_4 (
            .in0(_gnd_net_),
            .in1(N__20399),
            .in2(_gnd_net_),
            .in3(N__18620),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_7_5.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22665),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_8_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(N__23080),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_8_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__20473),
            .in2(N__18851),
            .in3(N__18590),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_8_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_8_2 (
            .in0(_gnd_net_),
            .in1(N__25871),
            .in2(N__20588),
            .in3(N__18587),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_8_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_8_3 (
            .in0(N__25310),
            .in1(N__20474),
            .in2(N__20537),
            .in3(N__18584),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_8_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_8_4 (
            .in0(_gnd_net_),
            .in1(N__20495),
            .in2(_gnd_net_),
            .in3(N__18581),
            .lcout(column_1_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9A68G8_2_LC_8_8_6.C_ON=1'b0;
    defparam beamY_RNI9A68G8_2_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI9A68G8_2_LC_8_8_6.LUT_INIT=16'b0110100101100110;
    LogicCell40 beamY_RNI9A68G8_2_LC_8_8_6 (
            .in0(N__20983),
            .in1(N__20933),
            .in2(N__20894),
            .in3(N__20672),
            .lcout(chary_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_8_8_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_8_8_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_8_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_i_LC_8_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22619),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFBK6ED_0_1_LC_8_9_0.C_ON=1'b0;
    defparam beamY_RNIFBK6ED_0_1_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIFBK6ED_0_1_LC_8_9_0.LUT_INIT=16'b0001001000100001;
    LogicCell40 beamY_RNIFBK6ED_0_1_LC_8_9_0 (
            .in0(N__20689),
            .in1(N__23300),
            .in2(N__18842),
            .in3(N__20892),
            .lcout(font_un64_pixel_ac0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_0_2_LC_8_9_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_0_2_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_0_2_LC_8_9_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 un113_pixel_4_0_15__g0_0_2_LC_8_9_1 (
            .in0(N__21625),
            .in1(N__18740),
            .in2(N__18827),
            .in3(N__18637),
            .lcout(un113_pixel_4_0_15__g0_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un57_pixel_LC_8_9_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un57_pixel_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un57_pixel_LC_8_9_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 un113_pixel_4_0_15__font_un57_pixel_LC_8_9_2 (
            .in0(N__18815),
            .in1(N__21624),
            .in2(N__18743),
            .in3(N__21289),
            .lcout(),
            .ltout(font_un57_pixel_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_3_LC_8_9_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_3_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_3_LC_8_9_3.LUT_INIT=16'b0000110000000000;
    LogicCell40 un113_pixel_4_0_15__font_un125_pixel_m_6_3_LC_8_9_3 (
            .in0(_gnd_net_),
            .in1(N__18803),
            .in2(N__18797),
            .in3(N__18794),
            .lcout(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3),
            .ltout(un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_LC_8_9_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un125_pixel_m_6_LC_8_9_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 un113_pixel_4_0_15__font_un125_pixel_m_6_LC_8_9_4 (
            .in0(N__18788),
            .in1(N__18779),
            .in2(N__18773),
            .in3(N__21258),
            .lcout(un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_5_LC_8_9_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_5_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_5_LC_8_9_5.LUT_INIT=16'b1111111011111111;
    LogicCell40 un113_pixel_4_0_15__g0_i_5_LC_8_9_5 (
            .in0(N__21259),
            .in1(N__18770),
            .in2(N__18758),
            .in3(N__21235),
            .lcout(),
            .ltout(un113_pixel_4_0_15__g0_iZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_1_1_LC_8_9_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_1_1_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_1_1_LC_8_9_6.LUT_INIT=16'b0000111000000100;
    LogicCell40 un113_pixel_4_0_15__g0_1_1_LC_8_9_6 (
            .in0(N__23348),
            .in1(N__18905),
            .in2(N__18746),
            .in3(N__21587),
            .lcout(g0_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__Pixel_6_iv_a3_0_LC_8_9_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__Pixel_6_iv_a3_0_LC_8_9_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__Pixel_6_iv_a3_0_LC_8_9_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 un113_pixel_4_0_15__Pixel_6_iv_a3_0_LC_8_9_7 (
            .in0(_gnd_net_),
            .in1(N__18741),
            .in2(_gnd_net_),
            .in3(N__18638),
            .lcout(un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un112_pixel_7_1_LC_8_10_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un112_pixel_7_1_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un112_pixel_7_1_LC_8_10_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 un113_pixel_4_0_15__un112_pixel_7_1_LC_8_10_0 (
            .in0(N__21325),
            .in1(N__25360),
            .in2(_gnd_net_),
            .in3(N__25585),
            .lcout(un112_pixel_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIOEPPEK1_0_LC_8_10_1.C_ON=1'b0;
    defparam beamY_RNIOEPPEK1_0_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIOEPPEK1_0_LC_8_10_1.LUT_INIT=16'b0000101000000000;
    LogicCell40 beamY_RNIOEPPEK1_0_LC_8_10_1 (
            .in0(N__25364),
            .in1(_gnd_net_),
            .in2(N__24852),
            .in3(N__21324),
            .lcout(),
            .ltout(beamY_RNIOEPPEK1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1G38U63_0_LC_8_10_2.C_ON=1'b0;
    defparam beamY_RNI1G38U63_0_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI1G38U63_0_LC_8_10_2.LUT_INIT=16'b0111110111010111;
    LogicCell40 beamY_RNI1G38U63_0_LC_8_10_2 (
            .in0(N__23879),
            .in1(N__23998),
            .in2(N__18920),
            .in3(N__24542),
            .lcout(),
            .ltout(N_3461_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_19_LC_8_10_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_19_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_19_LC_8_10_3.LUT_INIT=16'b0111001001010000;
    LogicCell40 un113_pixel_4_0_15__g0_19_LC_8_10_3 (
            .in0(N__24800),
            .in1(N__18917),
            .in2(N__18911),
            .in3(N__23443),
            .lcout(),
            .ltout(N_4568_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_18_LC_8_10_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_18_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_18_LC_8_10_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 un113_pixel_4_0_15__g0_18_LC_8_10_4 (
            .in0(N__21443),
            .in1(_gnd_net_),
            .in2(N__18908),
            .in3(N__24168),
            .lcout(N_1305_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_1_LC_8_10_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_1_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_1_LC_8_10_5.LUT_INIT=16'b1010100000001000;
    LogicCell40 un113_pixel_4_0_15__g0_1_LC_8_10_5 (
            .in0(N__18899),
            .in1(N__24242),
            .in2(N__23349),
            .in3(N__19808),
            .lcout(),
            .ltout(N_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_LC_8_10_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_LC_8_10_6.LUT_INIT=16'b0000000100000000;
    LogicCell40 un113_pixel_4_0_15__g0_LC_8_10_6 (
            .in0(N__18893),
            .in1(N__18881),
            .in2(N__18875),
            .in3(N__21206),
            .lcout(un113_pixel_4_0_15__g0_i_a3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un71_pixellto5_1_LC_8_10_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un71_pixellto5_1_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un71_pixellto5_1_LC_8_10_7.LUT_INIT=16'b0000000011101010;
    LogicCell40 un113_pixel_4_0_15__font_un71_pixellto5_1_LC_8_10_7 (
            .in0(N__23999),
            .in1(N__21326),
            .in2(N__25399),
            .in3(N__23880),
            .lcout(font_un71_pixellt7_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_1_LC_8_11_0.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_1_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_1_LC_8_11_0.LUT_INIT=16'b0101000101011011;
    LogicCell40 un113_pixel_3_0_11__currentchar_m7_0_m3_ns_1_LC_8_11_0 (
            .in0(N__25736),
            .in1(N__18872),
            .in2(N__25540),
            .in3(N__18863),
            .lcout(),
            .ltout(un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_LC_8_11_1.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_m7_0_m3_ns_LC_8_11_1.LUT_INIT=16'b1000111110000101;
    LogicCell40 un113_pixel_3_0_11__currentchar_m7_0_m3_ns_LC_8_11_1 (
            .in0(N__25525),
            .in1(N__19478),
            .in2(N__19469),
            .in3(N__19391),
            .lcout(un113_pixel_3_0_11__currentchar_N_13),
            .ltout(un113_pixel_3_0_11__currentchar_N_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_m7_0_1_LC_8_11_2.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_m7_0_1_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_m7_0_1_LC_8_11_2.LUT_INIT=16'b0101111111111111;
    LogicCell40 un113_pixel_3_0_11__currentchar_m7_0_1_LC_8_11_2 (
            .in0(N__25937),
            .in1(_gnd_net_),
            .in2(N__19466),
            .in3(N__25394),
            .lcout(un113_pixel_3_0_11__currentchar_m7_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_3_LC_8_11_4.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_3_LC_8_11_4.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_0_e_0_3_LC_8_11_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 ScreenBuffer_1_0_e_0_3_LC_8_11_4 (
            .in0(N__19462),
            .in1(N__19177),
            .in2(_gnd_net_),
            .in3(N__19432),
            .lcout(ScreenBuffer_1_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19979),
            .ce(N__18998),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_1_0_0_LC_8_11_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_1_0_0_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_1_0_0_LC_8_11_5.LUT_INIT=16'b1110000001000000;
    LogicCell40 un113_pixel_4_0_15__g0_1_0_0_LC_8_11_5 (
            .in0(N__25739),
            .in1(N__21404),
            .in2(N__25988),
            .in3(N__21386),
            .lcout(un113_pixel_4_0_15__g0_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_3_0_0_LC_8_11_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_3_0_0_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_3_0_0_LC_8_11_6.LUT_INIT=16'b1110000001000000;
    LogicCell40 un113_pixel_4_0_15__g0_3_0_0_LC_8_11_6 (
            .in0(N__25737),
            .in1(N__21437),
            .in2(N__25972),
            .in3(N__21422),
            .lcout(un113_pixel_4_0_15__g0_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_1_LC_8_11_7.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_1_LC_8_11_7.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_1_0_e_0_1_LC_8_11_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 ScreenBuffer_1_0_e_0_1_LC_8_11_7 (
            .in0(N__19368),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__19046),
            .lcout(ScreenBuffer_1_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19979),
            .ce(N__18998),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_12_RNIE3Q33F_0_LC_8_12_0.C_ON=1'b0;
    defparam ScreenBuffer_0_12_RNIE3Q33F_0_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_12_RNIE3Q33F_0_LC_8_12_0.LUT_INIT=16'b1110000001000000;
    LogicCell40 ScreenBuffer_0_12_RNIE3Q33F_0_LC_8_12_0 (
            .in0(N__25970),
            .in1(N__18974),
            .in2(N__23016),
            .in3(N__18959),
            .lcout(),
            .ltout(ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_6_RNIVTBDB12_0_LC_8_12_1.C_ON=1'b0;
    defparam ScreenBuffer_0_6_RNIVTBDB12_0_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_6_RNIVTBDB12_0_LC_8_12_1.LUT_INIT=16'b1110010010100000;
    LogicCell40 ScreenBuffer_0_6_RNIVTBDB12_0_LC_8_12_1 (
            .in0(N__25735),
            .in1(N__22990),
            .in2(N__18944),
            .in3(N__18941),
            .lcout(ScreenBuffer_0_6_RNIVTBDB12Z0Z_0),
            .ltout(ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNII0GVLQ_0_LC_8_12_2.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNII0GVLQ_0_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNII0GVLQ_0_LC_8_12_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 ScreenBuffer_0_7_RNII0GVLQ_0_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(N__25541),
            .in2(N__19553),
            .in3(N__25246),
            .lcout(ScreenBuffer_0_7_RNII0GVLQZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_m7_0_LC_8_12_3.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_m7_0_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_m7_0_LC_8_12_3.LUT_INIT=16'b1111011111111111;
    LogicCell40 un113_pixel_3_0_11__currentchar_m7_0_LC_8_12_3 (
            .in0(N__25386),
            .in1(N__25971),
            .in2(N__22986),
            .in3(N__19503),
            .lcout(currentchar_m7_0),
            .ltout(currentchar_m7_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m1_LC_8_12_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m1_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m1_LC_8_12_4.LUT_INIT=16'b1110000001000000;
    LogicCell40 un113_pixel_4_0_15__m1_LC_8_12_4 (
            .in0(N__25387),
            .in1(N__19598),
            .in2(N__19550),
            .in3(N__25586),
            .lcout(un113_pixel_4_0_15__N_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIN5F98I1_0_LC_8_12_5.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIN5F98I1_0_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIN5F98I1_0_LC_8_12_5.LUT_INIT=16'b1110000001000000;
    LogicCell40 ScreenBuffer_0_7_RNIN5F98I1_0_LC_8_12_5 (
            .in0(N__25734),
            .in1(N__19546),
            .in2(N__22985),
            .in3(N__19526),
            .lcout(ScreenBuffer_0_7_RNIN5F98I1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__un115_pixel_5_bm_7_LC_8_12_6.C_ON=1'b0;
    defparam un113_pixel_3_0_11__un115_pixel_5_bm_7_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__un115_pixel_5_bm_7_LC_8_12_6.LUT_INIT=16'b0001000110111011;
    LogicCell40 un113_pixel_3_0_11__un115_pixel_5_bm_7_LC_8_12_6 (
            .in0(N__24484),
            .in1(N__23425),
            .in2(_gnd_net_),
            .in3(N__25141),
            .lcout(un115_pixel_5_bm_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_0_LC_8_12_7.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_0_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIHMH43T2_0_0_LC_8_12_7.LUT_INIT=16'b0100011111011101;
    LogicCell40 ScreenBuffer_0_7_RNIHMH43T2_0_0_LC_8_12_7 (
            .in0(N__25140),
            .in1(N__25006),
            .in2(N__23439),
            .in3(N__24483),
            .lcout(ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_1_12_1_LC_8_13_0.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_1_12_1_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_1_12_1_LC_8_13_0.LUT_INIT=16'b1010100000001000;
    LogicCell40 un113_pixel_3_0_11__currentchar_1_12_1_LC_8_13_0 (
            .in0(N__25406),
            .in1(N__21359),
            .in2(N__25547),
            .in3(N__21341),
            .lcout(currentchar_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un112_pixel_1_2_ns_LC_8_13_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un112_pixel_1_2_ns_LC_8_13_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un112_pixel_1_2_ns_LC_8_13_1.LUT_INIT=16'b1111101101010001;
    LogicCell40 un113_pixel_4_0_15__un112_pixel_1_2_ns_LC_8_13_1 (
            .in0(N__19510),
            .in1(N__21523),
            .in2(N__23031),
            .in3(N__19487),
            .lcout(un112_pixel_2_8),
            .ltout(un112_pixel_2_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__m8_LC_8_13_2.C_ON=1'b0;
    defparam un113_pixel_7_1_7__m8_LC_8_13_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__m8_LC_8_13_2.LUT_INIT=16'b1110000000100000;
    LogicCell40 un113_pixel_7_1_7__m8_LC_8_13_2 (
            .in0(N__19600),
            .in1(N__25417),
            .in2(N__19481),
            .in3(N__25591),
            .lcout(un113_pixel_7_1_7__N_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_1_2_LC_8_13_3.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_1_2_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_1_2_LC_8_13_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 un113_pixel_3_0_11__currentchar_1_2_LC_8_13_3 (
            .in0(_gnd_net_),
            .in1(N__23019),
            .in2(_gnd_net_),
            .in3(N__21524),
            .lcout(currentchar_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_4_ns_7_LC_8_13_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_4_ns_7_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_4_ns_7_LC_8_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_4_ns_7_LC_8_13_4 (
            .in0(N__23322),
            .in1(N__19610),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(),
            .ltout(N_1287_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_7_LC_8_13_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_7_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_7_LC_8_13_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_6_ns_7_LC_8_13_5 (
            .in0(N__24154),
            .in1(_gnd_net_),
            .in2(N__19616),
            .in3(N__21539),
            .lcout(N_1289),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIR2AGB22_0_LC_8_13_6.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIR2AGB22_0_LC_8_13_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIR2AGB22_0_LC_8_13_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 ScreenBuffer_0_7_RNIR2AGB22_0_LC_8_13_6 (
            .in0(N__19599),
            .in1(N__25418),
            .in2(_gnd_net_),
            .in3(N__25590),
            .lcout(currentchar_1_0),
            .ltout(currentchar_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__m10_LC_8_13_7.C_ON=1'b0;
    defparam un113_pixel_7_1_7__m10_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__m10_LC_8_13_7.LUT_INIT=16'b1000001010100000;
    LogicCell40 un113_pixel_7_1_7__m10_LC_8_13_7 (
            .in0(N__23791),
            .in1(N__23020),
            .in2(N__19613),
            .in3(N__21525),
            .lcout(un113_pixel_7_1_7__N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_4_bm_7_LC_8_14_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_4_bm_7_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_4_bm_7_LC_8_14_0.LUT_INIT=16'b1100111111011111;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_4_bm_7_LC_8_14_0 (
            .in0(N__23958),
            .in1(N__25021),
            .in2(N__23881),
            .in3(N__24480),
            .lcout(un115_pixel_4_bm_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__m21_LC_8_14_1.C_ON=1'b0;
    defparam un113_pixel_3_0_11__m21_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__m21_LC_8_14_1.LUT_INIT=16'b1010100000001000;
    LogicCell40 un113_pixel_3_0_11__m21_LC_8_14_1 (
            .in0(N__25135),
            .in1(N__19604),
            .in2(N__25416),
            .in3(N__25592),
            .lcout(un113_pixel_1_0_3__N_10_mux),
            .ltout(un113_pixel_1_0_3__N_10_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_9_LC_8_14_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_9_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_9_LC_8_14_2.LUT_INIT=16'b0111010011111100;
    LogicCell40 un113_pixel_4_0_15__g0_9_LC_8_14_2 (
            .in0(N__23852),
            .in1(N__24153),
            .in2(N__19580),
            .in3(N__19658),
            .lcout(),
            .ltout(N_1285_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_i_m2_0_LC_8_14_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_i_m2_0_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_i_m2_0_LC_8_14_3.LUT_INIT=16'b0111010011010001;
    LogicCell40 un113_pixel_4_0_15__g0_i_m2_0_LC_8_14_3 (
            .in0(N__19559),
            .in1(N__23346),
            .in2(N__19577),
            .in3(N__19574),
            .lcout(N_1286_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__m14_LC_8_14_4.C_ON=1'b0;
    defparam un113_pixel_3_0_11__m14_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__m14_LC_8_14_4.LUT_INIT=16'b1001000001100000;
    LogicCell40 un113_pixel_3_0_11__m14_LC_8_14_4 (
            .in0(N__23959),
            .in1(N__25019),
            .in2(N__23882),
            .in3(N__24481),
            .lcout(m14),
            .ltout(m14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICJUESD2_1_0_LC_8_14_5.C_ON=1'b0;
    defparam beamY_RNICJUESD2_1_0_LC_8_14_5.SEQ_MODE=4'b0000;
    defparam beamY_RNICJUESD2_1_0_LC_8_14_5.LUT_INIT=16'b0001110100001100;
    LogicCell40 beamY_RNICJUESD2_1_0_LC_8_14_5 (
            .in0(N__25020),
            .in1(N__24837),
            .in2(N__19667),
            .in3(N__25205),
            .lcout(beamY_RNICJUESD2_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_4_LC_8_14_6.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_4_LC_8_14_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_4_LC_8_14_6.LUT_INIT=16'b0010111100100000;
    LogicCell40 un113_pixel_7_1_7__g0_4_LC_8_14_6 (
            .in0(N__25206),
            .in1(N__25025),
            .in2(N__21014),
            .in3(N__19664),
            .lcout(N_1327_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g0_6_LC_8_14_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g0_6_LC_8_14_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g0_6_LC_8_14_7.LUT_INIT=16'b0011101100001010;
    LogicCell40 un113_pixel_3_0_11__g0_6_LC_8_14_7 (
            .in0(N__24482),
            .in1(N__23017),
            .in2(N__25069),
            .in3(N__21529),
            .lcout(un113_pixel_3_0_11__g1_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_3_5_LC_8_15_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_3_5_LC_8_15_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_3_5_LC_8_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_3_5_LC_8_15_0 (
            .in0(N__24169),
            .in1(N__19652),
            .in2(_gnd_net_),
            .in3(N__19646),
            .lcout(),
            .ltout(N_1306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_17_LC_8_15_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_17_LC_8_15_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_17_LC_8_15_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_4_0_15__g0_17_LC_8_15_1 (
            .in0(_gnd_net_),
            .in1(N__23347),
            .in2(N__19640),
            .in3(N__19637),
            .lcout(N_4561_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m11_LC_8_15_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m11_LC_8_15_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m11_LC_8_15_2.LUT_INIT=16'b1000100000100010;
    LogicCell40 un113_pixel_4_0_15__m11_LC_8_15_2 (
            .in0(N__25145),
            .in1(N__25065),
            .in2(_gnd_net_),
            .in3(N__24525),
            .lcout(),
            .ltout(m11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_3_LC_8_15_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_3_LC_8_15_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_3_LC_8_15_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_5_ns_3_LC_8_15_3 (
            .in0(_gnd_net_),
            .in1(N__24838),
            .in2(N__19631),
            .in3(N__19628),
            .lcout(N_1322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m16_LC_8_15_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m16_LC_8_15_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m16_LC_8_15_4.LUT_INIT=16'b1000000001000000;
    LogicCell40 un113_pixel_4_0_15__m16_LC_8_15_4 (
            .in0(N__23987),
            .in1(N__25064),
            .in2(N__23883),
            .in3(N__24524),
            .lcout(un113_pixel_4_0_15__N_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_6_bm_2_LC_8_15_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_6_bm_2_LC_8_15_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_6_bm_2_LC_8_15_5.LUT_INIT=16'b1110110001001100;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_6_bm_2_LC_8_15_5 (
            .in0(N__25067),
            .in1(N__21650),
            .in2(N__24862),
            .in3(N__21944),
            .lcout(),
            .ltout(un115_pixel_6_bm_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_2_LC_8_15_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_2_LC_8_15_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_6_ns_2_LC_8_15_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_6_ns_2_LC_8_15_6 (
            .in0(N__24170),
            .in1(_gnd_net_),
            .in2(N__19811),
            .in3(N__19799),
            .lcout(N_1330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_6_am_2_LC_8_15_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_6_am_2_LC_8_15_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_6_am_2_LC_8_15_7.LUT_INIT=16'b0010001000110011;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_6_am_2_LC_8_15_7 (
            .in0(N__25066),
            .in1(N__24839),
            .in2(_gnd_net_),
            .in3(N__25214),
            .lcout(un115_pixel_6_am_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__SUM4_3_i_a2_LC_9_1_0.C_ON=1'b1;
    defparam un113_pixel_4_0_15__SUM4_3_i_a2_LC_9_1_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__SUM4_3_i_a2_LC_9_1_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 un113_pixel_4_0_15__SUM4_3_i_a2_LC_9_1_0 (
            .in0(_gnd_net_),
            .in1(N__22257),
            .in2(_gnd_net_),
            .in3(N__22319),
            .lcout(N_56),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DC_LC_9_1_1.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DC_LC_9_1_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DC_LC_9_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DC_LC_9_1_1 (
            .in0(_gnd_net_),
            .in1(N__19793),
            .in2(N__21746),
            .in3(N__19760),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDE_LC_9_1_2.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDE_LC_9_1_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDE_LC_9_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDE_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(N__21926),
            .in2(N__19682),
            .in3(N__19739),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS72T_LC_9_1_3.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS72T_LC_9_1_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS72T_LC_9_1_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS72T_LC_9_1_3 (
            .in0(N__19716),
            .in1(N__19688),
            .in2(N__21776),
            .in3(N__19724),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_LC_9_1_4.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_LC_9_1_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_LC_9_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_LC_9_1_4 (
            .in0(N__19681),
            .in1(N__21761),
            .in2(N__22094),
            .in3(N__19721),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_0_LC_9_1_5.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_0_LC_9_1_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_0_LC_9_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_0_LC_9_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19677),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_LC_9_1_6.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_LC_9_1_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_LC_9_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_LC_9_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21742),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_9_2_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_9_2_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_9_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_9_2_0 (
            .in0(_gnd_net_),
            .in1(N__22720),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_9_2_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_9_2_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_9_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_9_2_1 (
            .in0(_gnd_net_),
            .in1(N__19871),
            .in2(N__19832),
            .in3(N__19865),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_9_2_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_9_2_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_9_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_9_2_2 (
            .in0(_gnd_net_),
            .in1(N__19862),
            .in2(N__19856),
            .in3(N__19847),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_9_2_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_9_2_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_9_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_9_2_3 (
            .in0(_gnd_net_),
            .in1(N__19844),
            .in2(N__20234),
            .in3(N__19838),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_9_2_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_9_2_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_9_2_4.LUT_INIT=16'b0101010110101010;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_9_2_4 (
            .in0(N__22076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19835),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_9_2_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_9_2_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_9_2_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_2_LC_9_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22251),
            .lcout(un5_visiblex_i_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_2110_i_LC_9_3_1.C_ON=1'b0;
    defparam column_1_N_2110_i_LC_9_3_1.SEQ_MODE=4'b0000;
    defparam column_1_N_2110_i_LC_9_3_1.LUT_INIT=16'b0001000110111011;
    LogicCell40 column_1_N_2110_i_LC_9_3_1 (
            .in0(N__22023),
            .in1(N__22271),
            .in2(_gnd_net_),
            .in3(N__19820),
            .lcout(N_2110_i),
            .ltout(N_2110_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_9_3_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_9_3_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_9_3_2.LUT_INIT=16'b0000111111110000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_9_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19823),
            .in3(N__20246),
            .lcout(if_generate_plus_mult1_un54_sum_axb_2_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_9_3_3.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_9_3_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_m_5_LC_9_3_3 (
            .in0(N__22022),
            .in1(N__22270),
            .in2(_gnd_net_),
            .in3(N__19819),
            .lcout(if_generate_plus_mult1_un47_sum_m_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_9_3_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_9_3_4.LUT_INIT=16'b0011100101101100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_9_3_4 (
            .in0(N__22067),
            .in1(N__20337),
            .in2(N__22745),
            .in3(N__22730),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_9_3_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_9_3_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_9_3_5.LUT_INIT=16'b1110000101001011;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_9_3_5 (
            .in0(N__22024),
            .in1(N__22373),
            .in2(N__20349),
            .in3(N__20240),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_3_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_3_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_3_6.LUT_INIT=16'b0000010111111010;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_3_6 (
            .in0(N__22252),
            .in1(N__22162),
            .in2(N__22320),
            .in3(N__22021),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_9_3_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_9_3_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_9_3_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_9_3_7 (
            .in0(N__22025),
            .in1(N__20225),
            .in2(N__20350),
            .in3(N__22385),
            .lcout(if_generate_plus_mult1_un54_sum_axb_3_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_9_0_LC_9_4_0.C_ON=1'b0;
    defparam ScreenBuffer_0_9_0_LC_9_4_0.SEQ_MODE=4'b1000;
    defparam ScreenBuffer_0_9_0_LC_9_4_0.LUT_INIT=16'b1011111110000000;
    LogicCell40 ScreenBuffer_0_9_0_LC_9_4_0 (
            .in0(N__20216),
            .in1(N__20084),
            .in2(N__20039),
            .in3(N__20011),
            .lcout(ScreenBuffer_0_9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19983),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_9_4_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_9_4_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_9_4_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_9_4_2 (
            .in0(_gnd_net_),
            .in1(N__20278),
            .in2(_gnd_net_),
            .in3(N__19886),
            .lcout(if_generate_plus_mult1_un54_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_9_4_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_9_4_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_9_4_7.LUT_INIT=16'b1001100111000011;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_9_4_7 (
            .in0(N__19880),
            .in1(N__20344),
            .in2(N__22349),
            .in3(N__22032),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_9_5_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_9_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__22449),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_9_5_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_9_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__20363),
            .in2(N__20290),
            .in3(N__20354),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_5_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(N__20351),
            .in2(N__20312),
            .in3(N__20300),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_9_5_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_9_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_9_5_3 (
            .in0(N__20565),
            .in1(N__20297),
            .in2(N__20291),
            .in3(N__20267),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_9_5_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_9_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_s_5_LC_9_5_4 (
            .in0(_gnd_net_),
            .in1(N__20264),
            .in2(_gnd_net_),
            .in3(N__20258),
            .lcout(if_generate_plus_mult1_un54_sum_s_5),
            .ltout(if_generate_plus_mult1_un54_sum_s_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_9_5_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_9_5_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_9_5_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20255),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_0_LC_9_5_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_0_LC_9_5_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_0_LC_9_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_0_LC_9_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22492),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(N__23081),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PU8_LC_9_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PU8_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PU8_LC_9_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PU8_LC_9_6_1 (
            .in0(_gnd_net_),
            .in1(N__20464),
            .in2(N__20450),
            .in3(N__20252),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSC_LC_9_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSC_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSC_LC_9_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSC_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(N__22496),
            .in2(N__22562),
            .in3(N__20249),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIU5ODU_LC_9_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIU5ODU_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIU5ODU_LC_9_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIU5ODU_LC_9_6_3 (
            .in0(N__20620),
            .in1(N__20465),
            .in2(N__22544),
            .in3(N__20456),
            .lcout(charx_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_LC_9_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_LC_9_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_LC_9_6_4 (
            .in0(_gnd_net_),
            .in1(N__22514),
            .in2(_gnd_net_),
            .in3(N__20453),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_9_6_7.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_9_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_9_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22607),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_7_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_7_0 (
            .in0(_gnd_net_),
            .in1(N__22664),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RF_LC_9_7_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RF_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RF_LC_9_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RF_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(N__20602),
            .in2(N__20630),
            .in3(N__20432),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNO_LC_9_7_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNO_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNO_LC_9_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNO_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(N__20621),
            .in2(N__20429),
            .in3(N__20411),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI1QD7R1_LC_9_7_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI1QD7R1_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI1QD7R1_LC_9_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI1QD7R1_LC_9_7_3 (
            .in0(N__20380),
            .in1(N__20603),
            .in2(N__20408),
            .in3(N__20393),
            .lcout(charx_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHU_LC_9_7_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHU_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHU_LC_9_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHU_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__20390),
            .in2(_gnd_net_),
            .in3(N__20384),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_2096_i_LC_9_7_5.C_ON=1'b0;
    defparam column_1_N_2096_i_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam column_1_N_2096_i_LC_9_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_N_2096_i_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22461),
            .lcout(N_2096_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_7_6.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23089),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_0_LC_9_7_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_0_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_0_LC_9_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_0_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20619),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_8_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__22618),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_9_8_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_9_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__20594),
            .in2(N__20525),
            .in3(N__20579),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_9_8_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_9_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__20572),
            .in2(N__20549),
            .in3(N__20528),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_9_8_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_9_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_9_8_3 (
            .in0(N__25870),
            .in1(N__20524),
            .in2(N__20507),
            .in3(N__20489),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_9_8_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_9_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_s_5_LC_9_8_4 (
            .in0(_gnd_net_),
            .in1(N__20486),
            .in2(_gnd_net_),
            .in3(N__20477),
            .lcout(column_1_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_i_sbtinv_3_LC_9_8_5.C_ON=1'b0;
    defparam column_1_i_sbtinv_3_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam column_1_i_sbtinv_3_LC_9_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_i_sbtinv_3_LC_9_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25869),
            .lcout(column_1_i_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_9_9_0.C_ON=1'b0;
    defparam PixelZ0_LC_9_9_0.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_9_9_0.LUT_INIT=16'b0100000001010101;
    LogicCell40 PixelZ0_LC_9_9_0 (
            .in0(N__21095),
            .in1(N__21083),
            .in2(N__21278),
            .in3(N__21077),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21054),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_5_LC_9_9_1.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_5_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_5_LC_9_9_1.LUT_INIT=16'b0001100000000000;
    LogicCell40 un113_pixel_7_1_7__g0_5_LC_9_9_1 (
            .in0(N__21023),
            .in1(N__20691),
            .in2(N__20884),
            .in3(N__24725),
            .lcout(N_3078_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_i_sbtinv_2_LC_9_9_2.C_ON=1'b0;
    defparam column_1_i_sbtinv_2_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam column_1_i_sbtinv_2_LC_9_9_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_i_sbtinv_2_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25285),
            .lcout(column_1_i_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_12_LC_9_9_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_12_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_12_LC_9_9_3.LUT_INIT=16'b1100010111001111;
    LogicCell40 un113_pixel_4_0_15__g0_12_LC_9_9_3 (
            .in0(N__23877),
            .in1(N__21482),
            .in2(N__24853),
            .in3(N__21494),
            .lcout(),
            .ltout(N_1297_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_1_0_LC_9_9_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_1_0_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_1_0_LC_9_9_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 un113_pixel_4_0_15__g0_1_0_LC_9_9_4 (
            .in0(N__24117),
            .in1(_gnd_net_),
            .in2(N__20999),
            .in3(N__21458),
            .lcout(N_4564_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_14_LC_9_9_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_14_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_14_LC_9_9_5.LUT_INIT=16'b1000001000000000;
    LogicCell40 un113_pixel_4_0_15__g0_14_LC_9_9_5 (
            .in0(N__20900),
            .in1(N__20692),
            .in2(N__20885),
            .in3(N__23335),
            .lcout(font_un67_pixel_ac0_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_4_0_0_LC_9_9_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_4_0_0_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_4_0_0_LC_9_9_6.LUT_INIT=16'b0110011001100110;
    LogicCell40 un113_pixel_4_0_15__g0_4_0_0_LC_9_9_6 (
            .in0(N__20984),
            .in1(N__20939),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un113_pixel_4_0_15__g0_4_0Z0Z_0),
            .ltout(un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_13_LC_9_9_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_13_LC_9_9_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_13_LC_9_9_7.LUT_INIT=16'b0000000000101101;
    LogicCell40 un113_pixel_4_0_15__g0_13_LC_9_9_7 (
            .in0(N__20865),
            .in1(N__20693),
            .in2(N__20633),
            .in3(N__23336),
            .lcout(font_un64_pixel_ac0_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJIDRG11_0_0_LC_9_10_0.C_ON=1'b0;
    defparam beamY_RNIJIDRG11_0_0_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIJIDRG11_0_0_LC_9_10_0.LUT_INIT=16'b0010111100100000;
    LogicCell40 beamY_RNIJIDRG11_0_0_LC_9_10_0 (
            .in0(N__25035),
            .in1(N__24229),
            .in2(N__24804),
            .in3(N__25759),
            .lcout(beamY_RNIJIDRG11_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_4_LC_9_10_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_4_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_4_LC_9_10_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 un113_pixel_4_0_15__g0_4_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(N__21296),
            .in2(N__21104),
            .in3(N__21602),
            .lcout(N_1342),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_5_4_LC_9_10_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_5_4_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_5_4_LC_9_10_2.LUT_INIT=16'b1111111011111111;
    LogicCell40 un113_pixel_4_0_15__g0_5_4_LC_9_10_2 (
            .in0(N__21269),
            .in1(N__21260),
            .in2(N__21245),
            .in3(N__21236),
            .lcout(),
            .ltout(un113_pixel_4_0_15__g0_5Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_11_LC_9_10_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_11_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_11_LC_9_10_3.LUT_INIT=16'b1111001011110111;
    LogicCell40 un113_pixel_4_0_15__g0_11_LC_9_10_3 (
            .in0(N__21221),
            .in1(N__21185),
            .in2(N__21209),
            .in3(N__21173),
            .lcout(N_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g2_0_LC_9_10_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g2_0_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g2_0_LC_9_10_4.LUT_INIT=16'b0111011100110011;
    LogicCell40 un113_pixel_4_0_15__g2_0_LC_9_10_4 (
            .in0(N__25036),
            .in1(N__24752),
            .in2(_gnd_net_),
            .in3(N__25225),
            .lcout(),
            .ltout(un113_pixel_4_0_15__g2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_20_LC_9_10_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_20_LC_9_10_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_20_LC_9_10_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 un113_pixel_4_0_15__g0_20_LC_9_10_5 (
            .in0(N__21410),
            .in1(N__23343),
            .in2(N__21200),
            .in3(N__21197),
            .lcout(un115_pixel_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_0_0_LC_9_10_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_0_0_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_0_0_LC_9_10_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 un113_pixel_4_0_15__g0_0_0_LC_9_10_6 (
            .in0(N__23344),
            .in1(N__21692),
            .in2(_gnd_net_),
            .in3(N__21179),
            .lcout(N_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_10_LC_9_11_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_10_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_10_LC_9_11_0.LUT_INIT=16'b1110110101001000;
    LogicCell40 un113_pixel_4_0_15__g0_10_LC_9_11_0 (
            .in0(N__21167),
            .in1(N__21134),
            .in2(N__21122),
            .in3(N__24251),
            .lcout(N_2075),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_2_s_6_LC_9_11_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_2_s_6_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_2_s_6_LC_9_11_1.LUT_INIT=16'b0001000100110011;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_2_s_6_LC_9_11_1 (
            .in0(N__25398),
            .in1(N__24748),
            .in2(_gnd_net_),
            .in3(N__21316),
            .lcout(),
            .ltout(un115_pixel_2_s_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_2_d_0_6_LC_9_11_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_2_d_0_6_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_2_d_0_6_LC_9_11_2.LUT_INIT=16'b0101010101110010;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_2_d_0_6_LC_9_11_2 (
            .in0(N__23878),
            .in1(N__23994),
            .in2(N__21449),
            .in3(N__24540),
            .lcout(),
            .ltout(un115_pixel_2_d_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_3_bm_6_LC_9_11_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_3_bm_6_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_3_bm_6_LC_9_11_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_3_bm_6_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(N__21365),
            .in2(N__21446),
            .in3(N__25042),
            .lcout(un115_pixel_3_bm_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_RNIF16BSN1_1_LC_9_11_5.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_RNIF16BSN1_1_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_e_0_RNIF16BSN1_1_LC_9_11_5.LUT_INIT=16'b1110000001000000;
    LogicCell40 ScreenBuffer_1_0_e_0_RNIF16BSN1_1_LC_9_11_5 (
            .in0(N__25742),
            .in1(N__21436),
            .in2(N__23464),
            .in3(N__21421),
            .lcout(ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_23_LC_9_11_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_23_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_23_LC_9_11_6.LUT_INIT=16'b0000010000001100;
    LogicCell40 un113_pixel_4_0_15__g0_23_LC_9_11_6 (
            .in0(N__21302),
            .in1(N__24146),
            .in2(N__24827),
            .in3(N__23844),
            .lcout(N_1_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_RNIHFGISN1_1_LC_9_11_7.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_RNIHFGISN1_1_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_e_0_RNIHFGISN1_1_LC_9_11_7.LUT_INIT=16'b1110000001000000;
    LogicCell40 ScreenBuffer_1_1_e_0_RNIHFGISN1_1_LC_9_11_7 (
            .in0(N__25741),
            .in1(N__21403),
            .in2(N__23465),
            .in3(N__21385),
            .lcout(ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__m8_LC_9_12_0.C_ON=1'b0;
    defparam un113_pixel_3_0_11__m8_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__m8_LC_9_12_0.LUT_INIT=16'b0010101111101111;
    LogicCell40 un113_pixel_3_0_11__m8_LC_9_12_0 (
            .in0(N__24474),
            .in1(N__23790),
            .in2(N__24833),
            .in3(N__23956),
            .lcout(m8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_RNISDB6RM_1_LC_9_12_1.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_RNISDB6RM_1_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_e_0_RNISDB6RM_1_LC_9_12_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 ScreenBuffer_1_0_e_0_RNISDB6RM_1_LC_9_12_1 (
            .in0(N__25518),
            .in1(N__21355),
            .in2(_gnd_net_),
            .in3(N__21340),
            .lcout(ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1),
            .ltout(ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__un115_pixel_5_s_7_LC_9_12_2.C_ON=1'b0;
    defparam un113_pixel_3_0_11__un115_pixel_5_s_7_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__un115_pixel_5_s_7_LC_9_12_2.LUT_INIT=16'b1100000000000000;
    LogicCell40 un113_pixel_3_0_11__un115_pixel_5_s_7_LC_9_12_2 (
            .in0(_gnd_net_),
            .in1(N__23302),
            .in2(N__21305),
            .in3(N__25415),
            .lcout(un115_pixel_5_s_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__g1_LC_9_12_3.C_ON=1'b0;
    defparam un113_pixel_3_0_11__g1_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__g1_LC_9_12_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un113_pixel_3_0_11__g1_LC_9_12_3 (
            .in0(N__23957),
            .in1(N__24996),
            .in2(_gnd_net_),
            .in3(N__24475),
            .lcout(un113_pixel_3_0_11__gZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVDIFFI1_0_LC_9_12_4.C_ON=1'b0;
    defparam beamY_RNIVDIFFI1_0_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIVDIFFI1_0_LC_9_12_4.LUT_INIT=16'b1100101111000111;
    LogicCell40 beamY_RNIVDIFFI1_0_LC_9_12_4 (
            .in0(N__24473),
            .in1(N__23789),
            .in2(N__24832),
            .in3(N__23955),
            .lcout(beamY_RNIVDIFFI1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIB3R6U63_0_LC_9_12_5.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIB3R6U63_0_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIB3R6U63_0_LC_9_12_5.LUT_INIT=16'b1110000001010000;
    LogicCell40 ScreenBuffer_0_7_RNIB3R6U63_0_LC_9_12_5 (
            .in0(N__23954),
            .in1(N__24995),
            .in2(N__23845),
            .in3(N__24471),
            .lcout(ScreenBuffer_0_7_RNIB3R6U63Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__un115_pixel_5_am_7_LC_9_12_6.C_ON=1'b0;
    defparam un113_pixel_3_0_11__un115_pixel_5_am_7_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__un115_pixel_5_am_7_LC_9_12_6.LUT_INIT=16'b0101011111110010;
    LogicCell40 un113_pixel_3_0_11__un115_pixel_5_am_7_LC_9_12_6 (
            .in0(N__24472),
            .in1(N__23788),
            .in2(N__23345),
            .in3(N__23429),
            .lcout(),
            .ltout(un115_pixel_5_am_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__un115_pixel_5_ns_7_LC_9_12_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__un115_pixel_5_ns_7_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__un115_pixel_5_ns_7_LC_9_12_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_3_0_11__un115_pixel_5_ns_7_LC_9_12_7 (
            .in0(_gnd_net_),
            .in1(N__21554),
            .in2(N__21548),
            .in3(N__21545),
            .lcout(N_1288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g1_0_LC_9_13_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g1_0_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g1_0_LC_9_13_0.LUT_INIT=16'b0101100100000100;
    LogicCell40 un113_pixel_4_0_15__g1_0_LC_9_13_0 (
            .in0(N__25057),
            .in1(N__21533),
            .in2(N__23033),
            .in3(N__24510),
            .lcout(un113_pixel_4_0_15__g1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__m9_LC_9_13_1.C_ON=1'b0;
    defparam un113_pixel_7_1_7__m9_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__m9_LC_9_13_1.LUT_INIT=16'b1000000001100000;
    LogicCell40 un113_pixel_7_1_7__m9_LC_9_13_1 (
            .in0(N__24511),
            .in1(N__25056),
            .in2(N__23866),
            .in3(N__23971),
            .lcout(m9),
            .ltout(m9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICJUESD2_0_0_LC_9_13_2.C_ON=1'b0;
    defparam beamY_RNICJUESD2_0_0_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam beamY_RNICJUESD2_0_0_LC_9_13_2.LUT_INIT=16'b0000101001011111;
    LogicCell40 beamY_RNICJUESD2_0_0_LC_9_13_2 (
            .in0(N__24826),
            .in1(_gnd_net_),
            .in2(N__21470),
            .in3(N__21467),
            .lcout(beamY_RNICJUESD2_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m6_LC_9_13_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m6_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m6_LC_9_13_3.LUT_INIT=16'b1001000000100000;
    LogicCell40 un113_pixel_4_0_15__m6_LC_9_13_3 (
            .in0(N__24512),
            .in1(N__25058),
            .in2(N__23865),
            .in3(N__23970),
            .lcout(m6),
            .ltout(m6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICJUESD2_0_LC_9_13_4.C_ON=1'b0;
    defparam beamY_RNICJUESD2_0_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam beamY_RNICJUESD2_0_LC_9_13_4.LUT_INIT=16'b1010111100000101;
    LogicCell40 beamY_RNICJUESD2_0_LC_9_13_4 (
            .in0(N__24825),
            .in1(_gnd_net_),
            .in2(N__21461),
            .in3(N__21719),
            .lcout(beamY_RNICJUESD2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_8_LC_9_13_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_8_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_8_LC_9_13_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 un113_pixel_4_0_15__g0_8_LC_9_13_5 (
            .in0(N__24828),
            .in1(N__21644),
            .in2(_gnd_net_),
            .in3(N__21638),
            .lcout(),
            .ltout(N_4562_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_7_LC_9_13_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_7_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_7_LC_9_13_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_4_0_15__g0_7_LC_9_13_6 (
            .in0(_gnd_net_),
            .in1(N__21632),
            .in2(N__21605),
            .in3(N__21575),
            .lcout(N_1340_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1H36941_0_LC_9_13_7.C_ON=1'b0;
    defparam beamY_RNI1H36941_0_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI1H36941_0_LC_9_13_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 beamY_RNI1H36941_0_LC_9_13_7 (
            .in0(N__21560),
            .in1(_gnd_net_),
            .in2(N__24162),
            .in3(N__21593),
            .lcout(beamY_RNI1H36941Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x0_0_LC_9_14_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x0_0_LC_9_14_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x0_0_LC_9_14_0.LUT_INIT=16'b0101000101010101;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_5_ns_x0_0_LC_9_14_0 (
            .in0(N__24506),
            .in1(N__23434),
            .in2(N__24855),
            .in3(N__25030),
            .lcout(un115_pixel_5_ns_x0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x1_0_LC_9_14_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x1_0_LC_9_14_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_x1_0_LC_9_14_1.LUT_INIT=16'b1111000011110111;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_5_ns_x1_0_LC_9_14_1 (
            .in0(N__23435),
            .in1(N__25013),
            .in2(N__24856),
            .in3(N__24507),
            .lcout(un115_pixel_5_ns_x1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__font_un125_pixel_1_bm_LC_9_14_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__font_un125_pixel_1_bm_LC_9_14_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__font_un125_pixel_1_bm_LC_9_14_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 un113_pixel_4_0_15__font_un125_pixel_1_bm_LC_9_14_2 (
            .in0(N__23353),
            .in1(N__21656),
            .in2(_gnd_net_),
            .in3(N__21671),
            .lcout(font_un125_pixel_1_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_2_0_3__m7_LC_9_14_3.C_ON=1'b0;
    defparam un113_pixel_2_0_3__m7_LC_9_14_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_2_0_3__m7_LC_9_14_3.LUT_INIT=16'b0001000110101010;
    LogicCell40 un113_pixel_2_0_3__m7_LC_9_14_3 (
            .in0(N__23968),
            .in1(N__25014),
            .in2(_gnd_net_),
            .in3(N__24508),
            .lcout(un113_pixel_2_0_3__N_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_6_1_5__m10_LC_9_14_4.C_ON=1'b0;
    defparam un113_pixel_6_1_5__m10_LC_9_14_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_6_1_5__m10_LC_9_14_4.LUT_INIT=16'b0000000011100000;
    LogicCell40 un113_pixel_6_1_5__m10_LC_9_14_4 (
            .in0(N__24509),
            .in1(N__23969),
            .in2(N__23885),
            .in3(N__25031),
            .lcout(),
            .ltout(un113_pixel_6_1_5__N_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICJUESD2_2_0_LC_9_14_5.C_ON=1'b0;
    defparam beamY_RNICJUESD2_2_0_LC_9_14_5.SEQ_MODE=4'b0000;
    defparam beamY_RNICJUESD2_2_0_LC_9_14_5.LUT_INIT=16'b0000101001001110;
    LogicCell40 beamY_RNICJUESD2_2_0_LC_9_14_5 (
            .in0(N__24816),
            .in1(N__23864),
            .in2(N__21569),
            .in3(N__21566),
            .lcout(beamY_RNICJUESD2_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__m12_LC_9_14_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__m12_LC_9_14_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__m12_LC_9_14_6.LUT_INIT=16'b0111011100110011;
    LogicCell40 un113_pixel_4_0_15__m12_LC_9_14_6 (
            .in0(N__25012),
            .in1(N__23859),
            .in2(_gnd_net_),
            .in3(N__23967),
            .lcout(m12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__m17_LC_9_14_7.C_ON=1'b0;
    defparam un113_pixel_3_0_11__m17_LC_9_14_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__m17_LC_9_14_7.LUT_INIT=16'b0010000010010000;
    LogicCell40 un113_pixel_3_0_11__m17_LC_9_14_7 (
            .in0(N__23966),
            .in1(N__25011),
            .in2(N__23884),
            .in3(N__24505),
            .lcout(m17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_ns_0_LC_9_15_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_ns_0_LC_9_15_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_5_ns_ns_0_LC_9_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_5_ns_ns_0_LC_9_15_0 (
            .in0(N__21713),
            .in1(N__21707),
            .in2(_gnd_net_),
            .in3(N__21701),
            .lcout(),
            .ltout(N_1325_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_7_bm_0_LC_9_15_1.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_7_bm_0_LC_9_15_1.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_7_bm_0_LC_9_15_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_7_bm_0_LC_9_15_1 (
            .in0(_gnd_net_),
            .in1(N__24161),
            .in2(N__21695),
            .in3(N__21932),
            .lcout(un115_pixel_7_bm_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_4_3_LC_9_15_2.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_4_3_LC_9_15_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_4_3_LC_9_15_2.LUT_INIT=16'b0110011001010101;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_4_3_LC_9_15_2 (
            .in0(N__24821),
            .in1(N__25074),
            .in2(_gnd_net_),
            .in3(N__25212),
            .lcout(),
            .ltout(N_1315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_6_3_LC_9_15_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_6_3_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_6_3_LC_9_15_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_6_3_LC_9_15_3 (
            .in0(_gnd_net_),
            .in1(N__24160),
            .in2(N__21680),
            .in3(N__21677),
            .lcout(N_1329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_1_3_LC_9_15_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_1_3_LC_9_15_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_1_3_LC_9_15_4.LUT_INIT=16'b0111000010110000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_1_3_LC_9_15_4 (
            .in0(N__25070),
            .in1(N__25151),
            .in2(N__24857),
            .in3(N__24535),
            .lcout(),
            .ltout(N_1294_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_3_ns_3_LC_9_15_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_3_ns_3_LC_9_15_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_3_ns_3_LC_9_15_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_3_ns_3_LC_9_15_5 (
            .in0(_gnd_net_),
            .in1(N__24159),
            .in2(N__21665),
            .in3(N__21662),
            .lcout(N_1308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_5_d_2_LC_9_15_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_5_d_2_LC_9_15_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_5_d_2_LC_9_15_6.LUT_INIT=16'b0000000010000010;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_5_d_2_LC_9_15_6 (
            .in0(N__23860),
            .in1(N__24002),
            .in2(N__24858),
            .in3(N__24536),
            .lcout(un115_pixel_5_d_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMR86ES2_0_LC_9_15_7.C_ON=1'b0;
    defparam beamY_RNIMR86ES2_0_LC_9_15_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIMR86ES2_0_LC_9_15_7.LUT_INIT=16'b0011011111000100;
    LogicCell40 beamY_RNIMR86ES2_0_LC_9_15_7 (
            .in0(N__25213),
            .in1(N__24817),
            .in2(N__25082),
            .in3(N__21943),
            .lcout(beamY_RNIMR86ES2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_1_0.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_1_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_1_0 (
            .in0(_gnd_net_),
            .in1(N__22330),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9254_LC_11_1_1.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9254_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9254_LC_11_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9254_LC_11_1_1 (
            .in0(_gnd_net_),
            .in1(N__21731),
            .in2(_gnd_net_),
            .in3(N__21917),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIA464_LC_11_1_2.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIA464_LC_11_1_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIA464_LC_11_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIA464_LC_11_1_2 (
            .in0(_gnd_net_),
            .in1(N__21725),
            .in2(N__21904),
            .in3(N__21764),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_1_3.C_ON=1'b1;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_1_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_1_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_1_3 (
            .in0(_gnd_net_),
            .in1(N__22088),
            .in2(_gnd_net_),
            .in3(N__21752),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_1_4.C_ON=1'b0;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_1_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_1_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21749),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_11_1_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_11_1_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_11_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_3_LC_11_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22086),
            .lcout(chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_1_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_1_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_1_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_2_LC_11_1_6 (
            .in0(N__22087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_11_2_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_11_2_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_11_2_4.LUT_INIT=16'b0101010100110011;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_11_2_4 (
            .in0(N__22193),
            .in1(N__22163),
            .in2(_gnd_net_),
            .in3(N__22071),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_11_3_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_11_3_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_11_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_11_3_0 (
            .in0(_gnd_net_),
            .in1(N__22736),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_11_3_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_11_3_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_11_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_11_3_1 (
            .in0(_gnd_net_),
            .in1(N__22202),
            .in2(N__22092),
            .in3(N__22376),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_11_3_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_11_3_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_11_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_11_3_2 (
            .in0(_gnd_net_),
            .in1(N__22100),
            .in2(N__21953),
            .in3(N__22361),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_11_3_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_11_3_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_11_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_11_3_3 (
            .in0(_gnd_net_),
            .in1(N__22358),
            .in2(N__22093),
            .in3(N__22334),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_11_3_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_11_3_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_11_3_4.LUT_INIT=16'b1000000001111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_11_3_4 (
            .in0(N__22259),
            .in1(N__22084),
            .in2(N__22331),
            .in3(N__22274),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_11_3_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_11_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_3_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22258),
            .lcout(un5_visiblex_i_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_11_3_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_11_3_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_11_3_6.LUT_INIT=16'b0001000111101110;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_11_3_6 (
            .in0(N__22192),
            .in1(N__22158),
            .in2(_gnd_net_),
            .in3(N__22077),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_charx_if_generate_plus_mult1_un26_sum_axb_3_i_LC_11_4_2.C_ON=1'b0;
    defparam column_1_charx_if_generate_plus_mult1_un26_sum_axb_3_i_LC_11_4_2.SEQ_MODE=4'b0000;
    defparam column_1_charx_if_generate_plus_mult1_un26_sum_axb_3_i_LC_11_4_2.LUT_INIT=16'b0011001100110011;
    LogicCell40 column_1_charx_if_generate_plus_mult1_un26_sum_axb_3_i_LC_11_4_2 (
            .in0(_gnd_net_),
            .in1(N__22085),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un26_sum_axb_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(N__22620),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__22525),
            .in2(N__22472),
            .in3(N__22547),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__22813),
            .in2(N__22397),
            .in3(N__22529),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI0CRJF_LC_11_5_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI0CRJF_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI0CRJF_LC_11_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI0CRJF_LC_11_5_3 (
            .in0(N__22491),
            .in1(N__22526),
            .in2(N__22850),
            .in3(N__22502),
            .lcout(charx_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_LC_11_5_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_LC_11_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(N__22838),
            .in2(_gnd_net_),
            .in3(N__22499),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_11_5_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_11_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_11_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22463),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_11_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_11_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__22460),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_11_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_11_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__22406),
            .in2(N__22682),
            .in3(N__22388),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_11_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_11_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_11_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(N__22778),
            .in2(N__22862),
            .in3(N__22841),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNIU99G8_LC_11_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNIU99G8_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNIU99G8_LC_11_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNIU99G8_LC_11_6_3 (
            .in0(N__22812),
            .in1(N__22751),
            .in2(N__22793),
            .in3(N__22832),
            .lcout(charx_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_11_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_11_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(N__22829),
            .in2(_gnd_net_),
            .in3(N__22820),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINP73_LC_11_6_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINP73_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINP73_LC_11_6_5.LUT_INIT=16'b0011001100110011;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINP73_LC_11_6_5 (
            .in0(N__22792),
            .in1(N__22777),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_11_6_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_11_6_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_11_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_11_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22744),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_8_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__23146),
            .in2(_gnd_net_),
            .in3(N__25321),
            .lcout(if_generate_plus_mult1_un75_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_7.LUT_INIT=16'b0011001100110011;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_7 (
            .in0(_gnd_net_),
            .in1(N__22673),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_9_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(N__22672),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_9_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__22634),
            .in2(N__23042),
            .in3(N__22625),
            .lcout(if_generate_plus_mult1_un75_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_9_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__25400),
            .in2(N__23174),
            .in3(N__23159),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_9_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_9_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_9_3 (
            .in0(N__25688),
            .in1(N__23156),
            .in2(N__23150),
            .in3(N__23126),
            .lcout(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_9_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__23123),
            .in2(_gnd_net_),
            .in3(N__23111),
            .lcout(un6_rowlto1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un6_rowlto3_LC_11_9_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un6_rowlto3_LC_11_9_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un6_rowlto3_LC_11_9_5.LUT_INIT=16'b0000000100010001;
    LogicCell40 un113_pixel_4_0_15__un6_rowlto3_LC_11_9_5 (
            .in0(N__25401),
            .in1(N__25983),
            .in2(N__25512),
            .in3(N__25709),
            .lcout(un6_rowlt7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_11_9_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_11_9_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_11_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_i_LC_11_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23093),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPPD7L31_0_LC_11_10_1.C_ON=1'b0;
    defparam beamY_RNIPPD7L31_0_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIPPD7L31_0_LC_11_10_1.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_RNIPPD7L31_0_LC_11_10_1 (
            .in0(N__24834),
            .in1(N__23032),
            .in2(_gnd_net_),
            .in3(N__22919),
            .lcout(),
            .ltout(d_N_3_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2RNL4M2_0_LC_11_10_2.C_ON=1'b0;
    defparam beamY_RNI2RNL4M2_0_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2RNL4M2_0_LC_11_10_2.LUT_INIT=16'b0111000011111000;
    LogicCell40 beamY_RNI2RNL4M2_0_LC_11_10_2 (
            .in0(N__24001),
            .in1(N__23887),
            .in2(N__22907),
            .in3(N__24545),
            .lcout(beamY_RNI2RNL4M2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__currentchar_1_4_1_2_LC_11_10_3.C_ON=1'b0;
    defparam un113_pixel_3_0_11__currentchar_1_4_1_2_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__currentchar_1_4_1_2_LC_11_10_3.LUT_INIT=16'b1110111111100101;
    LogicCell40 un113_pixel_3_0_11__currentchar_1_4_1_2_LC_11_10_3 (
            .in0(N__25708),
            .in1(N__22904),
            .in2(N__25517),
            .in3(N__22889),
            .lcout(un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_10_RNIGDGIE9_0_LC_11_10_4.C_ON=1'b0;
    defparam ScreenBuffer_0_10_RNIGDGIE9_0_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_10_RNIGDGIE9_0_LC_11_10_4.LUT_INIT=16'b1001100100000000;
    LogicCell40 ScreenBuffer_0_10_RNIGDGIE9_0_LC_11_10_4 (
            .in0(N__23612),
            .in1(N__23529),
            .in2(_gnd_net_),
            .in3(N__23717),
            .lcout(ScreenBuffer_0_10_RNIGDGIE9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_11_RNI9RVK2F_0_LC_11_10_5.C_ON=1'b0;
    defparam ScreenBuffer_0_11_RNI9RVK2F_0_LC_11_10_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_11_RNI9RVK2F_0_LC_11_10_5.LUT_INIT=16'b0110011001101111;
    LogicCell40 ScreenBuffer_0_11_RNI9RVK2F_0_LC_11_10_5 (
            .in0(N__23530),
            .in1(N__23613),
            .in2(N__25987),
            .in3(N__23693),
            .lcout(),
            .ltout(currentchar_1_5_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_3_e_0_RNIR8DINK_0_LC_11_10_6.C_ON=1'b0;
    defparam ScreenBuffer_1_3_e_0_RNIR8DINK_0_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_3_e_0_RNIR8DINK_0_LC_11_10_6.LUT_INIT=16'b1000111110000101;
    LogicCell40 ScreenBuffer_1_3_e_0_RNIR8DINK_0_LC_11_10_6 (
            .in0(N__25968),
            .in1(N__23672),
            .in2(N__23660),
            .in3(N__23657),
            .lcout(ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_3_LC_11_11_0.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_3_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_3_LC_11_11_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 un113_pixel_7_1_7__g0_3_LC_11_11_0 (
            .in0(N__25078),
            .in1(N__23633),
            .in2(_gnd_net_),
            .in3(N__23621),
            .lcout(N_1303_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam currentchar_1_5_0_a2_0_1_LC_11_11_1.C_ON=1'b0;
    defparam currentchar_1_5_0_a2_0_1_LC_11_11_1.SEQ_MODE=4'b0000;
    defparam currentchar_1_5_0_a2_0_1_LC_11_11_1.LUT_INIT=16'b0011110000000000;
    LogicCell40 currentchar_1_5_0_a2_0_1_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(N__23614),
            .in2(N__23534),
            .in3(N__25969),
            .lcout(N_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_i_m2_LC_11_11_2.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_i_m2_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_i_m2_LC_11_11_2.LUT_INIT=16'b1011100011110000;
    LogicCell40 un113_pixel_7_1_7__g0_i_m2_LC_11_11_2 (
            .in0(N__25150),
            .in1(N__25080),
            .in2(N__23447),
            .in3(N__24544),
            .lcout(),
            .ltout(N_4581_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_0_LC_11_11_3.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_0_LC_11_11_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_0_LC_11_11_3.LUT_INIT=16'b1110001011110011;
    LogicCell40 un113_pixel_7_1_7__g0_0_LC_11_11_3 (
            .in0(N__25081),
            .in1(N__24835),
            .in2(N__23375),
            .in3(N__25226),
            .lcout(N_1296_0),
            .ltout(N_1296_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_16_x1_LC_11_11_4.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_16_x1_LC_11_11_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_16_x1_LC_11_11_4.LUT_INIT=16'b1111111000110010;
    LogicCell40 un113_pixel_4_0_15__g0_16_x1_LC_11_11_4 (
            .in0(N__24136),
            .in1(N__23359),
            .in2(N__23372),
            .in3(N__24010),
            .lcout(g0_16_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_16_x0_LC_11_11_5.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_16_x0_LC_11_11_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_16_x0_LC_11_11_5.LUT_INIT=16'b1010000010101100;
    LogicCell40 un113_pixel_4_0_15__g0_16_x0_LC_11_11_5 (
            .in0(N__24011),
            .in1(N__23369),
            .in2(N__23363),
            .in3(N__24137),
            .lcout(),
            .ltout(g0_16_x0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_16_ns_LC_11_11_6.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_16_ns_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_16_ns_LC_11_11_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 un113_pixel_4_0_15__g0_16_ns_LC_11_11_6 (
            .in0(_gnd_net_),
            .in1(N__24266),
            .in2(N__24260),
            .in3(N__24257),
            .lcout(N_4560_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_2_LC_11_12_0.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_2_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_2_LC_11_12_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 un113_pixel_4_0_15__g0_2_LC_11_12_0 (
            .in0(N__24135),
            .in1(N__24368),
            .in2(_gnd_net_),
            .in3(N__25157),
            .lcout(N_1309_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJIDRG11_0_LC_11_12_1.C_ON=1'b0;
    defparam beamY_RNIJIDRG11_0_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIJIDRG11_0_LC_11_12_1.LUT_INIT=16'b0111111101110000;
    LogicCell40 beamY_RNIJIDRG11_0_LC_11_12_1 (
            .in0(N__25075),
            .in1(N__24230),
            .in2(N__24854),
            .in3(N__25760),
            .lcout(),
            .ltout(beamY_RNIJIDRG11Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRG0LHO1_0_LC_11_12_2.C_ON=1'b0;
    defparam beamY_RNIRG0LHO1_0_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIRG0LHO1_0_LC_11_12_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNIRG0LHO1_0_LC_11_12_2 (
            .in0(_gnd_net_),
            .in1(N__24212),
            .in2(N__24200),
            .in3(N__24197),
            .lcout(beamY_RNIRG0LHO1Z0Z_0),
            .ltout(beamY_RNIRG0LHO1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_2_x0_LC_11_12_3.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_2_x0_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_2_x0_LC_11_12_3.LUT_INIT=16'b1101000111000000;
    LogicCell40 un113_pixel_7_1_7__g0_2_x0_LC_11_12_3 (
            .in0(N__24808),
            .in1(N__24131),
            .in2(N__24185),
            .in3(N__24181),
            .lcout(g0_2_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_2_x1_LC_11_12_4.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_2_x1_LC_11_12_4.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_2_x1_LC_11_12_4.LUT_INIT=16'b1111111000001110;
    LogicCell40 un113_pixel_7_1_7__g0_2_x1_LC_11_12_4 (
            .in0(N__24182),
            .in1(N__24809),
            .in2(N__24158),
            .in3(N__24035),
            .lcout(),
            .ltout(g0_2_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_7_1_7__g0_2_ns_LC_11_12_5.C_ON=1'b0;
    defparam un113_pixel_7_1_7__g0_2_ns_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam un113_pixel_7_1_7__g0_2_ns_LC_11_12_5.LUT_INIT=16'b1111001111000000;
    LogicCell40 un113_pixel_7_1_7__g0_2_ns_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(N__24029),
            .in2(N__24020),
            .in3(N__24017),
            .lcout(N_1331_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_3_0_11__m15_LC_11_12_6.C_ON=1'b0;
    defparam un113_pixel_3_0_11__m15_LC_11_12_6.SEQ_MODE=4'b0000;
    defparam un113_pixel_3_0_11__m15_LC_11_12_6.LUT_INIT=16'b1000000001010000;
    LogicCell40 un113_pixel_3_0_11__m15_LC_11_12_6 (
            .in0(N__24000),
            .in1(N__25076),
            .in2(N__23891),
            .in3(N__24543),
            .lcout(),
            .ltout(un113_pixel_3_0_11__N_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__g0_3_LC_11_12_7.C_ON=1'b0;
    defparam un113_pixel_4_0_15__g0_3_LC_11_12_7.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__g0_3_LC_11_12_7.LUT_INIT=16'b0001110100001100;
    LogicCell40 un113_pixel_4_0_15__g0_3_LC_11_12_7 (
            .in0(N__25077),
            .in1(N__24836),
            .in2(N__25229),
            .in3(N__25224),
            .lcout(N_4573_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un113_pixel_4_0_15__un115_pixel_3_am_2_LC_11_13_3.C_ON=1'b0;
    defparam un113_pixel_4_0_15__un115_pixel_3_am_2_LC_11_13_3.SEQ_MODE=4'b0000;
    defparam un113_pixel_4_0_15__un115_pixel_3_am_2_LC_11_13_3.LUT_INIT=16'b0111100011010000;
    LogicCell40 un113_pixel_4_0_15__un115_pixel_3_am_2_LC_11_13_3 (
            .in0(N__25149),
            .in1(N__25079),
            .in2(N__24863),
            .in3(N__24541),
            .lcout(un115_pixel_3_am_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_12_9_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_12_9_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_12_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_12_9_0 (
            .in0(_gnd_net_),
            .in1(N__24362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_12_9_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_12_9_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_12_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_12_9_1 (
            .in0(_gnd_net_),
            .in1(N__24305),
            .in2(N__24314),
            .in3(N__25686),
            .lcout(G_673),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_12_9_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_12_9_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_12_9_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_12_9_2 (
            .in0(_gnd_net_),
            .in1(N__25689),
            .in2(N__24299),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_12_9_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_12_9_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_12_9_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_12_9_3 (
            .in0(_gnd_net_),
            .in1(N__24281),
            .in2(N__24290),
            .in3(N__25687),
            .lcout(G_674),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_12_9_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_12_9_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_12_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_s_5_LC_12_9_4 (
            .in0(_gnd_net_),
            .in1(N__24275),
            .in2(_gnd_net_),
            .in3(N__24269),
            .lcout(un6_rowlto0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_LC_12_10_0.C_ON=1'b0;
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_LC_12_10_0.LUT_INIT=16'b1111101111101010;
    LogicCell40 ScreenBuffer_0_10_RNIB0Q4B12_0_LC_12_10_0 (
            .in0(N__25690),
            .in1(N__25966),
            .in2(N__25811),
            .in3(N__25819),
            .lcout(ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_0_LC_12_10_1.C_ON=1'b0;
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_0_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_10_RNIB0Q4B12_0_0_LC_12_10_1.LUT_INIT=16'b0011001000010000;
    LogicCell40 ScreenBuffer_0_10_RNIB0Q4B12_0_0_LC_12_10_1 (
            .in0(N__25967),
            .in1(N__25691),
            .in2(N__25823),
            .in3(N__25807),
            .lcout(),
            .ltout(ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_RNI1J74DN_0_LC_12_10_2.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_RNI1J74DN_0_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_e_0_RNI1J74DN_0_LC_12_10_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 ScreenBuffer_1_0_e_0_RNI1J74DN_0_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(N__25790),
            .in2(N__25781),
            .in3(N__25778),
            .lcout(ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_6_RNITJ4B17_0_LC_12_10_3.C_ON=1'b0;
    defparam ScreenBuffer_0_6_RNITJ4B17_0_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_6_RNITJ4B17_0_LC_12_10_3.LUT_INIT=16'b0000000010111111;
    LogicCell40 ScreenBuffer_0_6_RNITJ4B17_0_LC_12_10_3 (
            .in0(N__25397),
            .in1(N__25772),
            .in2(N__25513),
            .in3(N__25235),
            .lcout(ScreenBuffer_0_6_RNITJ4B17Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_LC_12_10_4.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_LC_12_10_4.LUT_INIT=16'b1111110111101100;
    LogicCell40 ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_LC_12_10_4 (
            .in0(N__25692),
            .in1(N__25478),
            .in2(N__25625),
            .in3(N__25633),
            .lcout(ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_0_LC_12_10_5.C_ON=1'b0;
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_0_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_0_LC_12_10_5.LUT_INIT=16'b0101010000010000;
    LogicCell40 ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_0_LC_12_10_5 (
            .in0(N__25477),
            .in1(N__25693),
            .in2(N__25637),
            .in3(N__25621),
            .lcout(),
            .ltout(ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_1_0_e_0_RNI3EKU1A_0_LC_12_10_6.C_ON=1'b0;
    defparam ScreenBuffer_1_0_e_0_RNI3EKU1A_0_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_1_0_e_0_RNI3EKU1A_0_LC_12_10_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 ScreenBuffer_1_0_e_0_RNI3EKU1A_0_LC_12_10_6 (
            .in0(_gnd_net_),
            .in1(N__25607),
            .in2(N__25601),
            .in3(N__25598),
            .lcout(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0),
            .ltout(ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ScreenBuffer_0_7_RNIS4U201_0_LC_12_10_7.C_ON=1'b0;
    defparam ScreenBuffer_0_7_RNIS4U201_0_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam ScreenBuffer_0_7_RNIS4U201_0_LC_12_10_7.LUT_INIT=16'b1101000111000000;
    LogicCell40 ScreenBuffer_0_7_RNIS4U201_0_LC_12_10_7 (
            .in0(N__25479),
            .in1(N__25402),
            .in2(N__25256),
            .in3(N__25253),
            .lcout(un115_pixel_5_am_sx_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
