// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 23 2015 17:44:05

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__14780;
    wire N__14779;
    wire N__14778;
    wire N__14771;
    wire N__14770;
    wire N__14769;
    wire N__14762;
    wire N__14761;
    wire N__14760;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14744;
    wire N__14743;
    wire N__14742;
    wire N__14735;
    wire N__14734;
    wire N__14733;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14700;
    wire N__14699;
    wire N__14698;
    wire N__14697;
    wire N__14696;
    wire N__14695;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14676;
    wire N__14671;
    wire N__14666;
    wire N__14663;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14631;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14623;
    wire N__14620;
    wire N__14619;
    wire N__14614;
    wire N__14611;
    wire N__14610;
    wire N__14609;
    wire N__14608;
    wire N__14607;
    wire N__14606;
    wire N__14601;
    wire N__14596;
    wire N__14595;
    wire N__14594;
    wire N__14593;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14545;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14494;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14411;
    wire N__14410;
    wire N__14409;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14384;
    wire N__14377;
    wire N__14376;
    wire N__14375;
    wire N__14374;
    wire N__14371;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14363;
    wire N__14362;
    wire N__14361;
    wire N__14360;
    wire N__14359;
    wire N__14358;
    wire N__14357;
    wire N__14356;
    wire N__14355;
    wire N__14352;
    wire N__14347;
    wire N__14344;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14326;
    wire N__14321;
    wire N__14316;
    wire N__14305;
    wire N__14296;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14262;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14148;
    wire N__14147;
    wire N__14140;
    wire N__14137;
    wire N__14136;
    wire N__14131;
    wire N__14128;
    wire N__14127;
    wire N__14124;
    wire N__14123;
    wire N__14120;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14102;
    wire N__14099;
    wire N__14092;
    wire N__14091;
    wire N__14090;
    wire N__14087;
    wire N__14086;
    wire N__14085;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14048;
    wire N__14041;
    wire N__14038;
    wire N__14037;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14002;
    wire N__13999;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13983;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13972;
    wire N__13971;
    wire N__13970;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13939;
    wire N__13930;
    wire N__13927;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13916;
    wire N__13913;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13892;
    wire N__13889;
    wire N__13882;
    wire N__13881;
    wire N__13880;
    wire N__13879;
    wire N__13876;
    wire N__13871;
    wire N__13870;
    wire N__13869;
    wire N__13868;
    wire N__13865;
    wire N__13860;
    wire N__13857;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13825;
    wire N__13820;
    wire N__13813;
    wire N__13810;
    wire N__13809;
    wire N__13808;
    wire N__13805;
    wire N__13804;
    wire N__13801;
    wire N__13800;
    wire N__13799;
    wire N__13796;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13777;
    wire N__13774;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13762;
    wire N__13761;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13710;
    wire N__13703;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13687;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13679;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13642;
    wire N__13641;
    wire N__13638;
    wire N__13637;
    wire N__13636;
    wire N__13635;
    wire N__13634;
    wire N__13633;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13607;
    wire N__13604;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire N__13572;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13547;
    wire N__13546;
    wire N__13543;
    wire N__13540;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13522;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13511;
    wire N__13510;
    wire N__13507;
    wire N__13504;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13500;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13482;
    wire N__13479;
    wire N__13474;
    wire N__13459;
    wire N__13456;
    wire N__13455;
    wire N__13454;
    wire N__13451;
    wire N__13450;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13426;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13418;
    wire N__13417;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13393;
    wire N__13390;
    wire N__13389;
    wire N__13388;
    wire N__13385;
    wire N__13384;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13314;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13293;
    wire N__13292;
    wire N__13291;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13276;
    wire N__13275;
    wire N__13274;
    wire N__13273;
    wire N__13272;
    wire N__13271;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13224;
    wire N__13223;
    wire N__13222;
    wire N__13221;
    wire N__13220;
    wire N__13219;
    wire N__13218;
    wire N__13217;
    wire N__13216;
    wire N__13215;
    wire N__13214;
    wire N__13213;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13179;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13168;
    wire N__13167;
    wire N__13166;
    wire N__13165;
    wire N__13164;
    wire N__13161;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13134;
    wire N__13131;
    wire N__13120;
    wire N__13119;
    wire N__13118;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13075;
    wire N__13074;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13067;
    wire N__13066;
    wire N__13061;
    wire N__13058;
    wire N__13057;
    wire N__13052;
    wire N__13049;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13024;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13008;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12907;
    wire N__12904;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12892;
    wire N__12889;
    wire N__12888;
    wire N__12887;
    wire N__12884;
    wire N__12879;
    wire N__12874;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12814;
    wire N__12811;
    wire N__12808;
    wire N__12805;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12766;
    wire N__12763;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12738;
    wire N__12737;
    wire N__12734;
    wire N__12729;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12690;
    wire N__12687;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12679;
    wire N__12678;
    wire N__12677;
    wire N__12674;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12662;
    wire N__12661;
    wire N__12658;
    wire N__12657;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12642;
    wire N__12637;
    wire N__12632;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12599;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12490;
    wire N__12487;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12343;
    wire N__12342;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12277;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12231;
    wire N__12228;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12204;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12189;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12168;
    wire N__12165;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12148;
    wire N__12147;
    wire N__12146;
    wire N__12145;
    wire N__12144;
    wire N__12139;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12115;
    wire N__12112;
    wire N__12107;
    wire N__12102;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12084;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12072;
    wire N__12069;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12049;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11995;
    wire N__11994;
    wire N__11991;
    wire N__11990;
    wire N__11987;
    wire N__11982;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11952;
    wire N__11951;
    wire N__11948;
    wire N__11947;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11917;
    wire N__11916;
    wire N__11915;
    wire N__11908;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11861;
    wire N__11858;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11811;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11797;
    wire N__11796;
    wire N__11795;
    wire N__11794;
    wire N__11793;
    wire N__11792;
    wire N__11791;
    wire N__11788;
    wire N__11787;
    wire N__11786;
    wire N__11781;
    wire N__11774;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11746;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11691;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11685;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11628;
    wire N__11625;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11422;
    wire N__11419;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11385;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11317;
    wire N__11314;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11199;
    wire N__11196;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11089;
    wire N__11088;
    wire N__11085;
    wire N__11078;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11044;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10988;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10952;
    wire N__10947;
    wire N__10942;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10919;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10912;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10885;
    wire N__10884;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10874;
    wire N__10871;
    wire N__10864;
    wire N__10861;
    wire N__10854;
    wire N__10851;
    wire N__10846;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10818;
    wire N__10817;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10799;
    wire N__10794;
    wire N__10793;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10713;
    wire N__10712;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10700;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10666;
    wire N__10665;
    wire N__10660;
    wire N__10655;
    wire N__10652;
    wire N__10645;
    wire N__10642;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10612;
    wire N__10607;
    wire N__10602;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10579;
    wire N__10576;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10555;
    wire N__10554;
    wire N__10553;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10545;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10533;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10500;
    wire N__10493;
    wire N__10474;
    wire N__10473;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10465;
    wire N__10464;
    wire N__10463;
    wire N__10462;
    wire N__10459;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10406;
    wire N__10399;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10363;
    wire N__10362;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10348;
    wire N__10345;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10329;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10248;
    wire N__10247;
    wire N__10244;
    wire N__10243;
    wire N__10240;
    wire N__10239;
    wire N__10236;
    wire N__10227;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10171;
    wire N__10170;
    wire N__10165;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10152;
    wire N__10151;
    wire N__10150;
    wire N__10149;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10144;
    wire N__10141;
    wire N__10140;
    wire N__10139;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10128;
    wire N__10127;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10110;
    wire N__10105;
    wire N__10100;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10083;
    wire N__10076;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10053;
    wire N__10042;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10018;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10002;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9979;
    wire N__9976;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9882;
    wire N__9881;
    wire N__9878;
    wire N__9877;
    wire N__9876;
    wire N__9873;
    wire N__9864;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9816;
    wire N__9813;
    wire N__9812;
    wire N__9811;
    wire N__9804;
    wire N__9801;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9736;
    wire N__9733;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9696;
    wire N__9693;
    wire N__9688;
    wire N__9681;
    wire N__9678;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9660;
    wire N__9657;
    wire N__9656;
    wire N__9653;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9635;
    wire N__9632;
    wire N__9627;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9594;
    wire N__9591;
    wire N__9590;
    wire N__9587;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9561;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9478;
    wire N__9477;
    wire N__9468;
    wire N__9465;
    wire N__9460;
    wire N__9447;
    wire N__9446;
    wire N__9445;
    wire N__9444;
    wire N__9443;
    wire N__9434;
    wire N__9433;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9429;
    wire N__9428;
    wire N__9427;
    wire N__9426;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9422;
    wire N__9415;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9388;
    wire N__9385;
    wire N__9372;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9366;
    wire N__9361;
    wire N__9354;
    wire N__9349;
    wire N__9336;
    wire N__9331;
    wire N__9328;
    wire N__9319;
    wire N__9316;
    wire N__9311;
    wire N__9292;
    wire N__9289;
    wire N__9288;
    wire N__9287;
    wire N__9286;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9277;
    wire N__9276;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9270;
    wire N__9269;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9265;
    wire N__9264;
    wire N__9263;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9259;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9251;
    wire N__9248;
    wire N__9247;
    wire N__9238;
    wire N__9229;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9213;
    wire N__9212;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9197;
    wire N__9194;
    wire N__9189;
    wire N__9184;
    wire N__9183;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9157;
    wire N__9150;
    wire N__9137;
    wire N__9134;
    wire N__9129;
    wire N__9118;
    wire N__9113;
    wire N__9110;
    wire N__9105;
    wire N__9098;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9032;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9007;
    wire N__8998;
    wire N__8997;
    wire N__8996;
    wire N__8995;
    wire N__8992;
    wire N__8991;
    wire N__8990;
    wire N__8989;
    wire N__8980;
    wire N__8977;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8958;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8943;
    wire N__8942;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8933;
    wire N__8928;
    wire N__8925;
    wire N__8918;
    wire N__8915;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8881;
    wire N__8876;
    wire N__8873;
    wire N__8872;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8864;
    wire N__8855;
    wire N__8844;
    wire N__8831;
    wire N__8822;
    wire N__8815;
    wire N__8812;
    wire N__8797;
    wire N__8796;
    wire N__8793;
    wire N__8792;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8755;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8739;
    wire N__8736;
    wire N__8735;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8719;
    wire N__8710;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8696;
    wire N__8695;
    wire N__8694;
    wire N__8693;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8688;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8668;
    wire N__8663;
    wire N__8658;
    wire N__8647;
    wire N__8642;
    wire N__8639;
    wire N__8624;
    wire N__8613;
    wire N__8610;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8573;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8567;
    wire N__8564;
    wire N__8563;
    wire N__8562;
    wire N__8561;
    wire N__8556;
    wire N__8553;
    wire N__8552;
    wire N__8549;
    wire N__8544;
    wire N__8541;
    wire N__8536;
    wire N__8533;
    wire N__8528;
    wire N__8527;
    wire N__8526;
    wire N__8523;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8510;
    wire N__8505;
    wire N__8502;
    wire N__8491;
    wire N__8486;
    wire N__8481;
    wire N__8476;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8455;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8403;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8358;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8331;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8262;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8196;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8178;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8090;
    wire N__8085;
    wire N__8082;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7974;
    wire N__7973;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7961;
    wire N__7954;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7918;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7891;
    wire N__7890;
    wire N__7885;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7872;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7853;
    wire N__7850;
    wire N__7845;
    wire N__7842;
    wire N__7837;
    wire N__7832;
    wire N__7829;
    wire N__7816;
    wire N__7815;
    wire N__7812;
    wire N__7811;
    wire N__7810;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7788;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7784;
    wire N__7779;
    wire N__7772;
    wire N__7763;
    wire N__7756;
    wire N__7755;
    wire N__7754;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7735;
    wire N__7732;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7699;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7691;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7620;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7605;
    wire N__7600;
    wire N__7597;
    wire N__7596;
    wire N__7593;
    wire N__7592;
    wire N__7589;
    wire N__7588;
    wire N__7587;
    wire N__7586;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7558;
    wire N__7555;
    wire N__7550;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7532;
    wire N__7527;
    wire N__7516;
    wire N__7515;
    wire N__7512;
    wire N__7511;
    wire N__7510;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7498;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7487;
    wire N__7486;
    wire N__7483;
    wire N__7482;
    wire N__7479;
    wire N__7472;
    wire N__7467;
    wire N__7466;
    wire N__7463;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7438;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7353;
    wire N__7350;
    wire N__7347;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7131;
    wire N__7128;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7108;
    wire N__7105;
    wire N__7104;
    wire N__7103;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7073;
    wire N__7070;
    wire N__7063;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7011;
    wire N__7010;
    wire N__7009;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6990;
    wire N__6989;
    wire N__6982;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6974;
    wire N__6963;
    wire N__6958;
    wire N__6957;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6953;
    wire N__6952;
    wire N__6941;
    wire N__6936;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6921;
    wire N__6920;
    wire N__6919;
    wire N__6914;
    wire N__6909;
    wire N__6904;
    wire N__6901;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6893;
    wire N__6888;
    wire N__6883;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6870;
    wire N__6867;
    wire N__6862;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6814;
    wire N__6813;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6771;
    wire N__6768;
    wire N__6767;
    wire N__6766;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6744;
    wire N__6741;
    wire N__6736;
    wire N__6731;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6660;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6483;
    wire N__6482;
    wire N__6481;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6463;
    wire N__6460;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6436;
    wire N__6435;
    wire N__6430;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6418;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6407;
    wire N__6406;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6392;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6368;
    wire N__6363;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6291;
    wire N__6286;
    wire N__6283;
    wire N__6282;
    wire N__6279;
    wire N__6278;
    wire N__6271;
    wire N__6268;
    wire N__6267;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6204;
    wire N__6203;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire Clock12MHz_c;
    wire \Clock50MHz.PixelClock ;
    wire GNDG0;
    wire VCCG0;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_;
    wire beamY_RNIQ8RJCCZ0Z_3_cascade_;
    wire beamY_RNIQ8RJCC_0Z0Z_3;
    wire font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9;
    wire font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_;
    wire beamY_RNI03RTE5Z0Z_4;
    wire beamY_RNI03RTE5_0Z0Z_4;
    wire font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1;
    wire Pixel_1_RNOZ0Z_34_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un68_sum_c4;
    wire beamY_RNIUAN5CR1Z0Z_3;
    wire font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i;
    wire beamY_fast_RNIEGGAZ0Z_6;
    wire font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0;
    wire font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_;
    wire beamY_RNIGBU92Z0Z_9_cascade_;
    wire beamY_RNIIDGN6_0Z0Z_7;
    wire beamY_RNIIDGN6Z0Z_7_cascade_;
    wire beamY_RNIPM0M5Z0Z_9_cascade_;
    wire beamY_RNIPM0M5_0Z0Z_9;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0;
    wire beamY_RNI1G0FH2Z0Z_3_cascade_;
    wire beamY_RNI1G0FH2_0Z0Z_3_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_;
    wire beamY_RNICCIKUQ_0Z0Z_3;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_c5;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i;
    wire font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un61_sum_c4;
    wire beamY_RNICCIKUQZ0Z_3;
    wire un4_beamylt6;
    wire un4_beamylt8_0_cascade_;
    wire un1_beamylto9_0;
    wire un1_beamylto9_3_cascade_;
    wire un5_beamx_4_cascade_;
    wire un117_pixel_6_ns_1_3_cascade_;
    wire N_192_0;
    wire N_192_0_cascade_;
    wire N_215_0;
    wire Pixel_1_RNOZ0Z_66_cascade_;
    wire un117_pixel_3_1_3;
    wire N_234_0;
    wire m3_0_cascade_;
    wire un115_pixel_2_0_5__N_9_cascade_;
    wire g0_3_1_cascade_;
    wire un115_pixel_0_a2_0_cascade_;
    wire N_281;
    wire N_231;
    wire Pixel_1_RNOZ0Z_62;
    wire N_275_0;
    wire un115_pixel_13_15__m3_a0Z0Z_0;
    wire un115_pixel_13_15__m3_a0Z0Z_0_cascade_;
    wire Pixel_1_RNOZ0Z_88;
    wire Pixel_1_RNOZ0Z_63;
    wire un115_pixel_2_0_5__N_14;
    wire bfn_4_12_0_;
    wire un4_pixel_if_generate_plus_mult1_un82_sum_cry_1;
    wire un4_pixel_if_generate_plus_mult1_un82_sum_cry_2;
    wire G_370;
    wire un4_pixel_if_generate_plus_mult1_un82_sum_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un82_sum_cry_4;
    wire un4_pixel_N_3_cascade_;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_iZ0;
    wire N_208_0_0_1;
    wire N_1260_0_0_1_cascade_;
    wire Z_decfrac2_1_0_0_0_cascade_;
    wire un115_pixel_3_0_3__N_8_0_0_0_cascade_;
    wire un117_pixel_3_1_0_1_4;
    wire m4_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1;
    wire font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_;
    wire beamY_fastZ0Z_4;
    wire beamY_fastZ0Z_9;
    wire beamY_fast_RNICEGAZ0Z_4;
    wire font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i;
    wire font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2;
    wire beamY_RNI9I1Q6Z0Z_9_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_;
    wire beamY_RNIQQREO1Z0Z_3;
    wire font_un36_pixel_if_generate_plus_mult1_un47_sum_c5;
    wire font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2;
    wire font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0;
    wire beamY_4_rep1_RNI9H1FZ0Z1;
    wire beamY_RNIHS041Z0Z_6;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0;
    wire beamY_RNIF8TM3Z0Z_9;
    wire beamY_RNIVD444Z0Z_9_cascade_;
    wire beamY_RNIGBU92Z0Z_9;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1;
    wire N_7_0_0_0_cascade_;
    wire un8_beamy_3_cascade_;
    wire Pixel_1_RNOZ0Z_43;
    wire Pixel_1_RNOZ0Z_42;
    wire N_282;
    wire font_un127_pixel_1_1_cascade_;
    wire N_336_0;
    wire un5_beamx_6;
    wire un8_beamy_3;
    wire g1_1;
    wire N_283_cascade_;
    wire N_285;
    wire font_un13_pixel_23;
    wire font_un73_pixellt7_0;
    wire font_un13_pixel_23_cascade_;
    wire Pixel_1_RNOZ0Z_60;
    wire Pixel_1_RNOZ0Z_39_cascade_;
    wire d_N_6_0;
    wire N_6;
    wire N_5_i_0;
    wire g1_0_0_cascade_;
    wire N_250_0_cascade_;
    wire N_266_0;
    wire N_242_0_cascade_;
    wire Pixel_1_RNOZ0Z_61;
    wire m3_0;
    wire Pixel_1_RNOZ0Z_69_cascade_;
    wire Pixel_1_RNOZ0Z_70;
    wire g0_35_1_cascade_;
    wire un115_pixel_13_15___m1_e_0Z0Z_1;
    wire un115_pixel_13_15__i2_mux;
    wire bfn_5_12_0_;
    wire if_generate_plus_mult1_un75_sum_cry_2_s;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire un7_pixel_1_axb1_cascade_;
    wire N_203_0_cascade_;
    wire N_268_0;
    wire g0_40_1;
    wire N_206;
    wire g0_6_1_1_cascade_;
    wire g0_6_1_cascade_;
    wire N_192_0_0;
    wire g1_3_1_cascade_;
    wire g1_3;
    wire g0_10_1_cascade_;
    wire N_309_0_cascade_;
    wire N_316_0;
    wire N_323_0_cascade_;
    wire N_302_0_0_0;
    wire N_5_0_0_0;
    wire bfn_6_3_0_;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7_c_RNIM7EZ0Z3;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire bfn_6_4_0_;
    wire un21_beamy_cry_8_c_RNIOAFZ0Z3;
    wire beamYZ0Z_3;
    wire beamYZ0Z_2;
    wire un11_visibleylto9_1;
    wire font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0;
    wire beamY_fastZ0Z_7;
    wire beamY_fastZ0Z_6;
    wire beamY_fastZ0Z_5;
    wire un11_visibleylto9_4;
    wire beamY_fast_RNI198KZ0Z_2_cascade_;
    wire font_un127_pixel_m_1;
    wire un21_beamy_cry_1_c_RNIALZ0Z73;
    wire beamY_fastZ0Z_8;
    wire beamY_fast_RNIG57DZ0Z_8;
    wire beamY_fast_RNIG57DZ0Z_8_cascade_;
    wire un5_visibley_c6_0_1;
    wire un21_beamy_cry_6_c_RNIK4DZ0Z3;
    wire un21_beamy_cry_2_c_RNICOZ0Z83;
    wire un21_beamy_cry_5_c_RNII1CZ0Z3;
    wire beamYZ0Z_4;
    wire beamY_RNI9DLCZ0Z_0;
    wire un21_beamy_cry_3_c_RNIERZ0Z93;
    wire un21_beamy_cry_4_c_RNIGUAZ0Z3;
    wire N_338_0_0_0;
    wire font_un127_pixel_m_cascade_;
    wire Pixel_c;
    wire font_un127_pixel_m_4;
    wire g0_0_1_cascade_;
    wire font_un69_pixellto3;
    wire g0_0_2;
    wire bfn_6_9_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_;
    wire Pixel_1_RNOZ0Z_82;
    wire font_un127_pixel_m_4_1_1_cascade_;
    wire font_un127_pixel_m_4_1;
    wire un7_pixel_1_c4_cascade_;
    wire font_un127_pixel_m_7_1_0;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_i;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2;
    wire N_307_0_0_1;
    wire font_un13_pixel_0_1_0_0_22_cascade_;
    wire beamY_RNIVV787O2Z0Z_2;
    wire Pixel_1_RNOZ0Z_47;
    wire N_1482_0_cascade_;
    wire bfn_6_11_0_;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_cry_1;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire un7_pixel_1_axb2_cascade_;
    wire un7_pixel_1_axb2_i;
    wire Pixel_1_RNOZ0Z_44;
    wire N_305_0_cascade_;
    wire N_326_0_0;
    wire g0_18_1;
    wire N_321_0_cascade_;
    wire N_314_0_0_0;
    wire N_328_0_0_0;
    wire g1_2_0_0_cascade_;
    wire N_192_0_1;
    wire un117_pixel_6_1_0_1_4_cascade_;
    wire N_219_0_0_1;
    wire un7_pixel_1_axb3_i;
    wire bfn_6_13_0_;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire un7_pixel_1_axb3;
    wire un7_pixel_1_axb3_cascade_;
    wire un7_pixel_1_axb1;
    wire N_532_i;
    wire un117_pixel_2_6_i3_mux;
    wire un7_pixel_1_axb2;
    wire un4_pixel_N_3;
    wire Pixel_1_RNOZ0Z_73_cascade_;
    wire Pixel_1_RNOZ0Z_72;
    wire font_un36_pixel_23;
    wire Pixel_1_RNOZ0Z_48_cascade_;
    wire N_234_0_0;
    wire d_N_3_0_0;
    wire un7_pixel_0_axb3_i;
    wire bfn_7_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum;
    wire bfn_7_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum;
    wire bfn_7_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_7;
    wire bfn_7_4_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6;
    wire Pixel_1_RNOZ0Z_18;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0;
    wire un43lto1;
    wire un43lto4_1_cascade_;
    wire un43lt10_cascade_;
    wire un1_beamY_26;
    wire un42lt10;
    wire un5_visibley_c7;
    wire bfn_7_6_0_;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_;
    wire Pixel_1_RNOZ0Z_19;
    wire un1_visiblex_27;
    wire un5_visibley_ac0_7;
    wire un5_visibley_ac0_7_cascade_;
    wire font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0;
    wire beamY_4_rep1_RNICDQEZ0_cascade_;
    wire beamY_fastZ0Z_3;
    wire un5_visibley_c2;
    wire un11_visibley;
    wire un44;
    wire Pixel_1_e_1;
    wire beamY_fastZ0Z_2;
    wire beamY_4_repZ0Z1;
    wire beamY_fast_RNIK8HHZ0Z_2;
    wire beamYZ0Z_6;
    wire beamYZ0Z_5;
    wire beamY_RNIKOP3Z0Z_7;
    wire bfn_7_8_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_i;
    wire beamYZ0Z_7;
    wire beamYZ0Z_9;
    wire un8_beamylto9_1;
    wire beamYZ0Z_8;
    wire bfn_7_9_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1;
    wire un14_visibleylt9_0;
    wire un14_visibleylt4_0;
    wire un3_beamx_5_cascade_;
    wire N_324_0_0_0;
    wire N_303_0_0_0;
    wire beamYZ0Z_0;
    wire g1_0_0_0_1;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0;
    wire g3_0_0_0_cascade_;
    wire g1_4_0_0_0;
    wire N_1869_0_0;
    wire N_1870_0_0;
    wire font_un127_pixel_6_ns_1_0_0_cascade_;
    wire font_un13_pixel_0_1_0_0_22;
    wire N_520;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i;
    wire un4_pixel_if_generate_plus_mult1_un68_sum_iZ0;
    wire beamY_RNIJ0DBZ0Z_8;
    wire VSync_c;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_iZ0;
    wire bfn_7_12_0_;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4;
    wire bfn_7_13_0_;
    wire un4_pixel_if_generate_plus_mult1_un47_sum0_2;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4;
    wire un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_;
    wire un4_pixel_if_generate_plus_mult1_un47_sum1_4;
    wire un4_pixel_if_generate_plus_mult1_un47_sum0_4;
    wire un7_pixel_0_axb4_cascade_;
    wire un4_pixel_if_generate_plus_mult1_un47_sum1_5;
    wire un4_pixel_if_generate_plus_mult1_un47_sum0_5;
    wire bfn_7_14_0_;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire un4_pixel_if_generate_plus_mult1_un54_sum_cry_1;
    wire un7_pixel_0_axb4;
    wire if_generate_plus_mult1_un47_sum_m_2;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire un4_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire un7_pixel_0_axb4_i;
    wire un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire un4_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire un4_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire un7_pixel_0_axb3;
    wire un4_pixel_if_generate_plus_mult1_un47_sum1_3;
    wire un4_pixel_if_generate_plus_mult1_un47_sum0_3;
    wire if_generate_plus_mult1_un47_sum_m_3;
    wire un1_beamY_if_generate_plus_mult1_un47_sum;
    wire bfn_8_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0;
    wire bfn_8_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un40_sum;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_0;
    wire bfn_8_4_0_;
    wire beamY_RNIALEQZ0Z_9;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2;
    wire beamY_RNIALEQ_1Z0Z_9;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_axb_6;
    wire un1_beamY_if_generate_plus_mult1_un33_sum;
    wire beamY_RNIQNF11_0Z0Z_8;
    wire beamY_i_2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0;
    wire un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4;
    wire bfn_8_6_0_;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i_8;
    wire bfn_8_7_0_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16;
    wire HSync_c;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i_8;
    wire bfn_8_8_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_i;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5;
    wire bfn_8_9_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un61_sum_i;
    wire bfn_8_10_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i;
    wire bfn_8_11_0_;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2;
    wire un5_visiblex_i_24;
    wire if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx;
    wire if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx;
    wire un5_visiblex_i_25;
    wire if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i;
    wire if_generate_plus_mult1_un47_sum_m_1;
    wire un5_visiblex_i_0_25;
    wire N_32;
    wire if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx;
    wire if_generate_plus_mult1_un47_sum_0_cry_3_ma;
    wire N_158_0_i;
    wire bfn_8_13_0_;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7;
    wire N_20_i;
    wire if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx;
    wire bfn_8_14_0_;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6;
    wire un18_beamylt4;
    wire un18_beamylto9_2_cascade_;
    wire un4_beamy_0;
    wire un18_beamylt10_0_cascade_;
    wire un8_beamy;
    wire un13_beamylt7;
    wire un15_beamy_2_cascade_;
    wire un15_beamy;
    wire un1_beamx_2_cascade_;
    wire un1_beamx;
    wire un1_beamxlt10_0;
    wire bfn_9_8_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62;
    wire font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_;
    wire font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5;
    wire font_un13_pixel_if_generate_plus_mult1_un40_sum_i;
    wire bfn_9_9_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_9_10_0_;
    wire un8_beamx_cry_9;
    wire beamXZ0Z_10;
    wire un3_beamx_7;
    wire un1_beamx_2;
    wire beamX_RNI5457Z0Z_5;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0;
    wire un3_beamx_g;
    wire font_un13_pixel_if_generate_plus_mult1_un33_sum_i;
    wire PixelClock_g;
    wire beamXZ0Z_0;
    wire bfn_9_11_0_;
    wire beamXZ0Z_1;
    wire font_un13_pixel_if_generate_plus_mult1_un75_sum;
    wire un5_visiblex_cry_0;
    wire beamXZ0Z_2;
    wire font_un13_pixel_if_generate_plus_mult1_un68_sum;
    wire un5_visiblex_cry_1;
    wire beamXZ0Z_3;
    wire un1_visiblex_24;
    wire un5_visiblex_cry_2;
    wire beamXZ0Z_4;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum;
    wire un5_visiblex_cry_3;
    wire beamXZ0Z_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum;
    wire un5_visiblex_cry_4;
    wire beamXZ0Z_6;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum;
    wire un5_visiblex_cry_5;
    wire beamXZ0Z_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire beamXZ0Z_8;
    wire bfn_9_12_0_;
    wire beamXZ0Z_9;
    wire un5_visiblex_cry_8;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_i_8;
    wire bfn_9_13_0_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum;
    wire bfn_11_12_0_;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1;
    wire CONSTANT_ONE_NET;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_1;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum;
    wire font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__6190),
            .RESETB(N__14610),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__14780),
            .DIN(N__14779),
            .DOUT(N__14778),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__14780),
            .PADOUT(N__14779),
            .PADIN(N__14778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11317),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__14771),
            .DIN(N__14770),
            .DOUT(N__14769),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__14771),
            .PADOUT(N__14770),
            .PADIN(N__14769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12366),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__14762),
            .DIN(N__14761),
            .DOUT(N__14760),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__14762),
            .PADOUT(N__14761),
            .PADIN(N__14760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8109),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__14753),
            .DIN(N__14752),
            .DOUT(N__14751),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__14753),
            .PADOUT(N__14752),
            .PADIN(N__14751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__14744),
            .DIN(N__14743),
            .DOUT(N__14742),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__14744),
            .PADOUT(N__14743),
            .PADIN(N__14742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__14735),
            .DIN(N__14734),
            .DOUT(N__14733),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__14735),
            .PADOUT(N__14734),
            .PADIN(N__14733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12373),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__14726),
            .DIN(N__14725),
            .DOUT(N__14724),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__14726),
            .PADOUT(N__14725),
            .PADIN(N__14724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8116),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__3380 (
            .O(N__14707),
            .I(N__14704));
    InMux I__3379 (
            .O(N__14704),
            .I(N__14701));
    LocalMux I__3378 (
            .O(N__14701),
            .I(N__14691));
    InMux I__3377 (
            .O(N__14700),
            .I(N__14688));
    InMux I__3376 (
            .O(N__14699),
            .I(N__14685));
    InMux I__3375 (
            .O(N__14698),
            .I(N__14682));
    InMux I__3374 (
            .O(N__14697),
            .I(N__14679));
    InMux I__3373 (
            .O(N__14696),
            .I(N__14676));
    InMux I__3372 (
            .O(N__14695),
            .I(N__14671));
    InMux I__3371 (
            .O(N__14694),
            .I(N__14671));
    Span4Mux_h I__3370 (
            .O(N__14691),
            .I(N__14666));
    LocalMux I__3369 (
            .O(N__14688),
            .I(N__14666));
    LocalMux I__3368 (
            .O(N__14685),
            .I(N__14663));
    LocalMux I__3367 (
            .O(N__14682),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    LocalMux I__3366 (
            .O(N__14679),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    LocalMux I__3365 (
            .O(N__14676),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    LocalMux I__3364 (
            .O(N__14671),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3363 (
            .O(N__14666),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3362 (
            .O(N__14663),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum));
    CascadeMux I__3361 (
            .O(N__14650),
            .I(N__14647));
    InMux I__3360 (
            .O(N__14647),
            .I(N__14644));
    LocalMux I__3359 (
            .O(N__14644),
            .I(N__14641));
    Span4Mux_h I__3358 (
            .O(N__14641),
            .I(N__14638));
    Odrv4 I__3357 (
            .O(N__14638),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0));
    InMux I__3356 (
            .O(N__14635),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1));
    InMux I__3355 (
            .O(N__14632),
            .I(N__14627));
    InMux I__3354 (
            .O(N__14631),
            .I(N__14624));
    CascadeMux I__3353 (
            .O(N__14630),
            .I(N__14620));
    LocalMux I__3352 (
            .O(N__14627),
            .I(N__14614));
    LocalMux I__3351 (
            .O(N__14624),
            .I(N__14614));
    InMux I__3350 (
            .O(N__14623),
            .I(N__14611));
    InMux I__3349 (
            .O(N__14620),
            .I(N__14601));
    InMux I__3348 (
            .O(N__14619),
            .I(N__14601));
    Span4Mux_v I__3347 (
            .O(N__14614),
            .I(N__14596));
    LocalMux I__3346 (
            .O(N__14611),
            .I(N__14596));
    IoInMux I__3345 (
            .O(N__14610),
            .I(N__14589));
    CascadeMux I__3344 (
            .O(N__14609),
            .I(N__14586));
    CascadeMux I__3343 (
            .O(N__14608),
            .I(N__14583));
    CascadeMux I__3342 (
            .O(N__14607),
            .I(N__14580));
    CascadeMux I__3341 (
            .O(N__14606),
            .I(N__14577));
    LocalMux I__3340 (
            .O(N__14601),
            .I(N__14572));
    Span4Mux_s3_h I__3339 (
            .O(N__14596),
            .I(N__14572));
    InMux I__3338 (
            .O(N__14595),
            .I(N__14569));
    InMux I__3337 (
            .O(N__14594),
            .I(N__14566));
    InMux I__3336 (
            .O(N__14593),
            .I(N__14563));
    InMux I__3335 (
            .O(N__14592),
            .I(N__14560));
    LocalMux I__3334 (
            .O(N__14589),
            .I(N__14557));
    InMux I__3333 (
            .O(N__14586),
            .I(N__14553));
    InMux I__3332 (
            .O(N__14583),
            .I(N__14550));
    InMux I__3331 (
            .O(N__14580),
            .I(N__14545));
    InMux I__3330 (
            .O(N__14577),
            .I(N__14545));
    Sp12to4 I__3329 (
            .O(N__14572),
            .I(N__14536));
    LocalMux I__3328 (
            .O(N__14569),
            .I(N__14536));
    LocalMux I__3327 (
            .O(N__14566),
            .I(N__14536));
    LocalMux I__3326 (
            .O(N__14563),
            .I(N__14536));
    LocalMux I__3325 (
            .O(N__14560),
            .I(N__14533));
    IoSpan4Mux I__3324 (
            .O(N__14557),
            .I(N__14530));
    CascadeMux I__3323 (
            .O(N__14556),
            .I(N__14527));
    LocalMux I__3322 (
            .O(N__14553),
            .I(N__14520));
    LocalMux I__3321 (
            .O(N__14550),
            .I(N__14520));
    LocalMux I__3320 (
            .O(N__14545),
            .I(N__14520));
    Span12Mux_v I__3319 (
            .O(N__14536),
            .I(N__14517));
    Span4Mux_v I__3318 (
            .O(N__14533),
            .I(N__14514));
    IoSpan4Mux I__3317 (
            .O(N__14530),
            .I(N__14511));
    InMux I__3316 (
            .O(N__14527),
            .I(N__14508));
    Span4Mux_v I__3315 (
            .O(N__14520),
            .I(N__14505));
    Odrv12 I__3314 (
            .O(N__14517),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3313 (
            .O(N__14514),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3312 (
            .O(N__14511),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3311 (
            .O(N__14508),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3310 (
            .O(N__14505),
            .I(CONSTANT_ONE_NET));
    InMux I__3309 (
            .O(N__14494),
            .I(N__14490));
    InMux I__3308 (
            .O(N__14493),
            .I(N__14487));
    LocalMux I__3307 (
            .O(N__14490),
            .I(N__14484));
    LocalMux I__3306 (
            .O(N__14487),
            .I(N__14481));
    Span4Mux_v I__3305 (
            .O(N__14484),
            .I(N__14478));
    Span4Mux_v I__3304 (
            .O(N__14481),
            .I(N__14475));
    Odrv4 I__3303 (
            .O(N__14478),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0));
    Odrv4 I__3302 (
            .O(N__14475),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0));
    InMux I__3301 (
            .O(N__14470),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__3300 (
            .O(N__14467),
            .I(N__14464));
    LocalMux I__3299 (
            .O(N__14464),
            .I(N__14461));
    Span4Mux_v I__3298 (
            .O(N__14461),
            .I(N__14458));
    Odrv4 I__3297 (
            .O(N__14458),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO));
    InMux I__3296 (
            .O(N__14455),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__3295 (
            .O(N__14452),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4));
    InMux I__3294 (
            .O(N__14449),
            .I(N__14445));
    InMux I__3293 (
            .O(N__14448),
            .I(N__14442));
    LocalMux I__3292 (
            .O(N__14445),
            .I(N__14437));
    LocalMux I__3291 (
            .O(N__14442),
            .I(N__14437));
    Span4Mux_h I__3290 (
            .O(N__14437),
            .I(N__14434));
    Odrv4 I__3289 (
            .O(N__14434),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    CascadeMux I__3288 (
            .O(N__14431),
            .I(N__14428));
    InMux I__3287 (
            .O(N__14428),
            .I(N__14425));
    LocalMux I__3286 (
            .O(N__14425),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_1));
    InMux I__3285 (
            .O(N__14422),
            .I(N__14418));
    CascadeMux I__3284 (
            .O(N__14421),
            .I(N__14415));
    LocalMux I__3283 (
            .O(N__14418),
            .I(N__14403));
    InMux I__3282 (
            .O(N__14415),
            .I(N__14400));
    CascadeMux I__3281 (
            .O(N__14414),
            .I(N__14397));
    InMux I__3280 (
            .O(N__14413),
            .I(N__14394));
    InMux I__3279 (
            .O(N__14412),
            .I(N__14391));
    InMux I__3278 (
            .O(N__14411),
            .I(N__14384));
    InMux I__3277 (
            .O(N__14410),
            .I(N__14384));
    InMux I__3276 (
            .O(N__14409),
            .I(N__14384));
    InMux I__3275 (
            .O(N__14408),
            .I(N__14377));
    InMux I__3274 (
            .O(N__14407),
            .I(N__14377));
    InMux I__3273 (
            .O(N__14406),
            .I(N__14377));
    Span4Mux_h I__3272 (
            .O(N__14403),
            .I(N__14371));
    LocalMux I__3271 (
            .O(N__14400),
            .I(N__14367));
    InMux I__3270 (
            .O(N__14397),
            .I(N__14364));
    LocalMux I__3269 (
            .O(N__14394),
            .I(N__14352));
    LocalMux I__3268 (
            .O(N__14391),
            .I(N__14347));
    LocalMux I__3267 (
            .O(N__14384),
            .I(N__14347));
    LocalMux I__3266 (
            .O(N__14377),
            .I(N__14344));
    InMux I__3265 (
            .O(N__14376),
            .I(N__14337));
    InMux I__3264 (
            .O(N__14375),
            .I(N__14337));
    InMux I__3263 (
            .O(N__14374),
            .I(N__14337));
    Span4Mux_v I__3262 (
            .O(N__14371),
            .I(N__14334));
    InMux I__3261 (
            .O(N__14370),
            .I(N__14331));
    Span4Mux_h I__3260 (
            .O(N__14367),
            .I(N__14326));
    LocalMux I__3259 (
            .O(N__14364),
            .I(N__14326));
    InMux I__3258 (
            .O(N__14363),
            .I(N__14321));
    InMux I__3257 (
            .O(N__14362),
            .I(N__14321));
    InMux I__3256 (
            .O(N__14361),
            .I(N__14316));
    InMux I__3255 (
            .O(N__14360),
            .I(N__14316));
    InMux I__3254 (
            .O(N__14359),
            .I(N__14305));
    InMux I__3253 (
            .O(N__14358),
            .I(N__14305));
    InMux I__3252 (
            .O(N__14357),
            .I(N__14305));
    InMux I__3251 (
            .O(N__14356),
            .I(N__14305));
    InMux I__3250 (
            .O(N__14355),
            .I(N__14305));
    Span4Mux_v I__3249 (
            .O(N__14352),
            .I(N__14296));
    Span4Mux_v I__3248 (
            .O(N__14347),
            .I(N__14296));
    Span4Mux_h I__3247 (
            .O(N__14344),
            .I(N__14296));
    LocalMux I__3246 (
            .O(N__14337),
            .I(N__14296));
    Odrv4 I__3245 (
            .O(N__14334),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    LocalMux I__3244 (
            .O(N__14331),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3243 (
            .O(N__14326),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    LocalMux I__3242 (
            .O(N__14321),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    LocalMux I__3241 (
            .O(N__14316),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    LocalMux I__3240 (
            .O(N__14305),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3239 (
            .O(N__14296),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum));
    CascadeMux I__3238 (
            .O(N__14281),
            .I(N__14278));
    InMux I__3237 (
            .O(N__14278),
            .I(N__14275));
    LocalMux I__3236 (
            .O(N__14275),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf));
    CascadeMux I__3235 (
            .O(N__14272),
            .I(N__14269));
    InMux I__3234 (
            .O(N__14269),
            .I(N__14266));
    LocalMux I__3233 (
            .O(N__14266),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_i));
    InMux I__3232 (
            .O(N__14263),
            .I(N__14257));
    InMux I__3231 (
            .O(N__14262),
            .I(N__14257));
    LocalMux I__3230 (
            .O(N__14257),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__3229 (
            .O(N__14254),
            .I(N__14251));
    InMux I__3228 (
            .O(N__14251),
            .I(N__14248));
    LocalMux I__3227 (
            .O(N__14248),
            .I(N__14245));
    Span4Mux_h I__3226 (
            .O(N__14245),
            .I(N__14242));
    Odrv4 I__3225 (
            .O(N__14242),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11));
    InMux I__3224 (
            .O(N__14239),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__3223 (
            .O(N__14236),
            .I(N__14233));
    InMux I__3222 (
            .O(N__14233),
            .I(N__14230));
    LocalMux I__3221 (
            .O(N__14230),
            .I(N__14227));
    Odrv4 I__3220 (
            .O(N__14227),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0));
    CascadeMux I__3219 (
            .O(N__14224),
            .I(N__14221));
    InMux I__3218 (
            .O(N__14221),
            .I(N__14218));
    LocalMux I__3217 (
            .O(N__14218),
            .I(N__14215));
    Odrv4 I__3216 (
            .O(N__14215),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1));
    InMux I__3215 (
            .O(N__14212),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5));
    CascadeMux I__3214 (
            .O(N__14209),
            .I(N__14206));
    InMux I__3213 (
            .O(N__14206),
            .I(N__14203));
    LocalMux I__3212 (
            .O(N__14203),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0));
    InMux I__3211 (
            .O(N__14200),
            .I(N__14197));
    LocalMux I__3210 (
            .O(N__14197),
            .I(N__14194));
    Odrv4 I__3209 (
            .O(N__14194),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__3208 (
            .O(N__14191),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__3207 (
            .O(N__14188),
            .I(N__14185));
    LocalMux I__3206 (
            .O(N__14185),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__3205 (
            .O(N__14182),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__3204 (
            .O(N__14179),
            .I(N__14176));
    LocalMux I__3203 (
            .O(N__14176),
            .I(N__14171));
    InMux I__3202 (
            .O(N__14175),
            .I(N__14168));
    InMux I__3201 (
            .O(N__14174),
            .I(N__14165));
    Odrv4 I__3200 (
            .O(N__14171),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1));
    LocalMux I__3199 (
            .O(N__14168),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1));
    LocalMux I__3198 (
            .O(N__14165),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1));
    CascadeMux I__3197 (
            .O(N__14158),
            .I(N__14155));
    InMux I__3196 (
            .O(N__14155),
            .I(N__14152));
    LocalMux I__3195 (
            .O(N__14152),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_i));
    InMux I__3194 (
            .O(N__14149),
            .I(N__14140));
    InMux I__3193 (
            .O(N__14148),
            .I(N__14140));
    InMux I__3192 (
            .O(N__14147),
            .I(N__14140));
    LocalMux I__3191 (
            .O(N__14140),
            .I(un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0));
    InMux I__3190 (
            .O(N__14137),
            .I(N__14131));
    InMux I__3189 (
            .O(N__14136),
            .I(N__14131));
    LocalMux I__3188 (
            .O(N__14131),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_i_8));
    InMux I__3187 (
            .O(N__14128),
            .I(N__14124));
    CascadeMux I__3186 (
            .O(N__14127),
            .I(N__14120));
    LocalMux I__3185 (
            .O(N__14124),
            .I(N__14116));
    InMux I__3184 (
            .O(N__14123),
            .I(N__14113));
    InMux I__3183 (
            .O(N__14120),
            .I(N__14110));
    InMux I__3182 (
            .O(N__14119),
            .I(N__14107));
    Span4Mux_v I__3181 (
            .O(N__14116),
            .I(N__14102));
    LocalMux I__3180 (
            .O(N__14113),
            .I(N__14102));
    LocalMux I__3179 (
            .O(N__14110),
            .I(N__14099));
    LocalMux I__3178 (
            .O(N__14107),
            .I(beamXZ0Z_2));
    Odrv4 I__3177 (
            .O(N__14102),
            .I(beamXZ0Z_2));
    Odrv4 I__3176 (
            .O(N__14099),
            .I(beamXZ0Z_2));
    InMux I__3175 (
            .O(N__14092),
            .I(N__14087));
    InMux I__3174 (
            .O(N__14091),
            .I(N__14080));
    InMux I__3173 (
            .O(N__14090),
            .I(N__14080));
    LocalMux I__3172 (
            .O(N__14087),
            .I(N__14077));
    InMux I__3171 (
            .O(N__14086),
            .I(N__14074));
    InMux I__3170 (
            .O(N__14085),
            .I(N__14071));
    LocalMux I__3169 (
            .O(N__14080),
            .I(N__14068));
    Span4Mux_h I__3168 (
            .O(N__14077),
            .I(N__14065));
    LocalMux I__3167 (
            .O(N__14074),
            .I(N__14062));
    LocalMux I__3166 (
            .O(N__14071),
            .I(N__14059));
    Span4Mux_v I__3165 (
            .O(N__14068),
            .I(N__14056));
    Span4Mux_h I__3164 (
            .O(N__14065),
            .I(N__14053));
    Span4Mux_v I__3163 (
            .O(N__14062),
            .I(N__14048));
    Span4Mux_v I__3162 (
            .O(N__14059),
            .I(N__14048));
    Odrv4 I__3161 (
            .O(N__14056),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3160 (
            .O(N__14053),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3159 (
            .O(N__14048),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum));
    InMux I__3158 (
            .O(N__14041),
            .I(un5_visiblex_cry_1));
    CascadeMux I__3157 (
            .O(N__14038),
            .I(N__14033));
    InMux I__3156 (
            .O(N__14037),
            .I(N__14029));
    CascadeMux I__3155 (
            .O(N__14036),
            .I(N__14026));
    InMux I__3154 (
            .O(N__14033),
            .I(N__14022));
    InMux I__3153 (
            .O(N__14032),
            .I(N__14019));
    LocalMux I__3152 (
            .O(N__14029),
            .I(N__14016));
    InMux I__3151 (
            .O(N__14026),
            .I(N__14013));
    InMux I__3150 (
            .O(N__14025),
            .I(N__14010));
    LocalMux I__3149 (
            .O(N__14022),
            .I(N__14007));
    LocalMux I__3148 (
            .O(N__14019),
            .I(N__14002));
    Span4Mux_h I__3147 (
            .O(N__14016),
            .I(N__14002));
    LocalMux I__3146 (
            .O(N__14013),
            .I(N__13999));
    LocalMux I__3145 (
            .O(N__14010),
            .I(beamXZ0Z_3));
    Odrv4 I__3144 (
            .O(N__14007),
            .I(beamXZ0Z_3));
    Odrv4 I__3143 (
            .O(N__14002),
            .I(beamXZ0Z_3));
    Odrv4 I__3142 (
            .O(N__13999),
            .I(beamXZ0Z_3));
    CascadeMux I__3141 (
            .O(N__13990),
            .I(N__13987));
    InMux I__3140 (
            .O(N__13987),
            .I(N__13984));
    LocalMux I__3139 (
            .O(N__13984),
            .I(N__13979));
    InMux I__3138 (
            .O(N__13983),
            .I(N__13976));
    InMux I__3137 (
            .O(N__13982),
            .I(N__13972));
    Span4Mux_v I__3136 (
            .O(N__13979),
            .I(N__13965));
    LocalMux I__3135 (
            .O(N__13976),
            .I(N__13965));
    InMux I__3134 (
            .O(N__13975),
            .I(N__13962));
    LocalMux I__3133 (
            .O(N__13972),
            .I(N__13959));
    InMux I__3132 (
            .O(N__13971),
            .I(N__13956));
    InMux I__3131 (
            .O(N__13970),
            .I(N__13953));
    Span4Mux_v I__3130 (
            .O(N__13965),
            .I(N__13950));
    LocalMux I__3129 (
            .O(N__13962),
            .I(N__13947));
    Span4Mux_h I__3128 (
            .O(N__13959),
            .I(N__13944));
    LocalMux I__3127 (
            .O(N__13956),
            .I(N__13939));
    LocalMux I__3126 (
            .O(N__13953),
            .I(N__13939));
    Odrv4 I__3125 (
            .O(N__13950),
            .I(un1_visiblex_24));
    Odrv4 I__3124 (
            .O(N__13947),
            .I(un1_visiblex_24));
    Odrv4 I__3123 (
            .O(N__13944),
            .I(un1_visiblex_24));
    Odrv4 I__3122 (
            .O(N__13939),
            .I(un1_visiblex_24));
    InMux I__3121 (
            .O(N__13930),
            .I(un5_visiblex_cry_2));
    InMux I__3120 (
            .O(N__13927),
            .I(N__13920));
    CascadeMux I__3119 (
            .O(N__13926),
            .I(N__13917));
    InMux I__3118 (
            .O(N__13925),
            .I(N__13913));
    InMux I__3117 (
            .O(N__13924),
            .I(N__13908));
    InMux I__3116 (
            .O(N__13923),
            .I(N__13908));
    LocalMux I__3115 (
            .O(N__13920),
            .I(N__13905));
    InMux I__3114 (
            .O(N__13917),
            .I(N__13902));
    InMux I__3113 (
            .O(N__13916),
            .I(N__13899));
    LocalMux I__3112 (
            .O(N__13913),
            .I(N__13892));
    LocalMux I__3111 (
            .O(N__13908),
            .I(N__13892));
    Span4Mux_h I__3110 (
            .O(N__13905),
            .I(N__13892));
    LocalMux I__3109 (
            .O(N__13902),
            .I(N__13889));
    LocalMux I__3108 (
            .O(N__13899),
            .I(beamXZ0Z_4));
    Odrv4 I__3107 (
            .O(N__13892),
            .I(beamXZ0Z_4));
    Odrv4 I__3106 (
            .O(N__13889),
            .I(beamXZ0Z_4));
    InMux I__3105 (
            .O(N__13882),
            .I(N__13876));
    InMux I__3104 (
            .O(N__13881),
            .I(N__13871));
    InMux I__3103 (
            .O(N__13880),
            .I(N__13871));
    CascadeMux I__3102 (
            .O(N__13879),
            .I(N__13865));
    LocalMux I__3101 (
            .O(N__13876),
            .I(N__13860));
    LocalMux I__3100 (
            .O(N__13871),
            .I(N__13860));
    InMux I__3099 (
            .O(N__13870),
            .I(N__13857));
    InMux I__3098 (
            .O(N__13869),
            .I(N__13853));
    InMux I__3097 (
            .O(N__13868),
            .I(N__13850));
    InMux I__3096 (
            .O(N__13865),
            .I(N__13847));
    Span4Mux_v I__3095 (
            .O(N__13860),
            .I(N__13842));
    LocalMux I__3094 (
            .O(N__13857),
            .I(N__13842));
    InMux I__3093 (
            .O(N__13856),
            .I(N__13839));
    LocalMux I__3092 (
            .O(N__13853),
            .I(N__13836));
    LocalMux I__3091 (
            .O(N__13850),
            .I(N__13833));
    LocalMux I__3090 (
            .O(N__13847),
            .I(N__13830));
    Span4Mux_v I__3089 (
            .O(N__13842),
            .I(N__13825));
    LocalMux I__3088 (
            .O(N__13839),
            .I(N__13825));
    Span4Mux_h I__3087 (
            .O(N__13836),
            .I(N__13820));
    Span4Mux_h I__3086 (
            .O(N__13833),
            .I(N__13820));
    Odrv4 I__3085 (
            .O(N__13830),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__3084 (
            .O(N__13825),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__3083 (
            .O(N__13820),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    InMux I__3082 (
            .O(N__13813),
            .I(un5_visiblex_cry_3));
    CascadeMux I__3081 (
            .O(N__13810),
            .I(N__13805));
    CascadeMux I__3080 (
            .O(N__13809),
            .I(N__13801));
    InMux I__3079 (
            .O(N__13808),
            .I(N__13796));
    InMux I__3078 (
            .O(N__13805),
            .I(N__13791));
    InMux I__3077 (
            .O(N__13804),
            .I(N__13791));
    InMux I__3076 (
            .O(N__13801),
            .I(N__13788));
    InMux I__3075 (
            .O(N__13800),
            .I(N__13785));
    InMux I__3074 (
            .O(N__13799),
            .I(N__13782));
    LocalMux I__3073 (
            .O(N__13796),
            .I(N__13777));
    LocalMux I__3072 (
            .O(N__13791),
            .I(N__13777));
    LocalMux I__3071 (
            .O(N__13788),
            .I(N__13774));
    LocalMux I__3070 (
            .O(N__13785),
            .I(beamXZ0Z_5));
    LocalMux I__3069 (
            .O(N__13782),
            .I(beamXZ0Z_5));
    Odrv4 I__3068 (
            .O(N__13777),
            .I(beamXZ0Z_5));
    Odrv4 I__3067 (
            .O(N__13774),
            .I(beamXZ0Z_5));
    InMux I__3066 (
            .O(N__13765),
            .I(N__13756));
    InMux I__3065 (
            .O(N__13764),
            .I(N__13753));
    InMux I__3064 (
            .O(N__13763),
            .I(N__13750));
    InMux I__3063 (
            .O(N__13762),
            .I(N__13747));
    InMux I__3062 (
            .O(N__13761),
            .I(N__13744));
    InMux I__3061 (
            .O(N__13760),
            .I(N__13741));
    InMux I__3060 (
            .O(N__13759),
            .I(N__13738));
    LocalMux I__3059 (
            .O(N__13756),
            .I(N__13735));
    LocalMux I__3058 (
            .O(N__13753),
            .I(N__13732));
    LocalMux I__3057 (
            .O(N__13750),
            .I(N__13729));
    LocalMux I__3056 (
            .O(N__13747),
            .I(N__13726));
    LocalMux I__3055 (
            .O(N__13744),
            .I(N__13723));
    LocalMux I__3054 (
            .O(N__13741),
            .I(N__13720));
    LocalMux I__3053 (
            .O(N__13738),
            .I(N__13717));
    Span4Mux_h I__3052 (
            .O(N__13735),
            .I(N__13710));
    Span4Mux_v I__3051 (
            .O(N__13732),
            .I(N__13710));
    Span4Mux_h I__3050 (
            .O(N__13729),
            .I(N__13710));
    Span4Mux_h I__3049 (
            .O(N__13726),
            .I(N__13703));
    Span4Mux_v I__3048 (
            .O(N__13723),
            .I(N__13703));
    Span4Mux_h I__3047 (
            .O(N__13720),
            .I(N__13703));
    Odrv4 I__3046 (
            .O(N__13717),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3045 (
            .O(N__13710),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3044 (
            .O(N__13703),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    InMux I__3043 (
            .O(N__13696),
            .I(un5_visiblex_cry_4));
    InMux I__3042 (
            .O(N__13693),
            .I(N__13690));
    LocalMux I__3041 (
            .O(N__13690),
            .I(N__13683));
    CascadeMux I__3040 (
            .O(N__13689),
            .I(N__13680));
    InMux I__3039 (
            .O(N__13688),
            .I(N__13674));
    InMux I__3038 (
            .O(N__13687),
            .I(N__13674));
    InMux I__3037 (
            .O(N__13686),
            .I(N__13671));
    Span4Mux_v I__3036 (
            .O(N__13683),
            .I(N__13668));
    InMux I__3035 (
            .O(N__13680),
            .I(N__13665));
    InMux I__3034 (
            .O(N__13679),
            .I(N__13662));
    LocalMux I__3033 (
            .O(N__13674),
            .I(N__13657));
    LocalMux I__3032 (
            .O(N__13671),
            .I(N__13657));
    Span4Mux_h I__3031 (
            .O(N__13668),
            .I(N__13654));
    LocalMux I__3030 (
            .O(N__13665),
            .I(N__13651));
    LocalMux I__3029 (
            .O(N__13662),
            .I(beamXZ0Z_6));
    Odrv4 I__3028 (
            .O(N__13657),
            .I(beamXZ0Z_6));
    Odrv4 I__3027 (
            .O(N__13654),
            .I(beamXZ0Z_6));
    Odrv4 I__3026 (
            .O(N__13651),
            .I(beamXZ0Z_6));
    InMux I__3025 (
            .O(N__13642),
            .I(N__13638));
    InMux I__3024 (
            .O(N__13641),
            .I(N__13629));
    LocalMux I__3023 (
            .O(N__13638),
            .I(N__13626));
    InMux I__3022 (
            .O(N__13637),
            .I(N__13623));
    InMux I__3021 (
            .O(N__13636),
            .I(N__13620));
    InMux I__3020 (
            .O(N__13635),
            .I(N__13617));
    InMux I__3019 (
            .O(N__13634),
            .I(N__13614));
    InMux I__3018 (
            .O(N__13633),
            .I(N__13611));
    CascadeMux I__3017 (
            .O(N__13632),
            .I(N__13608));
    LocalMux I__3016 (
            .O(N__13629),
            .I(N__13604));
    Span4Mux_h I__3015 (
            .O(N__13626),
            .I(N__13597));
    LocalMux I__3014 (
            .O(N__13623),
            .I(N__13597));
    LocalMux I__3013 (
            .O(N__13620),
            .I(N__13597));
    LocalMux I__3012 (
            .O(N__13617),
            .I(N__13594));
    LocalMux I__3011 (
            .O(N__13614),
            .I(N__13591));
    LocalMux I__3010 (
            .O(N__13611),
            .I(N__13588));
    InMux I__3009 (
            .O(N__13608),
            .I(N__13585));
    InMux I__3008 (
            .O(N__13607),
            .I(N__13582));
    Span4Mux_h I__3007 (
            .O(N__13604),
            .I(N__13579));
    Span4Mux_v I__3006 (
            .O(N__13597),
            .I(N__13572));
    Span4Mux_h I__3005 (
            .O(N__13594),
            .I(N__13572));
    Span4Mux_h I__3004 (
            .O(N__13591),
            .I(N__13572));
    Odrv12 I__3003 (
            .O(N__13588),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    LocalMux I__3002 (
            .O(N__13585),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    LocalMux I__3001 (
            .O(N__13582),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    Odrv4 I__3000 (
            .O(N__13579),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    Odrv4 I__2999 (
            .O(N__13572),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    InMux I__2998 (
            .O(N__13561),
            .I(un5_visiblex_cry_5));
    InMux I__2997 (
            .O(N__13558),
            .I(N__13547));
    InMux I__2996 (
            .O(N__13557),
            .I(N__13547));
    InMux I__2995 (
            .O(N__13556),
            .I(N__13547));
    InMux I__2994 (
            .O(N__13555),
            .I(N__13543));
    InMux I__2993 (
            .O(N__13554),
            .I(N__13540));
    LocalMux I__2992 (
            .O(N__13547),
            .I(N__13537));
    InMux I__2991 (
            .O(N__13546),
            .I(N__13534));
    LocalMux I__2990 (
            .O(N__13543),
            .I(N__13531));
    LocalMux I__2989 (
            .O(N__13540),
            .I(beamXZ0Z_7));
    Odrv4 I__2988 (
            .O(N__13537),
            .I(beamXZ0Z_7));
    LocalMux I__2987 (
            .O(N__13534),
            .I(beamXZ0Z_7));
    Odrv4 I__2986 (
            .O(N__13531),
            .I(beamXZ0Z_7));
    CascadeMux I__2985 (
            .O(N__13522),
            .I(N__13518));
    InMux I__2984 (
            .O(N__13521),
            .I(N__13515));
    InMux I__2983 (
            .O(N__13518),
            .I(N__13512));
    LocalMux I__2982 (
            .O(N__13515),
            .I(N__13507));
    LocalMux I__2981 (
            .O(N__13512),
            .I(N__13504));
    InMux I__2980 (
            .O(N__13511),
            .I(N__13496));
    InMux I__2979 (
            .O(N__13510),
            .I(N__13493));
    Span4Mux_v I__2978 (
            .O(N__13507),
            .I(N__13490));
    Span4Mux_h I__2977 (
            .O(N__13504),
            .I(N__13487));
    InMux I__2976 (
            .O(N__13503),
            .I(N__13482));
    InMux I__2975 (
            .O(N__13502),
            .I(N__13482));
    InMux I__2974 (
            .O(N__13501),
            .I(N__13479));
    InMux I__2973 (
            .O(N__13500),
            .I(N__13474));
    InMux I__2972 (
            .O(N__13499),
            .I(N__13474));
    LocalMux I__2971 (
            .O(N__13496),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__2970 (
            .O(N__13493),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    Odrv4 I__2969 (
            .O(N__13490),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    Odrv4 I__2968 (
            .O(N__13487),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__2967 (
            .O(N__13482),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__2966 (
            .O(N__13479),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__2965 (
            .O(N__13474),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    InMux I__2964 (
            .O(N__13459),
            .I(un5_visiblex_cry_6));
    CascadeMux I__2963 (
            .O(N__13456),
            .I(N__13451));
    InMux I__2962 (
            .O(N__13455),
            .I(N__13445));
    InMux I__2961 (
            .O(N__13454),
            .I(N__13445));
    InMux I__2960 (
            .O(N__13451),
            .I(N__13442));
    InMux I__2959 (
            .O(N__13450),
            .I(N__13439));
    LocalMux I__2958 (
            .O(N__13445),
            .I(N__13436));
    LocalMux I__2957 (
            .O(N__13442),
            .I(N__13433));
    LocalMux I__2956 (
            .O(N__13439),
            .I(beamXZ0Z_8));
    Odrv4 I__2955 (
            .O(N__13436),
            .I(beamXZ0Z_8));
    Odrv4 I__2954 (
            .O(N__13433),
            .I(beamXZ0Z_8));
    InMux I__2953 (
            .O(N__13426),
            .I(bfn_9_12_0_));
    CascadeMux I__2952 (
            .O(N__13423),
            .I(N__13419));
    InMux I__2951 (
            .O(N__13422),
            .I(N__13412));
    InMux I__2950 (
            .O(N__13419),
            .I(N__13412));
    InMux I__2949 (
            .O(N__13418),
            .I(N__13409));
    InMux I__2948 (
            .O(N__13417),
            .I(N__13406));
    LocalMux I__2947 (
            .O(N__13412),
            .I(N__13403));
    LocalMux I__2946 (
            .O(N__13409),
            .I(N__13400));
    LocalMux I__2945 (
            .O(N__13406),
            .I(beamXZ0Z_9));
    Odrv12 I__2944 (
            .O(N__13403),
            .I(beamXZ0Z_9));
    Odrv4 I__2943 (
            .O(N__13400),
            .I(beamXZ0Z_9));
    InMux I__2942 (
            .O(N__13393),
            .I(un5_visiblex_cry_8));
    CascadeMux I__2941 (
            .O(N__13390),
            .I(N__13385));
    InMux I__2940 (
            .O(N__13389),
            .I(N__13379));
    InMux I__2939 (
            .O(N__13388),
            .I(N__13379));
    InMux I__2938 (
            .O(N__13385),
            .I(N__13376));
    InMux I__2937 (
            .O(N__13384),
            .I(N__13373));
    LocalMux I__2936 (
            .O(N__13379),
            .I(N__13370));
    LocalMux I__2935 (
            .O(N__13376),
            .I(N__13367));
    LocalMux I__2934 (
            .O(N__13373),
            .I(beamXZ0Z_10));
    Odrv12 I__2933 (
            .O(N__13370),
            .I(beamXZ0Z_10));
    Odrv12 I__2932 (
            .O(N__13367),
            .I(beamXZ0Z_10));
    InMux I__2931 (
            .O(N__13360),
            .I(N__13357));
    LocalMux I__2930 (
            .O(N__13357),
            .I(N__13354));
    Odrv4 I__2929 (
            .O(N__13354),
            .I(un3_beamx_7));
    CascadeMux I__2928 (
            .O(N__13351),
            .I(N__13348));
    InMux I__2927 (
            .O(N__13348),
            .I(N__13344));
    InMux I__2926 (
            .O(N__13347),
            .I(N__13341));
    LocalMux I__2925 (
            .O(N__13344),
            .I(N__13338));
    LocalMux I__2924 (
            .O(N__13341),
            .I(un1_beamx_2));
    Odrv12 I__2923 (
            .O(N__13338),
            .I(un1_beamx_2));
    IoInMux I__2922 (
            .O(N__13333),
            .I(N__13330));
    LocalMux I__2921 (
            .O(N__13330),
            .I(N__13327));
    Span4Mux_s0_h I__2920 (
            .O(N__13327),
            .I(N__13324));
    Span4Mux_h I__2919 (
            .O(N__13324),
            .I(N__13321));
    Span4Mux_h I__2918 (
            .O(N__13321),
            .I(N__13318));
    Odrv4 I__2917 (
            .O(N__13318),
            .I(beamX_RNI5457Z0Z_5));
    InMux I__2916 (
            .O(N__13315),
            .I(N__13309));
    InMux I__2915 (
            .O(N__13314),
            .I(N__13309));
    LocalMux I__2914 (
            .O(N__13309),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9));
    CascadeMux I__2913 (
            .O(N__13306),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_));
    CascadeMux I__2912 (
            .O(N__13303),
            .I(N__13300));
    InMux I__2911 (
            .O(N__13300),
            .I(N__13297));
    LocalMux I__2910 (
            .O(N__13297),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0));
    InMux I__2909 (
            .O(N__13294),
            .I(N__13287));
    InMux I__2908 (
            .O(N__13293),
            .I(N__13284));
    InMux I__2907 (
            .O(N__13292),
            .I(N__13281));
    InMux I__2906 (
            .O(N__13291),
            .I(N__13276));
    InMux I__2905 (
            .O(N__13290),
            .I(N__13276));
    LocalMux I__2904 (
            .O(N__13287),
            .I(N__13267));
    LocalMux I__2903 (
            .O(N__13284),
            .I(N__13264));
    LocalMux I__2902 (
            .O(N__13281),
            .I(N__13261));
    LocalMux I__2901 (
            .O(N__13276),
            .I(N__13258));
    CEMux I__2900 (
            .O(N__13275),
            .I(N__13237));
    CEMux I__2899 (
            .O(N__13274),
            .I(N__13237));
    CEMux I__2898 (
            .O(N__13273),
            .I(N__13237));
    CEMux I__2897 (
            .O(N__13272),
            .I(N__13237));
    CEMux I__2896 (
            .O(N__13271),
            .I(N__13237));
    CEMux I__2895 (
            .O(N__13270),
            .I(N__13237));
    Glb2LocalMux I__2894 (
            .O(N__13267),
            .I(N__13237));
    Glb2LocalMux I__2893 (
            .O(N__13264),
            .I(N__13237));
    Glb2LocalMux I__2892 (
            .O(N__13261),
            .I(N__13237));
    Glb2LocalMux I__2891 (
            .O(N__13258),
            .I(N__13237));
    GlobalMux I__2890 (
            .O(N__13237),
            .I(N__13234));
    gio2CtrlBuf I__2889 (
            .O(N__13234),
            .I(un3_beamx_g));
    InMux I__2888 (
            .O(N__13231),
            .I(N__13228));
    LocalMux I__2887 (
            .O(N__13228),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_i));
    ClkMux I__2886 (
            .O(N__13225),
            .I(N__13186));
    ClkMux I__2885 (
            .O(N__13224),
            .I(N__13186));
    ClkMux I__2884 (
            .O(N__13223),
            .I(N__13186));
    ClkMux I__2883 (
            .O(N__13222),
            .I(N__13186));
    ClkMux I__2882 (
            .O(N__13221),
            .I(N__13186));
    ClkMux I__2881 (
            .O(N__13220),
            .I(N__13186));
    ClkMux I__2880 (
            .O(N__13219),
            .I(N__13186));
    ClkMux I__2879 (
            .O(N__13218),
            .I(N__13186));
    ClkMux I__2878 (
            .O(N__13217),
            .I(N__13186));
    ClkMux I__2877 (
            .O(N__13216),
            .I(N__13186));
    ClkMux I__2876 (
            .O(N__13215),
            .I(N__13186));
    ClkMux I__2875 (
            .O(N__13214),
            .I(N__13186));
    ClkMux I__2874 (
            .O(N__13213),
            .I(N__13186));
    GlobalMux I__2873 (
            .O(N__13186),
            .I(N__13183));
    gio2CtrlBuf I__2872 (
            .O(N__13183),
            .I(PixelClock_g));
    InMux I__2871 (
            .O(N__13180),
            .I(N__13175));
    InMux I__2870 (
            .O(N__13179),
            .I(N__13172));
    InMux I__2869 (
            .O(N__13178),
            .I(N__13169));
    LocalMux I__2868 (
            .O(N__13175),
            .I(N__13161));
    LocalMux I__2867 (
            .O(N__13172),
            .I(N__13156));
    LocalMux I__2866 (
            .O(N__13169),
            .I(N__13156));
    InMux I__2865 (
            .O(N__13168),
            .I(N__13153));
    CascadeMux I__2864 (
            .O(N__13167),
            .I(N__13150));
    InMux I__2863 (
            .O(N__13166),
            .I(N__13145));
    InMux I__2862 (
            .O(N__13165),
            .I(N__13145));
    InMux I__2861 (
            .O(N__13164),
            .I(N__13142));
    Span4Mux_h I__2860 (
            .O(N__13161),
            .I(N__13139));
    Span4Mux_v I__2859 (
            .O(N__13156),
            .I(N__13134));
    LocalMux I__2858 (
            .O(N__13153),
            .I(N__13134));
    InMux I__2857 (
            .O(N__13150),
            .I(N__13131));
    LocalMux I__2856 (
            .O(N__13145),
            .I(beamXZ0Z_0));
    LocalMux I__2855 (
            .O(N__13142),
            .I(beamXZ0Z_0));
    Odrv4 I__2854 (
            .O(N__13139),
            .I(beamXZ0Z_0));
    Odrv4 I__2853 (
            .O(N__13134),
            .I(beamXZ0Z_0));
    LocalMux I__2852 (
            .O(N__13131),
            .I(beamXZ0Z_0));
    InMux I__2851 (
            .O(N__13120),
            .I(N__13115));
    CascadeMux I__2850 (
            .O(N__13119),
            .I(N__13110));
    InMux I__2849 (
            .O(N__13118),
            .I(N__13107));
    LocalMux I__2848 (
            .O(N__13115),
            .I(N__13104));
    CascadeMux I__2847 (
            .O(N__13114),
            .I(N__13101));
    InMux I__2846 (
            .O(N__13113),
            .I(N__13098));
    InMux I__2845 (
            .O(N__13110),
            .I(N__13095));
    LocalMux I__2844 (
            .O(N__13107),
            .I(N__13092));
    Span4Mux_h I__2843 (
            .O(N__13104),
            .I(N__13089));
    InMux I__2842 (
            .O(N__13101),
            .I(N__13086));
    LocalMux I__2841 (
            .O(N__13098),
            .I(beamXZ0Z_1));
    LocalMux I__2840 (
            .O(N__13095),
            .I(beamXZ0Z_1));
    Odrv4 I__2839 (
            .O(N__13092),
            .I(beamXZ0Z_1));
    Odrv4 I__2838 (
            .O(N__13089),
            .I(beamXZ0Z_1));
    LocalMux I__2837 (
            .O(N__13086),
            .I(beamXZ0Z_1));
    InMux I__2836 (
            .O(N__13075),
            .I(N__13061));
    InMux I__2835 (
            .O(N__13074),
            .I(N__13061));
    InMux I__2834 (
            .O(N__13073),
            .I(N__13058));
    InMux I__2833 (
            .O(N__13072),
            .I(N__13052));
    InMux I__2832 (
            .O(N__13071),
            .I(N__13052));
    InMux I__2831 (
            .O(N__13070),
            .I(N__13049));
    InMux I__2830 (
            .O(N__13069),
            .I(N__13040));
    InMux I__2829 (
            .O(N__13068),
            .I(N__13040));
    InMux I__2828 (
            .O(N__13067),
            .I(N__13040));
    InMux I__2827 (
            .O(N__13066),
            .I(N__13040));
    LocalMux I__2826 (
            .O(N__13061),
            .I(N__13037));
    LocalMux I__2825 (
            .O(N__13058),
            .I(N__13034));
    InMux I__2824 (
            .O(N__13057),
            .I(N__13031));
    LocalMux I__2823 (
            .O(N__13052),
            .I(N__13024));
    LocalMux I__2822 (
            .O(N__13049),
            .I(N__13024));
    LocalMux I__2821 (
            .O(N__13040),
            .I(N__13024));
    Span4Mux_v I__2820 (
            .O(N__13037),
            .I(N__13019));
    Span4Mux_v I__2819 (
            .O(N__13034),
            .I(N__13019));
    LocalMux I__2818 (
            .O(N__13031),
            .I(N__13016));
    Span4Mux_h I__2817 (
            .O(N__13024),
            .I(N__13013));
    Sp12to4 I__2816 (
            .O(N__13019),
            .I(N__13008));
    Span12Mux_s5_v I__2815 (
            .O(N__13016),
            .I(N__13008));
    Odrv4 I__2814 (
            .O(N__13013),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum));
    Odrv12 I__2813 (
            .O(N__13008),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum));
    InMux I__2812 (
            .O(N__13003),
            .I(un5_visiblex_cry_0));
    InMux I__2811 (
            .O(N__13000),
            .I(un8_beamx_cry_1));
    InMux I__2810 (
            .O(N__12997),
            .I(un8_beamx_cry_2));
    InMux I__2809 (
            .O(N__12994),
            .I(un8_beamx_cry_3));
    InMux I__2808 (
            .O(N__12991),
            .I(un8_beamx_cry_4));
    InMux I__2807 (
            .O(N__12988),
            .I(un8_beamx_cry_5));
    InMux I__2806 (
            .O(N__12985),
            .I(un8_beamx_cry_6));
    InMux I__2805 (
            .O(N__12982),
            .I(un8_beamx_cry_7));
    InMux I__2804 (
            .O(N__12979),
            .I(bfn_9_10_0_));
    InMux I__2803 (
            .O(N__12976),
            .I(un8_beamx_cry_9));
    CascadeMux I__2802 (
            .O(N__12973),
            .I(N__12970));
    InMux I__2801 (
            .O(N__12970),
            .I(N__12967));
    LocalMux I__2800 (
            .O(N__12967),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63));
    InMux I__2799 (
            .O(N__12964),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1));
    CascadeMux I__2798 (
            .O(N__12961),
            .I(N__12958));
    InMux I__2797 (
            .O(N__12958),
            .I(N__12955));
    LocalMux I__2796 (
            .O(N__12955),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1));
    InMux I__2795 (
            .O(N__12952),
            .I(N__12949));
    LocalMux I__2794 (
            .O(N__12949),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4));
    InMux I__2793 (
            .O(N__12946),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__2792 (
            .O(N__12943),
            .I(N__12940));
    LocalMux I__2791 (
            .O(N__12940),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62));
    InMux I__2790 (
            .O(N__12937),
            .I(N__12934));
    LocalMux I__2789 (
            .O(N__12934),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__2788 (
            .O(N__12931),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__2787 (
            .O(N__12928),
            .I(N__12925));
    LocalMux I__2786 (
            .O(N__12925),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__2785 (
            .O(N__12922),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__2784 (
            .O(N__12919),
            .I(N__12915));
    InMux I__2783 (
            .O(N__12918),
            .I(N__12912));
    LocalMux I__2782 (
            .O(N__12915),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5));
    LocalMux I__2781 (
            .O(N__12912),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5));
    CascadeMux I__2780 (
            .O(N__12907),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_));
    CascadeMux I__2779 (
            .O(N__12904),
            .I(N__12900));
    CascadeMux I__2778 (
            .O(N__12903),
            .I(N__12897));
    InMux I__2777 (
            .O(N__12900),
            .I(N__12892));
    InMux I__2776 (
            .O(N__12897),
            .I(N__12892));
    LocalMux I__2775 (
            .O(N__12892),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__2774 (
            .O(N__12889),
            .I(N__12884));
    InMux I__2773 (
            .O(N__12888),
            .I(N__12879));
    InMux I__2772 (
            .O(N__12887),
            .I(N__12879));
    LocalMux I__2771 (
            .O(N__12884),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2));
    LocalMux I__2770 (
            .O(N__12879),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2));
    CascadeMux I__2769 (
            .O(N__12874),
            .I(N__12870));
    CascadeMux I__2768 (
            .O(N__12873),
            .I(N__12867));
    InMux I__2767 (
            .O(N__12870),
            .I(N__12862));
    InMux I__2766 (
            .O(N__12867),
            .I(N__12862));
    LocalMux I__2765 (
            .O(N__12862),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5));
    InMux I__2764 (
            .O(N__12859),
            .I(N__12856));
    LocalMux I__2763 (
            .O(N__12856),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_i));
    InMux I__2762 (
            .O(N__12853),
            .I(N__12850));
    LocalMux I__2761 (
            .O(N__12850),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO));
    InMux I__2760 (
            .O(N__12847),
            .I(un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6));
    CascadeMux I__2759 (
            .O(N__12844),
            .I(N__12841));
    InMux I__2758 (
            .O(N__12841),
            .I(N__12837));
    InMux I__2757 (
            .O(N__12840),
            .I(N__12834));
    LocalMux I__2756 (
            .O(N__12837),
            .I(N__12829));
    LocalMux I__2755 (
            .O(N__12834),
            .I(N__12829));
    Span4Mux_h I__2754 (
            .O(N__12829),
            .I(N__12826));
    Odrv4 I__2753 (
            .O(N__12826),
            .I(un18_beamylt4));
    CascadeMux I__2752 (
            .O(N__12823),
            .I(un18_beamylto9_2_cascade_));
    InMux I__2751 (
            .O(N__12820),
            .I(N__12817));
    LocalMux I__2750 (
            .O(N__12817),
            .I(N__12814));
    Odrv12 I__2749 (
            .O(N__12814),
            .I(un4_beamy_0));
    CascadeMux I__2748 (
            .O(N__12811),
            .I(un18_beamylt10_0_cascade_));
    InMux I__2747 (
            .O(N__12808),
            .I(N__12805));
    LocalMux I__2746 (
            .O(N__12805),
            .I(N__12802));
    Span4Mux_h I__2745 (
            .O(N__12802),
            .I(N__12799));
    Odrv4 I__2744 (
            .O(N__12799),
            .I(un8_beamy));
    InMux I__2743 (
            .O(N__12796),
            .I(N__12793));
    LocalMux I__2742 (
            .O(N__12793),
            .I(un13_beamylt7));
    CascadeMux I__2741 (
            .O(N__12790),
            .I(un15_beamy_2_cascade_));
    InMux I__2740 (
            .O(N__12787),
            .I(N__12784));
    LocalMux I__2739 (
            .O(N__12784),
            .I(N__12780));
    InMux I__2738 (
            .O(N__12783),
            .I(N__12777));
    Span4Mux_v I__2737 (
            .O(N__12780),
            .I(N__12774));
    LocalMux I__2736 (
            .O(N__12777),
            .I(N__12771));
    Odrv4 I__2735 (
            .O(N__12774),
            .I(un15_beamy));
    Odrv12 I__2734 (
            .O(N__12771),
            .I(un15_beamy));
    CascadeMux I__2733 (
            .O(N__12766),
            .I(un1_beamx_2_cascade_));
    InMux I__2732 (
            .O(N__12763),
            .I(N__12759));
    InMux I__2731 (
            .O(N__12762),
            .I(N__12756));
    LocalMux I__2730 (
            .O(N__12759),
            .I(N__12751));
    LocalMux I__2729 (
            .O(N__12756),
            .I(N__12751));
    Odrv12 I__2728 (
            .O(N__12751),
            .I(un1_beamx));
    InMux I__2727 (
            .O(N__12748),
            .I(N__12745));
    LocalMux I__2726 (
            .O(N__12745),
            .I(un1_beamxlt10_0));
    InMux I__2725 (
            .O(N__12742),
            .I(N__12739));
    LocalMux I__2724 (
            .O(N__12739),
            .I(N__12734));
    InMux I__2723 (
            .O(N__12738),
            .I(N__12729));
    InMux I__2722 (
            .O(N__12737),
            .I(N__12729));
    Odrv12 I__2721 (
            .O(N__12734),
            .I(N_32));
    LocalMux I__2720 (
            .O(N__12729),
            .I(N_32));
    InMux I__2719 (
            .O(N__12724),
            .I(N__12721));
    LocalMux I__2718 (
            .O(N__12721),
            .I(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx));
    CascadeMux I__2717 (
            .O(N__12718),
            .I(N__12715));
    InMux I__2716 (
            .O(N__12715),
            .I(N__12712));
    LocalMux I__2715 (
            .O(N__12712),
            .I(if_generate_plus_mult1_un47_sum_0_cry_3_ma));
    InMux I__2714 (
            .O(N__12709),
            .I(N__12706));
    LocalMux I__2713 (
            .O(N__12706),
            .I(N_158_0_i));
    InMux I__2712 (
            .O(N__12703),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__2711 (
            .O(N__12700),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__2710 (
            .O(N__12697),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__2709 (
            .O(N__12694),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7));
    InMux I__2708 (
            .O(N__12691),
            .I(N__12687));
    InMux I__2707 (
            .O(N__12690),
            .I(N__12683));
    LocalMux I__2706 (
            .O(N__12687),
            .I(N__12680));
    InMux I__2705 (
            .O(N__12686),
            .I(N__12674));
    LocalMux I__2704 (
            .O(N__12683),
            .I(N__12669));
    Span4Mux_v I__2703 (
            .O(N__12680),
            .I(N__12669));
    InMux I__2702 (
            .O(N__12679),
            .I(N__12666));
    CascadeMux I__2701 (
            .O(N__12678),
            .I(N__12663));
    CascadeMux I__2700 (
            .O(N__12677),
            .I(N__12658));
    LocalMux I__2699 (
            .O(N__12674),
            .I(N__12653));
    Span4Mux_v I__2698 (
            .O(N__12669),
            .I(N__12650));
    LocalMux I__2697 (
            .O(N__12666),
            .I(N__12647));
    InMux I__2696 (
            .O(N__12663),
            .I(N__12642));
    InMux I__2695 (
            .O(N__12662),
            .I(N__12642));
    InMux I__2694 (
            .O(N__12661),
            .I(N__12637));
    InMux I__2693 (
            .O(N__12658),
            .I(N__12637));
    InMux I__2692 (
            .O(N__12657),
            .I(N__12632));
    InMux I__2691 (
            .O(N__12656),
            .I(N__12632));
    Odrv4 I__2690 (
            .O(N__12653),
            .I(N_20_i));
    Odrv4 I__2689 (
            .O(N__12650),
            .I(N_20_i));
    Odrv4 I__2688 (
            .O(N__12647),
            .I(N_20_i));
    LocalMux I__2687 (
            .O(N__12642),
            .I(N_20_i));
    LocalMux I__2686 (
            .O(N__12637),
            .I(N_20_i));
    LocalMux I__2685 (
            .O(N__12632),
            .I(N_20_i));
    CascadeMux I__2684 (
            .O(N__12619),
            .I(N__12616));
    InMux I__2683 (
            .O(N__12616),
            .I(N__12613));
    LocalMux I__2682 (
            .O(N__12613),
            .I(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx));
    InMux I__2681 (
            .O(N__12610),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__2680 (
            .O(N__12607),
            .I(N__12603));
    InMux I__2679 (
            .O(N__12606),
            .I(N__12600));
    LocalMux I__2678 (
            .O(N__12603),
            .I(N__12594));
    LocalMux I__2677 (
            .O(N__12600),
            .I(N__12594));
    InMux I__2676 (
            .O(N__12599),
            .I(N__12591));
    Span4Mux_h I__2675 (
            .O(N__12594),
            .I(N__12588));
    LocalMux I__2674 (
            .O(N__12591),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2));
    Odrv4 I__2673 (
            .O(N__12588),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2));
    CascadeMux I__2672 (
            .O(N__12583),
            .I(N__12580));
    InMux I__2671 (
            .O(N__12580),
            .I(N__12577));
    LocalMux I__2670 (
            .O(N__12577),
            .I(un5_visiblex_i_24));
    CascadeMux I__2669 (
            .O(N__12574),
            .I(N__12571));
    InMux I__2668 (
            .O(N__12571),
            .I(N__12568));
    LocalMux I__2667 (
            .O(N__12568),
            .I(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx));
    InMux I__2666 (
            .O(N__12565),
            .I(N__12562));
    LocalMux I__2665 (
            .O(N__12562),
            .I(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx));
    CascadeMux I__2664 (
            .O(N__12559),
            .I(N__12556));
    InMux I__2663 (
            .O(N__12556),
            .I(N__12553));
    LocalMux I__2662 (
            .O(N__12553),
            .I(un5_visiblex_i_25));
    InMux I__2661 (
            .O(N__12550),
            .I(N__12547));
    LocalMux I__2660 (
            .O(N__12547),
            .I(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx));
    CascadeMux I__2659 (
            .O(N__12544),
            .I(N__12541));
    InMux I__2658 (
            .O(N__12541),
            .I(N__12538));
    LocalMux I__2657 (
            .O(N__12538),
            .I(font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i));
    InMux I__2656 (
            .O(N__12535),
            .I(N__12532));
    LocalMux I__2655 (
            .O(N__12532),
            .I(N__12529));
    Span4Mux_h I__2654 (
            .O(N__12529),
            .I(N__12526));
    Odrv4 I__2653 (
            .O(N__12526),
            .I(if_generate_plus_mult1_un47_sum_m_1));
    CascadeMux I__2652 (
            .O(N__12523),
            .I(N__12520));
    InMux I__2651 (
            .O(N__12520),
            .I(N__12517));
    LocalMux I__2650 (
            .O(N__12517),
            .I(un5_visiblex_i_0_25));
    InMux I__2649 (
            .O(N__12514),
            .I(N__12511));
    LocalMux I__2648 (
            .O(N__12511),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__2647 (
            .O(N__12508),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__2646 (
            .O(N__12505),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4));
    InMux I__2645 (
            .O(N__12502),
            .I(N__12498));
    InMux I__2644 (
            .O(N__12501),
            .I(N__12495));
    LocalMux I__2643 (
            .O(N__12498),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251));
    LocalMux I__2642 (
            .O(N__12495),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251));
    CascadeMux I__2641 (
            .O(N__12490),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_));
    CascadeMux I__2640 (
            .O(N__12487),
            .I(N__12483));
    CascadeMux I__2639 (
            .O(N__12486),
            .I(N__12480));
    InMux I__2638 (
            .O(N__12483),
            .I(N__12475));
    InMux I__2637 (
            .O(N__12480),
            .I(N__12475));
    LocalMux I__2636 (
            .O(N__12475),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5));
    CascadeMux I__2635 (
            .O(N__12472),
            .I(N__12469));
    InMux I__2634 (
            .O(N__12469),
            .I(N__12466));
    LocalMux I__2633 (
            .O(N__12466),
            .I(N__12463));
    Odrv12 I__2632 (
            .O(N__12463),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__2631 (
            .O(N__12460),
            .I(N__12457));
    InMux I__2630 (
            .O(N__12457),
            .I(N__12454));
    LocalMux I__2629 (
            .O(N__12454),
            .I(N__12451));
    Span4Mux_h I__2628 (
            .O(N__12451),
            .I(N__12448));
    Odrv4 I__2627 (
            .O(N__12448),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1));
    InMux I__2626 (
            .O(N__12445),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__2625 (
            .O(N__12442),
            .I(N__12439));
    InMux I__2624 (
            .O(N__12439),
            .I(N__12436));
    LocalMux I__2623 (
            .O(N__12436),
            .I(N__12433));
    Odrv12 I__2622 (
            .O(N__12433),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2));
    InMux I__2621 (
            .O(N__12430),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__2620 (
            .O(N__12427),
            .I(N__12424));
    LocalMux I__2619 (
            .O(N__12424),
            .I(N__12421));
    Odrv12 I__2618 (
            .O(N__12421),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__2617 (
            .O(N__12418),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__2616 (
            .O(N__12415),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1));
    InMux I__2615 (
            .O(N__12412),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__2614 (
            .O(N__12409),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__2613 (
            .O(N__12406),
            .I(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__2612 (
            .O(N__12403),
            .I(N__12400));
    LocalMux I__2611 (
            .O(N__12400),
            .I(N__12397));
    Odrv4 I__2610 (
            .O(N__12397),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_i));
    CascadeMux I__2609 (
            .O(N__12394),
            .I(N__12391));
    InMux I__2608 (
            .O(N__12391),
            .I(N__12388));
    LocalMux I__2607 (
            .O(N__12388),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0));
    InMux I__2606 (
            .O(N__12385),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1));
    InMux I__2605 (
            .O(N__12382),
            .I(N__12379));
    LocalMux I__2604 (
            .O(N__12379),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41));
    InMux I__2603 (
            .O(N__12376),
            .I(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    IoInMux I__2602 (
            .O(N__12373),
            .I(N__12370));
    LocalMux I__2601 (
            .O(N__12370),
            .I(N__12367));
    Span4Mux_s2_v I__2600 (
            .O(N__12367),
            .I(N__12363));
    IoInMux I__2599 (
            .O(N__12366),
            .I(N__12360));
    Span4Mux_h I__2598 (
            .O(N__12363),
            .I(N__12357));
    LocalMux I__2597 (
            .O(N__12360),
            .I(N__12354));
    Span4Mux_v I__2596 (
            .O(N__12357),
            .I(N__12351));
    Span4Mux_s3_v I__2595 (
            .O(N__12354),
            .I(N__12348));
    Odrv4 I__2594 (
            .O(N__12351),
            .I(HSync_c));
    Odrv4 I__2593 (
            .O(N__12348),
            .I(HSync_c));
    InMux I__2592 (
            .O(N__12343),
            .I(N__12337));
    InMux I__2591 (
            .O(N__12342),
            .I(N__12337));
    LocalMux I__2590 (
            .O(N__12337),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__2589 (
            .O(N__12334),
            .I(N__12331));
    InMux I__2588 (
            .O(N__12331),
            .I(N__12328));
    LocalMux I__2587 (
            .O(N__12328),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156));
    InMux I__2586 (
            .O(N__12325),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__2585 (
            .O(N__12322),
            .I(N__12319));
    LocalMux I__2584 (
            .O(N__12319),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99));
    InMux I__2583 (
            .O(N__12316),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__2582 (
            .O(N__12313),
            .I(N__12310));
    LocalMux I__2581 (
            .O(N__12310),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__2580 (
            .O(N__12307),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2579 (
            .O(N__12304),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2578 (
            .O(N__12301),
            .I(N__12298));
    LocalMux I__2577 (
            .O(N__12298),
            .I(font_un13_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__2576 (
            .O(N__12295),
            .I(N__12290));
    InMux I__2575 (
            .O(N__12294),
            .I(N__12287));
    InMux I__2574 (
            .O(N__12293),
            .I(N__12284));
    LocalMux I__2573 (
            .O(N__12290),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0));
    LocalMux I__2572 (
            .O(N__12287),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0));
    LocalMux I__2571 (
            .O(N__12284),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0));
    CascadeMux I__2570 (
            .O(N__12277),
            .I(N__12273));
    CascadeMux I__2569 (
            .O(N__12276),
            .I(N__12270));
    InMux I__2568 (
            .O(N__12273),
            .I(N__12265));
    InMux I__2567 (
            .O(N__12270),
            .I(N__12265));
    LocalMux I__2566 (
            .O(N__12265),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__2565 (
            .O(N__12262),
            .I(N__12259));
    LocalMux I__2564 (
            .O(N__12259),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0));
    CascadeMux I__2563 (
            .O(N__12256),
            .I(N__12253));
    InMux I__2562 (
            .O(N__12253),
            .I(N__12250));
    LocalMux I__2561 (
            .O(N__12250),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i));
    InMux I__2560 (
            .O(N__12247),
            .I(N__12244));
    LocalMux I__2559 (
            .O(N__12244),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__2558 (
            .O(N__12241),
            .I(N__12238));
    LocalMux I__2557 (
            .O(N__12238),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983));
    InMux I__2556 (
            .O(N__12235),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2555 (
            .O(N__12232),
            .I(N__12228));
    InMux I__2554 (
            .O(N__12231),
            .I(N__12223));
    InMux I__2553 (
            .O(N__12228),
            .I(N__12223));
    LocalMux I__2552 (
            .O(N__12223),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4));
    InMux I__2551 (
            .O(N__12220),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__2550 (
            .O(N__12217),
            .I(N__12214));
    LocalMux I__2549 (
            .O(N__12214),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__2548 (
            .O(N__12211),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__2547 (
            .O(N__12208),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__2546 (
            .O(N__12205),
            .I(N__12201));
    InMux I__2545 (
            .O(N__12204),
            .I(N__12196));
    InMux I__2544 (
            .O(N__12201),
            .I(N__12189));
    InMux I__2543 (
            .O(N__12200),
            .I(N__12189));
    InMux I__2542 (
            .O(N__12199),
            .I(N__12189));
    LocalMux I__2541 (
            .O(N__12196),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16));
    LocalMux I__2540 (
            .O(N__12189),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16));
    InMux I__2539 (
            .O(N__12184),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__2538 (
            .O(N__12181),
            .I(N__12178));
    LocalMux I__2537 (
            .O(N__12178),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    CascadeMux I__2536 (
            .O(N__12175),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    CascadeMux I__2535 (
            .O(N__12172),
            .I(N__12169));
    InMux I__2534 (
            .O(N__12169),
            .I(N__12165));
    InMux I__2533 (
            .O(N__12168),
            .I(N__12161));
    LocalMux I__2532 (
            .O(N__12165),
            .I(N__12158));
    InMux I__2531 (
            .O(N__12164),
            .I(N__12155));
    LocalMux I__2530 (
            .O(N__12161),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    Odrv4 I__2529 (
            .O(N__12158),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__2528 (
            .O(N__12155),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    InMux I__2527 (
            .O(N__12148),
            .I(N__12139));
    InMux I__2526 (
            .O(N__12147),
            .I(N__12139));
    InMux I__2525 (
            .O(N__12146),
            .I(N__12136));
    InMux I__2524 (
            .O(N__12145),
            .I(N__12126));
    InMux I__2523 (
            .O(N__12144),
            .I(N__12126));
    LocalMux I__2522 (
            .O(N__12139),
            .I(N__12123));
    LocalMux I__2521 (
            .O(N__12136),
            .I(N__12120));
    InMux I__2520 (
            .O(N__12135),
            .I(N__12115));
    InMux I__2519 (
            .O(N__12134),
            .I(N__12115));
    InMux I__2518 (
            .O(N__12133),
            .I(N__12112));
    InMux I__2517 (
            .O(N__12132),
            .I(N__12107));
    InMux I__2516 (
            .O(N__12131),
            .I(N__12107));
    LocalMux I__2515 (
            .O(N__12126),
            .I(N__12102));
    Span4Mux_v I__2514 (
            .O(N__12123),
            .I(N__12102));
    Odrv4 I__2513 (
            .O(N__12120),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__2512 (
            .O(N__12115),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__2511 (
            .O(N__12112),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__2510 (
            .O(N__12107),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2509 (
            .O(N__12102),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    InMux I__2508 (
            .O(N__12091),
            .I(N__12088));
    LocalMux I__2507 (
            .O(N__12088),
            .I(beamY_RNIQNF11_0Z0Z_8));
    InMux I__2506 (
            .O(N__12085),
            .I(N__12081));
    CascadeMux I__2505 (
            .O(N__12084),
            .I(N__12076));
    LocalMux I__2504 (
            .O(N__12081),
            .I(N__12073));
    InMux I__2503 (
            .O(N__12080),
            .I(N__12069));
    InMux I__2502 (
            .O(N__12079),
            .I(N__12064));
    InMux I__2501 (
            .O(N__12076),
            .I(N__12064));
    Span4Mux_h I__2500 (
            .O(N__12073),
            .I(N__12061));
    InMux I__2499 (
            .O(N__12072),
            .I(N__12058));
    LocalMux I__2498 (
            .O(N__12069),
            .I(beamY_i_2));
    LocalMux I__2497 (
            .O(N__12064),
            .I(beamY_i_2));
    Odrv4 I__2496 (
            .O(N__12061),
            .I(beamY_i_2));
    LocalMux I__2495 (
            .O(N__12058),
            .I(beamY_i_2));
    InMux I__2494 (
            .O(N__12049),
            .I(N__12045));
    InMux I__2493 (
            .O(N__12048),
            .I(N__12042));
    LocalMux I__2492 (
            .O(N__12045),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0));
    LocalMux I__2491 (
            .O(N__12042),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0));
    InMux I__2490 (
            .O(N__12037),
            .I(N__12034));
    LocalMux I__2489 (
            .O(N__12034),
            .I(un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4));
    InMux I__2488 (
            .O(N__12031),
            .I(N__12028));
    LocalMux I__2487 (
            .O(N__12028),
            .I(N__12025));
    Odrv4 I__2486 (
            .O(N__12025),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6));
    InMux I__2485 (
            .O(N__12022),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__2484 (
            .O(N__12019),
            .I(N__12016));
    InMux I__2483 (
            .O(N__12016),
            .I(N__12013));
    LocalMux I__2482 (
            .O(N__12013),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9));
    InMux I__2481 (
            .O(N__12010),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__2480 (
            .O(N__12007),
            .I(N__12004));
    LocalMux I__2479 (
            .O(N__12004),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__2478 (
            .O(N__12001),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__2477 (
            .O(N__11998),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__2476 (
            .O(N__11995),
            .I(N__11991));
    InMux I__2475 (
            .O(N__11994),
            .I(N__11987));
    InMux I__2474 (
            .O(N__11991),
            .I(N__11982));
    InMux I__2473 (
            .O(N__11990),
            .I(N__11982));
    LocalMux I__2472 (
            .O(N__11987),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0));
    LocalMux I__2471 (
            .O(N__11982),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0));
    CascadeMux I__2470 (
            .O(N__11977),
            .I(N__11974));
    InMux I__2469 (
            .O(N__11974),
            .I(N__11971));
    LocalMux I__2468 (
            .O(N__11971),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51));
    InMux I__2467 (
            .O(N__11968),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__2466 (
            .O(N__11965),
            .I(N__11962));
    LocalMux I__2465 (
            .O(N__11962),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__2464 (
            .O(N__11959),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__2463 (
            .O(N__11956),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__2462 (
            .O(N__11953),
            .I(N__11948));
    InMux I__2461 (
            .O(N__11952),
            .I(N__11938));
    InMux I__2460 (
            .O(N__11951),
            .I(N__11938));
    InMux I__2459 (
            .O(N__11948),
            .I(N__11938));
    InMux I__2458 (
            .O(N__11947),
            .I(N__11938));
    LocalMux I__2457 (
            .O(N__11938),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0));
    CascadeMux I__2456 (
            .O(N__11935),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_));
    InMux I__2455 (
            .O(N__11932),
            .I(N__11929));
    LocalMux I__2454 (
            .O(N__11929),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_7));
    CascadeMux I__2453 (
            .O(N__11926),
            .I(N__11921));
    InMux I__2452 (
            .O(N__11925),
            .I(N__11908));
    InMux I__2451 (
            .O(N__11924),
            .I(N__11908));
    InMux I__2450 (
            .O(N__11921),
            .I(N__11908));
    InMux I__2449 (
            .O(N__11920),
            .I(N__11901));
    InMux I__2448 (
            .O(N__11919),
            .I(N__11901));
    InMux I__2447 (
            .O(N__11918),
            .I(N__11901));
    InMux I__2446 (
            .O(N__11917),
            .I(N__11893));
    InMux I__2445 (
            .O(N__11916),
            .I(N__11893));
    InMux I__2444 (
            .O(N__11915),
            .I(N__11890));
    LocalMux I__2443 (
            .O(N__11908),
            .I(N__11887));
    LocalMux I__2442 (
            .O(N__11901),
            .I(N__11884));
    InMux I__2441 (
            .O(N__11900),
            .I(N__11881));
    InMux I__2440 (
            .O(N__11899),
            .I(N__11876));
    InMux I__2439 (
            .O(N__11898),
            .I(N__11876));
    LocalMux I__2438 (
            .O(N__11893),
            .I(N__11873));
    LocalMux I__2437 (
            .O(N__11890),
            .I(N__11870));
    Span4Mux_v I__2436 (
            .O(N__11887),
            .I(N__11861));
    Span4Mux_v I__2435 (
            .O(N__11884),
            .I(N__11861));
    LocalMux I__2434 (
            .O(N__11881),
            .I(N__11861));
    LocalMux I__2433 (
            .O(N__11876),
            .I(N__11861));
    Span4Mux_s2_v I__2432 (
            .O(N__11873),
            .I(N__11858));
    Odrv4 I__2431 (
            .O(N__11870),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2430 (
            .O(N__11861),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2429 (
            .O(N__11858),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    CascadeMux I__2428 (
            .O(N__11851),
            .I(N__11848));
    InMux I__2427 (
            .O(N__11848),
            .I(N__11845));
    LocalMux I__2426 (
            .O(N__11845),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__2425 (
            .O(N__11842),
            .I(N__11839));
    LocalMux I__2424 (
            .O(N__11839),
            .I(beamY_RNIALEQZ0Z_9));
    InMux I__2423 (
            .O(N__11836),
            .I(N__11833));
    LocalMux I__2422 (
            .O(N__11833),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151));
    InMux I__2421 (
            .O(N__11830),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__2420 (
            .O(N__11827),
            .I(N__11824));
    LocalMux I__2419 (
            .O(N__11824),
            .I(beamY_RNIALEQ_1Z0Z_9));
    InMux I__2418 (
            .O(N__11821),
            .I(N__11818));
    LocalMux I__2417 (
            .O(N__11818),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251));
    InMux I__2416 (
            .O(N__11815),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__2415 (
            .O(N__11812),
            .I(N__11807));
    InMux I__2414 (
            .O(N__11811),
            .I(N__11804));
    InMux I__2413 (
            .O(N__11810),
            .I(N__11801));
    LocalMux I__2412 (
            .O(N__11807),
            .I(N__11798));
    LocalMux I__2411 (
            .O(N__11804),
            .I(N__11788));
    LocalMux I__2410 (
            .O(N__11801),
            .I(N__11781));
    Span4Mux_s2_v I__2409 (
            .O(N__11798),
            .I(N__11781));
    InMux I__2408 (
            .O(N__11797),
            .I(N__11774));
    InMux I__2407 (
            .O(N__11796),
            .I(N__11774));
    InMux I__2406 (
            .O(N__11795),
            .I(N__11774));
    InMux I__2405 (
            .O(N__11794),
            .I(N__11765));
    InMux I__2404 (
            .O(N__11793),
            .I(N__11765));
    InMux I__2403 (
            .O(N__11792),
            .I(N__11765));
    InMux I__2402 (
            .O(N__11791),
            .I(N__11765));
    Span4Mux_s2_v I__2401 (
            .O(N__11788),
            .I(N__11762));
    InMux I__2400 (
            .O(N__11787),
            .I(N__11759));
    InMux I__2399 (
            .O(N__11786),
            .I(N__11756));
    Span4Mux_v I__2398 (
            .O(N__11781),
            .I(N__11753));
    LocalMux I__2397 (
            .O(N__11774),
            .I(N__11746));
    LocalMux I__2396 (
            .O(N__11765),
            .I(N__11746));
    Span4Mux_h I__2395 (
            .O(N__11762),
            .I(N__11746));
    LocalMux I__2394 (
            .O(N__11759),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    LocalMux I__2393 (
            .O(N__11756),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2392 (
            .O(N__11753),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2391 (
            .O(N__11746),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    InMux I__2390 (
            .O(N__11737),
            .I(N__11734));
    LocalMux I__2389 (
            .O(N__11734),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0));
    InMux I__2388 (
            .O(N__11731),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__2387 (
            .O(N__11728),
            .I(N__11725));
    InMux I__2386 (
            .O(N__11725),
            .I(N__11722));
    LocalMux I__2385 (
            .O(N__11722),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1));
    InMux I__2384 (
            .O(N__11719),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3));
    CascadeMux I__2383 (
            .O(N__11716),
            .I(N__11713));
    InMux I__2382 (
            .O(N__11713),
            .I(N__11710));
    LocalMux I__2381 (
            .O(N__11710),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1));
    InMux I__2380 (
            .O(N__11707),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__2379 (
            .O(N__11704),
            .I(N__11701));
    LocalMux I__2378 (
            .O(N__11701),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__2377 (
            .O(N__11698),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__2376 (
            .O(N__11695),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__2375 (
            .O(N__11692),
            .I(N__11688));
    InMux I__2374 (
            .O(N__11691),
            .I(N__11678));
    InMux I__2373 (
            .O(N__11688),
            .I(N__11678));
    InMux I__2372 (
            .O(N__11687),
            .I(N__11678));
    InMux I__2371 (
            .O(N__11686),
            .I(N__11675));
    InMux I__2370 (
            .O(N__11685),
            .I(N__11672));
    LocalMux I__2369 (
            .O(N__11678),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    LocalMux I__2368 (
            .O(N__11675),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    LocalMux I__2367 (
            .O(N__11672),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    InMux I__2366 (
            .O(N__11665),
            .I(N__11662));
    LocalMux I__2365 (
            .O(N__11662),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921));
    InMux I__2364 (
            .O(N__11659),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__2363 (
            .O(N__11656),
            .I(N__11653));
    InMux I__2362 (
            .O(N__11653),
            .I(N__11650));
    LocalMux I__2361 (
            .O(N__11650),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51));
    InMux I__2360 (
            .O(N__11647),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__2359 (
            .O(N__11644),
            .I(N__11641));
    LocalMux I__2358 (
            .O(N__11641),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum1_4));
    InMux I__2357 (
            .O(N__11638),
            .I(N__11635));
    LocalMux I__2356 (
            .O(N__11635),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum0_4));
    CascadeMux I__2355 (
            .O(N__11632),
            .I(un7_pixel_0_axb4_cascade_));
    CascadeMux I__2354 (
            .O(N__11629),
            .I(N__11625));
    InMux I__2353 (
            .O(N__11628),
            .I(N__11620));
    InMux I__2352 (
            .O(N__11625),
            .I(N__11620));
    LocalMux I__2351 (
            .O(N__11620),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum1_5));
    InMux I__2350 (
            .O(N__11617),
            .I(N__11614));
    LocalMux I__2349 (
            .O(N__11614),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum0_5));
    CascadeMux I__2348 (
            .O(N__11611),
            .I(N__11608));
    InMux I__2347 (
            .O(N__11608),
            .I(N__11605));
    LocalMux I__2346 (
            .O(N__11605),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    InMux I__2345 (
            .O(N__11602),
            .I(un4_pixel_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__2344 (
            .O(N__11599),
            .I(N__11596));
    LocalMux I__2343 (
            .O(N__11596),
            .I(N__11593));
    Span4Mux_v I__2342 (
            .O(N__11593),
            .I(N__11589));
    InMux I__2341 (
            .O(N__11592),
            .I(N__11586));
    Odrv4 I__2340 (
            .O(N__11589),
            .I(un7_pixel_0_axb4));
    LocalMux I__2339 (
            .O(N__11586),
            .I(un7_pixel_0_axb4));
    CascadeMux I__2338 (
            .O(N__11581),
            .I(N__11578));
    InMux I__2337 (
            .O(N__11578),
            .I(N__11575));
    LocalMux I__2336 (
            .O(N__11575),
            .I(N__11572));
    Odrv12 I__2335 (
            .O(N__11572),
            .I(if_generate_plus_mult1_un47_sum_m_2));
    CascadeMux I__2334 (
            .O(N__11569),
            .I(N__11566));
    InMux I__2333 (
            .O(N__11566),
            .I(N__11563));
    LocalMux I__2332 (
            .O(N__11563),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__2331 (
            .O(N__11560),
            .I(un4_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__2330 (
            .O(N__11557),
            .I(N__11553));
    CascadeMux I__2329 (
            .O(N__11556),
            .I(N__11550));
    InMux I__2328 (
            .O(N__11553),
            .I(N__11545));
    InMux I__2327 (
            .O(N__11550),
            .I(N__11545));
    LocalMux I__2326 (
            .O(N__11545),
            .I(un7_pixel_0_axb4_i));
    InMux I__2325 (
            .O(N__11542),
            .I(N__11539));
    LocalMux I__2324 (
            .O(N__11539),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__2323 (
            .O(N__11536),
            .I(un4_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2322 (
            .O(N__11533),
            .I(N__11530));
    LocalMux I__2321 (
            .O(N__11530),
            .I(un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__2320 (
            .O(N__11527),
            .I(un4_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2319 (
            .O(N__11524),
            .I(N__11521));
    LocalMux I__2318 (
            .O(N__11521),
            .I(N__11518));
    Span4Mux_h I__2317 (
            .O(N__11518),
            .I(N__11512));
    InMux I__2316 (
            .O(N__11517),
            .I(N__11509));
    InMux I__2315 (
            .O(N__11516),
            .I(N__11506));
    InMux I__2314 (
            .O(N__11515),
            .I(N__11503));
    Odrv4 I__2313 (
            .O(N__11512),
            .I(un7_pixel_0_axb3));
    LocalMux I__2312 (
            .O(N__11509),
            .I(un7_pixel_0_axb3));
    LocalMux I__2311 (
            .O(N__11506),
            .I(un7_pixel_0_axb3));
    LocalMux I__2310 (
            .O(N__11503),
            .I(un7_pixel_0_axb3));
    InMux I__2309 (
            .O(N__11494),
            .I(N__11491));
    LocalMux I__2308 (
            .O(N__11491),
            .I(N__11488));
    Odrv4 I__2307 (
            .O(N__11488),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum1_3));
    InMux I__2306 (
            .O(N__11485),
            .I(N__11482));
    LocalMux I__2305 (
            .O(N__11482),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum0_3));
    InMux I__2304 (
            .O(N__11479),
            .I(N__11476));
    LocalMux I__2303 (
            .O(N__11476),
            .I(if_generate_plus_mult1_un47_sum_m_3));
    InMux I__2302 (
            .O(N__11473),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2));
    InMux I__2301 (
            .O(N__11470),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3));
    InMux I__2300 (
            .O(N__11467),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4));
    InMux I__2299 (
            .O(N__11464),
            .I(N__11461));
    LocalMux I__2298 (
            .O(N__11461),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum0_2));
    InMux I__2297 (
            .O(N__11458),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1));
    InMux I__2296 (
            .O(N__11455),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2));
    InMux I__2295 (
            .O(N__11452),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3));
    InMux I__2294 (
            .O(N__11449),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4));
    CascadeMux I__2293 (
            .O(N__11446),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_));
    InMux I__2292 (
            .O(N__11443),
            .I(N__11440));
    LocalMux I__2291 (
            .O(N__11440),
            .I(g1_0_0_0_1));
    InMux I__2290 (
            .O(N__11437),
            .I(N__11430));
    InMux I__2289 (
            .O(N__11436),
            .I(N__11427));
    InMux I__2288 (
            .O(N__11435),
            .I(N__11422));
    InMux I__2287 (
            .O(N__11434),
            .I(N__11422));
    InMux I__2286 (
            .O(N__11433),
            .I(N__11419));
    LocalMux I__2285 (
            .O(N__11430),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0));
    LocalMux I__2284 (
            .O(N__11427),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0));
    LocalMux I__2283 (
            .O(N__11422),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0));
    LocalMux I__2282 (
            .O(N__11419),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0));
    CascadeMux I__2281 (
            .O(N__11410),
            .I(g3_0_0_0_cascade_));
    InMux I__2280 (
            .O(N__11407),
            .I(N__11404));
    LocalMux I__2279 (
            .O(N__11404),
            .I(g1_4_0_0_0));
    InMux I__2278 (
            .O(N__11401),
            .I(N__11398));
    LocalMux I__2277 (
            .O(N__11398),
            .I(N_1869_0_0));
    InMux I__2276 (
            .O(N__11395),
            .I(N__11392));
    LocalMux I__2275 (
            .O(N__11392),
            .I(N_1870_0_0));
    CascadeMux I__2274 (
            .O(N__11389),
            .I(font_un127_pixel_6_ns_1_0_0_cascade_));
    InMux I__2273 (
            .O(N__11386),
            .I(N__11380));
    InMux I__2272 (
            .O(N__11385),
            .I(N__11380));
    LocalMux I__2271 (
            .O(N__11380),
            .I(font_un13_pixel_0_1_0_0_22));
    InMux I__2270 (
            .O(N__11377),
            .I(N__11374));
    LocalMux I__2269 (
            .O(N__11374),
            .I(N__11371));
    Odrv4 I__2268 (
            .O(N__11371),
            .I(N_520));
    CascadeMux I__2267 (
            .O(N__11368),
            .I(N__11365));
    InMux I__2266 (
            .O(N__11365),
            .I(N__11362));
    LocalMux I__2265 (
            .O(N__11362),
            .I(N__11359));
    Span4Mux_v I__2264 (
            .O(N__11359),
            .I(N__11356));
    Odrv4 I__2263 (
            .O(N__11356),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__2262 (
            .O(N__11353),
            .I(N__11350));
    InMux I__2261 (
            .O(N__11350),
            .I(N__11347));
    LocalMux I__2260 (
            .O(N__11347),
            .I(N__11344));
    Span4Mux_h I__2259 (
            .O(N__11344),
            .I(N__11341));
    Odrv4 I__2258 (
            .O(N__11341),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_iZ0));
    InMux I__2257 (
            .O(N__11338),
            .I(N__11334));
    SRMux I__2256 (
            .O(N__11337),
            .I(N__11331));
    LocalMux I__2255 (
            .O(N__11334),
            .I(N__11328));
    LocalMux I__2254 (
            .O(N__11331),
            .I(N__11325));
    Span4Mux_h I__2253 (
            .O(N__11328),
            .I(N__11322));
    Odrv4 I__2252 (
            .O(N__11325),
            .I(beamY_RNIJ0DBZ0Z_8));
    Odrv4 I__2251 (
            .O(N__11322),
            .I(beamY_RNIJ0DBZ0Z_8));
    IoInMux I__2250 (
            .O(N__11317),
            .I(N__11314));
    LocalMux I__2249 (
            .O(N__11314),
            .I(N__11310));
    IoInMux I__2248 (
            .O(N__11313),
            .I(N__11307));
    Span4Mux_s2_v I__2247 (
            .O(N__11310),
            .I(N__11304));
    LocalMux I__2246 (
            .O(N__11307),
            .I(N__11301));
    Span4Mux_v I__2245 (
            .O(N__11304),
            .I(N__11298));
    Span4Mux_s1_v I__2244 (
            .O(N__11301),
            .I(N__11295));
    Span4Mux_v I__2243 (
            .O(N__11298),
            .I(N__11292));
    Span4Mux_v I__2242 (
            .O(N__11295),
            .I(N__11289));
    Odrv4 I__2241 (
            .O(N__11292),
            .I(VSync_c));
    Odrv4 I__2240 (
            .O(N__11289),
            .I(VSync_c));
    CascadeMux I__2239 (
            .O(N__11284),
            .I(N__11281));
    InMux I__2238 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__2237 (
            .O(N__11278),
            .I(N__11275));
    Odrv4 I__2236 (
            .O(N__11275),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_iZ0));
    InMux I__2235 (
            .O(N__11272),
            .I(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1));
    InMux I__2234 (
            .O(N__11269),
            .I(N__11266));
    LocalMux I__2233 (
            .O(N__11266),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0));
    CascadeMux I__2232 (
            .O(N__11263),
            .I(N__11260));
    InMux I__2231 (
            .O(N__11260),
            .I(N__11256));
    InMux I__2230 (
            .O(N__11259),
            .I(N__11253));
    LocalMux I__2229 (
            .O(N__11256),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0));
    LocalMux I__2228 (
            .O(N__11253),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0));
    InMux I__2227 (
            .O(N__11248),
            .I(N__11245));
    LocalMux I__2226 (
            .O(N__11245),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321));
    InMux I__2225 (
            .O(N__11242),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__2224 (
            .O(N__11239),
            .I(N__11236));
    LocalMux I__2223 (
            .O(N__11236),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0));
    CascadeMux I__2222 (
            .O(N__11233),
            .I(N__11229));
    CascadeMux I__2221 (
            .O(N__11232),
            .I(N__11226));
    InMux I__2220 (
            .O(N__11229),
            .I(N__11221));
    InMux I__2219 (
            .O(N__11226),
            .I(N__11221));
    LocalMux I__2218 (
            .O(N__11221),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5));
    InMux I__2217 (
            .O(N__11218),
            .I(N__11215));
    LocalMux I__2216 (
            .O(N__11215),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__2215 (
            .O(N__11212),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__2214 (
            .O(N__11209),
            .I(N__11206));
    LocalMux I__2213 (
            .O(N__11206),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__2212 (
            .O(N__11203),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__2211 (
            .O(N__11200),
            .I(N__11196));
    InMux I__2210 (
            .O(N__11199),
            .I(N__11192));
    InMux I__2209 (
            .O(N__11196),
            .I(N__11187));
    InMux I__2208 (
            .O(N__11195),
            .I(N__11187));
    LocalMux I__2207 (
            .O(N__11192),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1));
    LocalMux I__2206 (
            .O(N__11187),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1));
    CascadeMux I__2205 (
            .O(N__11182),
            .I(N__11179));
    InMux I__2204 (
            .O(N__11179),
            .I(N__11176));
    LocalMux I__2203 (
            .O(N__11176),
            .I(N__11173));
    Span4Mux_v I__2202 (
            .O(N__11173),
            .I(N__11170));
    Odrv4 I__2201 (
            .O(N__11170),
            .I(un14_visibleylt9_0));
    CascadeMux I__2200 (
            .O(N__11167),
            .I(N__11164));
    InMux I__2199 (
            .O(N__11164),
            .I(N__11161));
    LocalMux I__2198 (
            .O(N__11161),
            .I(un14_visibleylt4_0));
    CascadeMux I__2197 (
            .O(N__11158),
            .I(un3_beamx_5_cascade_));
    InMux I__2196 (
            .O(N__11155),
            .I(N__11152));
    LocalMux I__2195 (
            .O(N__11152),
            .I(N__11149));
    Span4Mux_h I__2194 (
            .O(N__11149),
            .I(N__11146));
    Odrv4 I__2193 (
            .O(N__11146),
            .I(N_324_0_0_0));
    InMux I__2192 (
            .O(N__11143),
            .I(N__11140));
    LocalMux I__2191 (
            .O(N__11140),
            .I(N__11137));
    Span4Mux_h I__2190 (
            .O(N__11137),
            .I(N__11134));
    Odrv4 I__2189 (
            .O(N__11134),
            .I(N_303_0_0_0));
    CascadeMux I__2188 (
            .O(N__11131),
            .I(N__11125));
    CascadeMux I__2187 (
            .O(N__11130),
            .I(N__11120));
    CascadeMux I__2186 (
            .O(N__11129),
            .I(N__11116));
    CascadeMux I__2185 (
            .O(N__11128),
            .I(N__11113));
    InMux I__2184 (
            .O(N__11125),
            .I(N__11109));
    InMux I__2183 (
            .O(N__11124),
            .I(N__11106));
    InMux I__2182 (
            .O(N__11123),
            .I(N__11103));
    InMux I__2181 (
            .O(N__11120),
            .I(N__11100));
    InMux I__2180 (
            .O(N__11119),
            .I(N__11095));
    InMux I__2179 (
            .O(N__11116),
            .I(N__11095));
    InMux I__2178 (
            .O(N__11113),
            .I(N__11092));
    InMux I__2177 (
            .O(N__11112),
            .I(N__11085));
    LocalMux I__2176 (
            .O(N__11109),
            .I(N__11078));
    LocalMux I__2175 (
            .O(N__11106),
            .I(N__11078));
    LocalMux I__2174 (
            .O(N__11103),
            .I(N__11078));
    LocalMux I__2173 (
            .O(N__11100),
            .I(N__11073));
    LocalMux I__2172 (
            .O(N__11095),
            .I(N__11073));
    LocalMux I__2171 (
            .O(N__11092),
            .I(N__11070));
    InMux I__2170 (
            .O(N__11091),
            .I(N__11067));
    InMux I__2169 (
            .O(N__11090),
            .I(N__11064));
    InMux I__2168 (
            .O(N__11089),
            .I(N__11061));
    InMux I__2167 (
            .O(N__11088),
            .I(N__11058));
    LocalMux I__2166 (
            .O(N__11085),
            .I(N__11055));
    Span4Mux_v I__2165 (
            .O(N__11078),
            .I(N__11052));
    Span4Mux_v I__2164 (
            .O(N__11073),
            .I(N__11049));
    Span12Mux_s7_h I__2163 (
            .O(N__11070),
            .I(N__11044));
    LocalMux I__2162 (
            .O(N__11067),
            .I(N__11044));
    LocalMux I__2161 (
            .O(N__11064),
            .I(beamYZ0Z_0));
    LocalMux I__2160 (
            .O(N__11061),
            .I(beamYZ0Z_0));
    LocalMux I__2159 (
            .O(N__11058),
            .I(beamYZ0Z_0));
    Odrv4 I__2158 (
            .O(N__11055),
            .I(beamYZ0Z_0));
    Odrv4 I__2157 (
            .O(N__11052),
            .I(beamYZ0Z_0));
    Odrv4 I__2156 (
            .O(N__11049),
            .I(beamYZ0Z_0));
    Odrv12 I__2155 (
            .O(N__11044),
            .I(beamYZ0Z_0));
    InMux I__2154 (
            .O(N__11029),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__2153 (
            .O(N__11026),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__2152 (
            .O(N__11023),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__2151 (
            .O(N__11020),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2150 (
            .O(N__11017),
            .I(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_));
    InMux I__2149 (
            .O(N__11014),
            .I(N__11011));
    LocalMux I__2148 (
            .O(N__11011),
            .I(font_un13_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__2147 (
            .O(N__11008),
            .I(N__11001));
    InMux I__2146 (
            .O(N__11007),
            .I(N__10998));
    InMux I__2145 (
            .O(N__11006),
            .I(N__10993));
    InMux I__2144 (
            .O(N__11005),
            .I(N__10993));
    InMux I__2143 (
            .O(N__11004),
            .I(N__10988));
    LocalMux I__2142 (
            .O(N__11001),
            .I(N__10982));
    LocalMux I__2141 (
            .O(N__10998),
            .I(N__10979));
    LocalMux I__2140 (
            .O(N__10993),
            .I(N__10976));
    InMux I__2139 (
            .O(N__10992),
            .I(N__10973));
    CascadeMux I__2138 (
            .O(N__10991),
            .I(N__10970));
    LocalMux I__2137 (
            .O(N__10988),
            .I(N__10966));
    InMux I__2136 (
            .O(N__10987),
            .I(N__10963));
    InMux I__2135 (
            .O(N__10986),
            .I(N__10960));
    InMux I__2134 (
            .O(N__10985),
            .I(N__10957));
    Span4Mux_h I__2133 (
            .O(N__10982),
            .I(N__10952));
    Span4Mux_h I__2132 (
            .O(N__10979),
            .I(N__10952));
    Span4Mux_h I__2131 (
            .O(N__10976),
            .I(N__10947));
    LocalMux I__2130 (
            .O(N__10973),
            .I(N__10947));
    InMux I__2129 (
            .O(N__10970),
            .I(N__10942));
    InMux I__2128 (
            .O(N__10969),
            .I(N__10942));
    Odrv12 I__2127 (
            .O(N__10966),
            .I(beamYZ0Z_7));
    LocalMux I__2126 (
            .O(N__10963),
            .I(beamYZ0Z_7));
    LocalMux I__2125 (
            .O(N__10960),
            .I(beamYZ0Z_7));
    LocalMux I__2124 (
            .O(N__10957),
            .I(beamYZ0Z_7));
    Odrv4 I__2123 (
            .O(N__10952),
            .I(beamYZ0Z_7));
    Odrv4 I__2122 (
            .O(N__10947),
            .I(beamYZ0Z_7));
    LocalMux I__2121 (
            .O(N__10942),
            .I(beamYZ0Z_7));
    InMux I__2120 (
            .O(N__10927),
            .I(N__10919));
    InMux I__2119 (
            .O(N__10926),
            .I(N__10919));
    InMux I__2118 (
            .O(N__10925),
            .I(N__10916));
    InMux I__2117 (
            .O(N__10924),
            .I(N__10908));
    LocalMux I__2116 (
            .O(N__10919),
            .I(N__10905));
    LocalMux I__2115 (
            .O(N__10916),
            .I(N__10902));
    InMux I__2114 (
            .O(N__10915),
            .I(N__10899));
    InMux I__2113 (
            .O(N__10914),
            .I(N__10896));
    InMux I__2112 (
            .O(N__10913),
            .I(N__10893));
    InMux I__2111 (
            .O(N__10912),
            .I(N__10888));
    InMux I__2110 (
            .O(N__10911),
            .I(N__10888));
    LocalMux I__2109 (
            .O(N__10908),
            .I(N__10881));
    Span4Mux_v I__2108 (
            .O(N__10905),
            .I(N__10874));
    Span4Mux_v I__2107 (
            .O(N__10902),
            .I(N__10874));
    LocalMux I__2106 (
            .O(N__10899),
            .I(N__10871));
    LocalMux I__2105 (
            .O(N__10896),
            .I(N__10864));
    LocalMux I__2104 (
            .O(N__10893),
            .I(N__10864));
    LocalMux I__2103 (
            .O(N__10888),
            .I(N__10864));
    InMux I__2102 (
            .O(N__10887),
            .I(N__10861));
    InMux I__2101 (
            .O(N__10886),
            .I(N__10854));
    InMux I__2100 (
            .O(N__10885),
            .I(N__10854));
    InMux I__2099 (
            .O(N__10884),
            .I(N__10854));
    Span4Mux_h I__2098 (
            .O(N__10881),
            .I(N__10851));
    InMux I__2097 (
            .O(N__10880),
            .I(N__10846));
    InMux I__2096 (
            .O(N__10879),
            .I(N__10846));
    Odrv4 I__2095 (
            .O(N__10874),
            .I(beamYZ0Z_9));
    Odrv4 I__2094 (
            .O(N__10871),
            .I(beamYZ0Z_9));
    Odrv4 I__2093 (
            .O(N__10864),
            .I(beamYZ0Z_9));
    LocalMux I__2092 (
            .O(N__10861),
            .I(beamYZ0Z_9));
    LocalMux I__2091 (
            .O(N__10854),
            .I(beamYZ0Z_9));
    Odrv4 I__2090 (
            .O(N__10851),
            .I(beamYZ0Z_9));
    LocalMux I__2089 (
            .O(N__10846),
            .I(beamYZ0Z_9));
    CascadeMux I__2088 (
            .O(N__10831),
            .I(N__10828));
    InMux I__2087 (
            .O(N__10828),
            .I(N__10825));
    LocalMux I__2086 (
            .O(N__10825),
            .I(N__10822));
    Odrv4 I__2085 (
            .O(N__10822),
            .I(un8_beamylto9_1));
    InMux I__2084 (
            .O(N__10819),
            .I(N__10814));
    InMux I__2083 (
            .O(N__10818),
            .I(N__10806));
    InMux I__2082 (
            .O(N__10817),
            .I(N__10806));
    LocalMux I__2081 (
            .O(N__10814),
            .I(N__10803));
    InMux I__2080 (
            .O(N__10813),
            .I(N__10800));
    InMux I__2079 (
            .O(N__10812),
            .I(N__10794));
    InMux I__2078 (
            .O(N__10811),
            .I(N__10794));
    LocalMux I__2077 (
            .O(N__10806),
            .I(N__10788));
    Span4Mux_h I__2076 (
            .O(N__10803),
            .I(N__10788));
    LocalMux I__2075 (
            .O(N__10800),
            .I(N__10785));
    InMux I__2074 (
            .O(N__10799),
            .I(N__10782));
    LocalMux I__2073 (
            .O(N__10794),
            .I(N__10778));
    InMux I__2072 (
            .O(N__10793),
            .I(N__10775));
    Span4Mux_v I__2071 (
            .O(N__10788),
            .I(N__10772));
    Span4Mux_v I__2070 (
            .O(N__10785),
            .I(N__10767));
    LocalMux I__2069 (
            .O(N__10782),
            .I(N__10767));
    InMux I__2068 (
            .O(N__10781),
            .I(N__10764));
    Span4Mux_v I__2067 (
            .O(N__10778),
            .I(N__10761));
    LocalMux I__2066 (
            .O(N__10775),
            .I(beamYZ0Z_8));
    Odrv4 I__2065 (
            .O(N__10772),
            .I(beamYZ0Z_8));
    Odrv4 I__2064 (
            .O(N__10767),
            .I(beamYZ0Z_8));
    LocalMux I__2063 (
            .O(N__10764),
            .I(beamYZ0Z_8));
    Odrv4 I__2062 (
            .O(N__10761),
            .I(beamYZ0Z_8));
    InMux I__2061 (
            .O(N__10750),
            .I(N__10747));
    LocalMux I__2060 (
            .O(N__10747),
            .I(N__10744));
    Odrv4 I__2059 (
            .O(N__10744),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0));
    InMux I__2058 (
            .O(N__10741),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__2057 (
            .O(N__10738),
            .I(un5_visibley_ac0_7_cascade_));
    InMux I__2056 (
            .O(N__10735),
            .I(N__10726));
    InMux I__2055 (
            .O(N__10734),
            .I(N__10726));
    InMux I__2054 (
            .O(N__10733),
            .I(N__10726));
    LocalMux I__2053 (
            .O(N__10726),
            .I(N__10723));
    Span4Mux_h I__2052 (
            .O(N__10723),
            .I(N__10720));
    Odrv4 I__2051 (
            .O(N__10720),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0));
    CascadeMux I__2050 (
            .O(N__10717),
            .I(beamY_4_rep1_RNICDQEZ0_cascade_));
    InMux I__2049 (
            .O(N__10714),
            .I(N__10708));
    InMux I__2048 (
            .O(N__10713),
            .I(N__10705));
    InMux I__2047 (
            .O(N__10712),
            .I(N__10700));
    InMux I__2046 (
            .O(N__10711),
            .I(N__10700));
    LocalMux I__2045 (
            .O(N__10708),
            .I(beamY_fastZ0Z_3));
    LocalMux I__2044 (
            .O(N__10705),
            .I(beamY_fastZ0Z_3));
    LocalMux I__2043 (
            .O(N__10700),
            .I(beamY_fastZ0Z_3));
    InMux I__2042 (
            .O(N__10693),
            .I(N__10688));
    InMux I__2041 (
            .O(N__10692),
            .I(N__10685));
    InMux I__2040 (
            .O(N__10691),
            .I(N__10682));
    LocalMux I__2039 (
            .O(N__10688),
            .I(N__10677));
    LocalMux I__2038 (
            .O(N__10685),
            .I(N__10674));
    LocalMux I__2037 (
            .O(N__10682),
            .I(N__10671));
    InMux I__2036 (
            .O(N__10681),
            .I(N__10666));
    InMux I__2035 (
            .O(N__10680),
            .I(N__10666));
    Span4Mux_h I__2034 (
            .O(N__10677),
            .I(N__10660));
    Span4Mux_h I__2033 (
            .O(N__10674),
            .I(N__10660));
    Span4Mux_v I__2032 (
            .O(N__10671),
            .I(N__10655));
    LocalMux I__2031 (
            .O(N__10666),
            .I(N__10655));
    InMux I__2030 (
            .O(N__10665),
            .I(N__10652));
    Odrv4 I__2029 (
            .O(N__10660),
            .I(un5_visibley_c2));
    Odrv4 I__2028 (
            .O(N__10655),
            .I(un5_visibley_c2));
    LocalMux I__2027 (
            .O(N__10652),
            .I(un5_visibley_c2));
    CascadeMux I__2026 (
            .O(N__10645),
            .I(N__10642));
    InMux I__2025 (
            .O(N__10642),
            .I(N__10638));
    InMux I__2024 (
            .O(N__10641),
            .I(N__10635));
    LocalMux I__2023 (
            .O(N__10638),
            .I(un11_visibley));
    LocalMux I__2022 (
            .O(N__10635),
            .I(un11_visibley));
    InMux I__2021 (
            .O(N__10630),
            .I(N__10627));
    LocalMux I__2020 (
            .O(N__10627),
            .I(N__10624));
    Odrv4 I__2019 (
            .O(N__10624),
            .I(un44));
    InMux I__2018 (
            .O(N__10621),
            .I(N__10618));
    LocalMux I__2017 (
            .O(N__10618),
            .I(Pixel_1_e_1));
    InMux I__2016 (
            .O(N__10615),
            .I(N__10607));
    InMux I__2015 (
            .O(N__10614),
            .I(N__10607));
    InMux I__2014 (
            .O(N__10613),
            .I(N__10602));
    InMux I__2013 (
            .O(N__10612),
            .I(N__10602));
    LocalMux I__2012 (
            .O(N__10607),
            .I(beamY_fastZ0Z_2));
    LocalMux I__2011 (
            .O(N__10602),
            .I(beamY_fastZ0Z_2));
    CascadeMux I__2010 (
            .O(N__10597),
            .I(N__10590));
    InMux I__2009 (
            .O(N__10596),
            .I(N__10587));
    InMux I__2008 (
            .O(N__10595),
            .I(N__10584));
    InMux I__2007 (
            .O(N__10594),
            .I(N__10579));
    InMux I__2006 (
            .O(N__10593),
            .I(N__10579));
    InMux I__2005 (
            .O(N__10590),
            .I(N__10576));
    LocalMux I__2004 (
            .O(N__10587),
            .I(beamY_4_repZ0Z1));
    LocalMux I__2003 (
            .O(N__10584),
            .I(beamY_4_repZ0Z1));
    LocalMux I__2002 (
            .O(N__10579),
            .I(beamY_4_repZ0Z1));
    LocalMux I__2001 (
            .O(N__10576),
            .I(beamY_4_repZ0Z1));
    CascadeMux I__2000 (
            .O(N__10567),
            .I(N__10564));
    InMux I__1999 (
            .O(N__10564),
            .I(N__10561));
    LocalMux I__1998 (
            .O(N__10561),
            .I(beamY_fast_RNIK8HHZ0Z_2));
    InMux I__1997 (
            .O(N__10558),
            .I(N__10549));
    InMux I__1996 (
            .O(N__10557),
            .I(N__10546));
    InMux I__1995 (
            .O(N__10556),
            .I(N__10540));
    InMux I__1994 (
            .O(N__10555),
            .I(N__10540));
    CascadeMux I__1993 (
            .O(N__10554),
            .I(N__10537));
    InMux I__1992 (
            .O(N__10553),
            .I(N__10534));
    CascadeMux I__1991 (
            .O(N__10552),
            .I(N__10529));
    LocalMux I__1990 (
            .O(N__10549),
            .I(N__10523));
    LocalMux I__1989 (
            .O(N__10546),
            .I(N__10520));
    InMux I__1988 (
            .O(N__10545),
            .I(N__10517));
    LocalMux I__1987 (
            .O(N__10540),
            .I(N__10514));
    InMux I__1986 (
            .O(N__10537),
            .I(N__10511));
    LocalMux I__1985 (
            .O(N__10534),
            .I(N__10508));
    InMux I__1984 (
            .O(N__10533),
            .I(N__10505));
    InMux I__1983 (
            .O(N__10532),
            .I(N__10500));
    InMux I__1982 (
            .O(N__10529),
            .I(N__10500));
    InMux I__1981 (
            .O(N__10528),
            .I(N__10493));
    InMux I__1980 (
            .O(N__10527),
            .I(N__10493));
    InMux I__1979 (
            .O(N__10526),
            .I(N__10493));
    Odrv12 I__1978 (
            .O(N__10523),
            .I(beamYZ0Z_6));
    Odrv4 I__1977 (
            .O(N__10520),
            .I(beamYZ0Z_6));
    LocalMux I__1976 (
            .O(N__10517),
            .I(beamYZ0Z_6));
    Odrv4 I__1975 (
            .O(N__10514),
            .I(beamYZ0Z_6));
    LocalMux I__1974 (
            .O(N__10511),
            .I(beamYZ0Z_6));
    Odrv4 I__1973 (
            .O(N__10508),
            .I(beamYZ0Z_6));
    LocalMux I__1972 (
            .O(N__10505),
            .I(beamYZ0Z_6));
    LocalMux I__1971 (
            .O(N__10500),
            .I(beamYZ0Z_6));
    LocalMux I__1970 (
            .O(N__10493),
            .I(beamYZ0Z_6));
    InMux I__1969 (
            .O(N__10474),
            .I(N__10469));
    InMux I__1968 (
            .O(N__10473),
            .I(N__10466));
    InMux I__1967 (
            .O(N__10472),
            .I(N__10459));
    LocalMux I__1966 (
            .O(N__10469),
            .I(N__10455));
    LocalMux I__1965 (
            .O(N__10466),
            .I(N__10448));
    InMux I__1964 (
            .O(N__10465),
            .I(N__10445));
    InMux I__1963 (
            .O(N__10464),
            .I(N__10440));
    InMux I__1962 (
            .O(N__10463),
            .I(N__10440));
    CascadeMux I__1961 (
            .O(N__10462),
            .I(N__10436));
    LocalMux I__1960 (
            .O(N__10459),
            .I(N__10432));
    InMux I__1959 (
            .O(N__10458),
            .I(N__10429));
    Span12Mux_s6_v I__1958 (
            .O(N__10455),
            .I(N__10426));
    InMux I__1957 (
            .O(N__10454),
            .I(N__10423));
    InMux I__1956 (
            .O(N__10453),
            .I(N__10420));
    InMux I__1955 (
            .O(N__10452),
            .I(N__10417));
    InMux I__1954 (
            .O(N__10451),
            .I(N__10414));
    Span4Mux_h I__1953 (
            .O(N__10448),
            .I(N__10411));
    LocalMux I__1952 (
            .O(N__10445),
            .I(N__10406));
    LocalMux I__1951 (
            .O(N__10440),
            .I(N__10406));
    InMux I__1950 (
            .O(N__10439),
            .I(N__10399));
    InMux I__1949 (
            .O(N__10436),
            .I(N__10399));
    InMux I__1948 (
            .O(N__10435),
            .I(N__10399));
    Odrv4 I__1947 (
            .O(N__10432),
            .I(beamYZ0Z_5));
    LocalMux I__1946 (
            .O(N__10429),
            .I(beamYZ0Z_5));
    Odrv12 I__1945 (
            .O(N__10426),
            .I(beamYZ0Z_5));
    LocalMux I__1944 (
            .O(N__10423),
            .I(beamYZ0Z_5));
    LocalMux I__1943 (
            .O(N__10420),
            .I(beamYZ0Z_5));
    LocalMux I__1942 (
            .O(N__10417),
            .I(beamYZ0Z_5));
    LocalMux I__1941 (
            .O(N__10414),
            .I(beamYZ0Z_5));
    Odrv4 I__1940 (
            .O(N__10411),
            .I(beamYZ0Z_5));
    Odrv12 I__1939 (
            .O(N__10406),
            .I(beamYZ0Z_5));
    LocalMux I__1938 (
            .O(N__10399),
            .I(beamYZ0Z_5));
    InMux I__1937 (
            .O(N__10378),
            .I(N__10375));
    LocalMux I__1936 (
            .O(N__10375),
            .I(beamY_RNIKOP3Z0Z_7));
    InMux I__1935 (
            .O(N__10372),
            .I(N__10369));
    LocalMux I__1934 (
            .O(N__10369),
            .I(un42lt10));
    InMux I__1933 (
            .O(N__10366),
            .I(N__10358));
    InMux I__1932 (
            .O(N__10365),
            .I(N__10355));
    InMux I__1931 (
            .O(N__10364),
            .I(N__10348));
    InMux I__1930 (
            .O(N__10363),
            .I(N__10348));
    InMux I__1929 (
            .O(N__10362),
            .I(N__10348));
    InMux I__1928 (
            .O(N__10361),
            .I(N__10345));
    LocalMux I__1927 (
            .O(N__10358),
            .I(un5_visibley_c7));
    LocalMux I__1926 (
            .O(N__10355),
            .I(un5_visibley_c7));
    LocalMux I__1925 (
            .O(N__10348),
            .I(un5_visibley_c7));
    LocalMux I__1924 (
            .O(N__10345),
            .I(un5_visibley_c7));
    InMux I__1923 (
            .O(N__10336),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1922 (
            .O(N__10333),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__1921 (
            .O(N__10330),
            .I(N__10324));
    InMux I__1920 (
            .O(N__10329),
            .I(N__10324));
    LocalMux I__1919 (
            .O(N__10324),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__1918 (
            .O(N__10321),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__1917 (
            .O(N__10318),
            .I(N__10315));
    LocalMux I__1916 (
            .O(N__10315),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0));
    InMux I__1915 (
            .O(N__10312),
            .I(N__10308));
    InMux I__1914 (
            .O(N__10311),
            .I(N__10305));
    LocalMux I__1913 (
            .O(N__10308),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5));
    LocalMux I__1912 (
            .O(N__10305),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5));
    CascadeMux I__1911 (
            .O(N__10300),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_));
    InMux I__1910 (
            .O(N__10297),
            .I(N__10294));
    LocalMux I__1909 (
            .O(N__10294),
            .I(Pixel_1_RNOZ0Z_19));
    InMux I__1908 (
            .O(N__10291),
            .I(N__10288));
    LocalMux I__1907 (
            .O(N__10288),
            .I(un1_visiblex_27));
    CascadeMux I__1906 (
            .O(N__10285),
            .I(N__10282));
    InMux I__1905 (
            .O(N__10282),
            .I(N__10279));
    LocalMux I__1904 (
            .O(N__10279),
            .I(N__10276));
    Span4Mux_h I__1903 (
            .O(N__10276),
            .I(N__10273));
    Odrv4 I__1902 (
            .O(N__10273),
            .I(un5_visibley_ac0_7));
    InMux I__1901 (
            .O(N__10270),
            .I(N__10267));
    LocalMux I__1900 (
            .O(N__10267),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8));
    InMux I__1899 (
            .O(N__10264),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1898 (
            .O(N__10261),
            .I(N__10258));
    InMux I__1897 (
            .O(N__10258),
            .I(N__10255));
    LocalMux I__1896 (
            .O(N__10255),
            .I(N__10252));
    Odrv4 I__1895 (
            .O(N__10252),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299));
    CascadeMux I__1894 (
            .O(N__10249),
            .I(N__10244));
    CascadeMux I__1893 (
            .O(N__10248),
            .I(N__10240));
    InMux I__1892 (
            .O(N__10247),
            .I(N__10236));
    InMux I__1891 (
            .O(N__10244),
            .I(N__10227));
    InMux I__1890 (
            .O(N__10243),
            .I(N__10227));
    InMux I__1889 (
            .O(N__10240),
            .I(N__10227));
    InMux I__1888 (
            .O(N__10239),
            .I(N__10227));
    LocalMux I__1887 (
            .O(N__10236),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0));
    LocalMux I__1886 (
            .O(N__10227),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0));
    InMux I__1885 (
            .O(N__10222),
            .I(N__10219));
    LocalMux I__1884 (
            .O(N__10219),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__1883 (
            .O(N__10216),
            .I(N__10213));
    LocalMux I__1882 (
            .O(N__10213),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__1881 (
            .O(N__10210),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__1880 (
            .O(N__10207),
            .I(N__10204));
    LocalMux I__1879 (
            .O(N__10204),
            .I(Pixel_1_RNOZ0Z_18));
    CascadeMux I__1878 (
            .O(N__10201),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_));
    InMux I__1877 (
            .O(N__10198),
            .I(N__10195));
    LocalMux I__1876 (
            .O(N__10195),
            .I(N__10191));
    InMux I__1875 (
            .O(N__10194),
            .I(N__10188));
    Odrv4 I__1874 (
            .O(N__10191),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf));
    LocalMux I__1873 (
            .O(N__10188),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf));
    InMux I__1872 (
            .O(N__10183),
            .I(N__10179));
    InMux I__1871 (
            .O(N__10182),
            .I(N__10176));
    LocalMux I__1870 (
            .O(N__10179),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0));
    LocalMux I__1869 (
            .O(N__10176),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0));
    InMux I__1868 (
            .O(N__10171),
            .I(N__10165));
    InMux I__1867 (
            .O(N__10170),
            .I(N__10165));
    LocalMux I__1866 (
            .O(N__10165),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0));
    InMux I__1865 (
            .O(N__10162),
            .I(N__10157));
    CascadeMux I__1864 (
            .O(N__10161),
            .I(N__10154));
    InMux I__1863 (
            .O(N__10160),
            .I(N__10141));
    LocalMux I__1862 (
            .O(N__10157),
            .I(N__10130));
    InMux I__1861 (
            .O(N__10154),
            .I(N__10120));
    InMux I__1860 (
            .O(N__10153),
            .I(N__10117));
    InMux I__1859 (
            .O(N__10152),
            .I(N__10110));
    InMux I__1858 (
            .O(N__10151),
            .I(N__10110));
    InMux I__1857 (
            .O(N__10150),
            .I(N__10110));
    InMux I__1856 (
            .O(N__10149),
            .I(N__10105));
    InMux I__1855 (
            .O(N__10148),
            .I(N__10105));
    InMux I__1854 (
            .O(N__10147),
            .I(N__10100));
    InMux I__1853 (
            .O(N__10146),
            .I(N__10100));
    InMux I__1852 (
            .O(N__10145),
            .I(N__10097));
    InMux I__1851 (
            .O(N__10144),
            .I(N__10092));
    LocalMux I__1850 (
            .O(N__10141),
            .I(N__10089));
    InMux I__1849 (
            .O(N__10140),
            .I(N__10076));
    InMux I__1848 (
            .O(N__10139),
            .I(N__10076));
    InMux I__1847 (
            .O(N__10138),
            .I(N__10076));
    InMux I__1846 (
            .O(N__10137),
            .I(N__10071));
    InMux I__1845 (
            .O(N__10136),
            .I(N__10071));
    InMux I__1844 (
            .O(N__10135),
            .I(N__10068));
    CascadeMux I__1843 (
            .O(N__10134),
            .I(N__10065));
    InMux I__1842 (
            .O(N__10133),
            .I(N__10061));
    Span4Mux_h I__1841 (
            .O(N__10130),
            .I(N__10058));
    InMux I__1840 (
            .O(N__10129),
            .I(N__10053));
    InMux I__1839 (
            .O(N__10128),
            .I(N__10053));
    InMux I__1838 (
            .O(N__10127),
            .I(N__10042));
    InMux I__1837 (
            .O(N__10126),
            .I(N__10042));
    InMux I__1836 (
            .O(N__10125),
            .I(N__10042));
    InMux I__1835 (
            .O(N__10124),
            .I(N__10042));
    InMux I__1834 (
            .O(N__10123),
            .I(N__10042));
    LocalMux I__1833 (
            .O(N__10120),
            .I(N__10029));
    LocalMux I__1832 (
            .O(N__10117),
            .I(N__10029));
    LocalMux I__1831 (
            .O(N__10110),
            .I(N__10029));
    LocalMux I__1830 (
            .O(N__10105),
            .I(N__10029));
    LocalMux I__1829 (
            .O(N__10100),
            .I(N__10029));
    LocalMux I__1828 (
            .O(N__10097),
            .I(N__10029));
    InMux I__1827 (
            .O(N__10096),
            .I(N__10026));
    InMux I__1826 (
            .O(N__10095),
            .I(N__10023));
    LocalMux I__1825 (
            .O(N__10092),
            .I(N__10018));
    Span4Mux_v I__1824 (
            .O(N__10089),
            .I(N__10018));
    InMux I__1823 (
            .O(N__10088),
            .I(N__10013));
    InMux I__1822 (
            .O(N__10087),
            .I(N__10013));
    InMux I__1821 (
            .O(N__10086),
            .I(N__10010));
    InMux I__1820 (
            .O(N__10085),
            .I(N__10007));
    InMux I__1819 (
            .O(N__10084),
            .I(N__10002));
    InMux I__1818 (
            .O(N__10083),
            .I(N__10002));
    LocalMux I__1817 (
            .O(N__10076),
            .I(N__9995));
    LocalMux I__1816 (
            .O(N__10071),
            .I(N__9995));
    LocalMux I__1815 (
            .O(N__10068),
            .I(N__9995));
    InMux I__1814 (
            .O(N__10065),
            .I(N__9992));
    InMux I__1813 (
            .O(N__10064),
            .I(N__9989));
    LocalMux I__1812 (
            .O(N__10061),
            .I(N__9986));
    Span4Mux_v I__1811 (
            .O(N__10058),
            .I(N__9979));
    LocalMux I__1810 (
            .O(N__10053),
            .I(N__9979));
    LocalMux I__1809 (
            .O(N__10042),
            .I(N__9979));
    Span4Mux_v I__1808 (
            .O(N__10029),
            .I(N__9976));
    LocalMux I__1807 (
            .O(N__10026),
            .I(un43lto1));
    LocalMux I__1806 (
            .O(N__10023),
            .I(un43lto1));
    Odrv4 I__1805 (
            .O(N__10018),
            .I(un43lto1));
    LocalMux I__1804 (
            .O(N__10013),
            .I(un43lto1));
    LocalMux I__1803 (
            .O(N__10010),
            .I(un43lto1));
    LocalMux I__1802 (
            .O(N__10007),
            .I(un43lto1));
    LocalMux I__1801 (
            .O(N__10002),
            .I(un43lto1));
    Odrv4 I__1800 (
            .O(N__9995),
            .I(un43lto1));
    LocalMux I__1799 (
            .O(N__9992),
            .I(un43lto1));
    LocalMux I__1798 (
            .O(N__9989),
            .I(un43lto1));
    Odrv12 I__1797 (
            .O(N__9986),
            .I(un43lto1));
    Odrv4 I__1796 (
            .O(N__9979),
            .I(un43lto1));
    Odrv4 I__1795 (
            .O(N__9976),
            .I(un43lto1));
    CascadeMux I__1794 (
            .O(N__9949),
            .I(un43lto4_1_cascade_));
    CascadeMux I__1793 (
            .O(N__9946),
            .I(un43lt10_cascade_));
    InMux I__1792 (
            .O(N__9943),
            .I(N__9940));
    LocalMux I__1791 (
            .O(N__9940),
            .I(un1_beamY_26));
    CascadeMux I__1790 (
            .O(N__9937),
            .I(N__9934));
    InMux I__1789 (
            .O(N__9934),
            .I(N__9931));
    LocalMux I__1788 (
            .O(N__9931),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__1787 (
            .O(N__9928),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1786 (
            .O(N__9925),
            .I(N__9922));
    LocalMux I__1785 (
            .O(N__9922),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93));
    InMux I__1784 (
            .O(N__9919),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__1783 (
            .O(N__9916),
            .I(N__9913));
    InMux I__1782 (
            .O(N__9913),
            .I(N__9910));
    LocalMux I__1781 (
            .O(N__9910),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3));
    InMux I__1780 (
            .O(N__9907),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1779 (
            .O(N__9904),
            .I(N__9901));
    InMux I__1778 (
            .O(N__9901),
            .I(N__9898));
    LocalMux I__1777 (
            .O(N__9898),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94));
    InMux I__1776 (
            .O(N__9895),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1775 (
            .O(N__9892),
            .I(N__9889));
    LocalMux I__1774 (
            .O(N__9889),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__1773 (
            .O(N__9886),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__1772 (
            .O(N__9883),
            .I(N__9878));
    InMux I__1771 (
            .O(N__9882),
            .I(N__9873));
    InMux I__1770 (
            .O(N__9881),
            .I(N__9864));
    InMux I__1769 (
            .O(N__9878),
            .I(N__9864));
    InMux I__1768 (
            .O(N__9877),
            .I(N__9864));
    InMux I__1767 (
            .O(N__9876),
            .I(N__9864));
    LocalMux I__1766 (
            .O(N__9873),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5));
    LocalMux I__1765 (
            .O(N__9864),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5));
    InMux I__1764 (
            .O(N__9859),
            .I(N__9856));
    LocalMux I__1763 (
            .O(N__9856),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__1762 (
            .O(N__9853),
            .I(N__9850));
    LocalMux I__1761 (
            .O(N__9850),
            .I(N__9847));
    Odrv4 I__1760 (
            .O(N__9847),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__1759 (
            .O(N__9844),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__1758 (
            .O(N__9841),
            .I(N__9838));
    InMux I__1757 (
            .O(N__9838),
            .I(N__9835));
    LocalMux I__1756 (
            .O(N__9835),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5));
    InMux I__1755 (
            .O(N__9832),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__1754 (
            .O(N__9829),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__1753 (
            .O(N__9826),
            .I(N__9823));
    LocalMux I__1752 (
            .O(N__9823),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0));
    InMux I__1751 (
            .O(N__9820),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__1750 (
            .O(N__9817),
            .I(N__9813));
    InMux I__1749 (
            .O(N__9816),
            .I(N__9804));
    InMux I__1748 (
            .O(N__9813),
            .I(N__9804));
    InMux I__1747 (
            .O(N__9812),
            .I(N__9804));
    InMux I__1746 (
            .O(N__9811),
            .I(N__9801));
    LocalMux I__1745 (
            .O(N__9804),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2));
    LocalMux I__1744 (
            .O(N__9801),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2));
    CascadeMux I__1743 (
            .O(N__9796),
            .I(N__9793));
    InMux I__1742 (
            .O(N__9793),
            .I(N__9790));
    LocalMux I__1741 (
            .O(N__9790),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1));
    InMux I__1740 (
            .O(N__9787),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__1739 (
            .O(N__9784),
            .I(N__9781));
    LocalMux I__1738 (
            .O(N__9781),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_7));
    CascadeMux I__1737 (
            .O(N__9778),
            .I(N__9775));
    InMux I__1736 (
            .O(N__9775),
            .I(N__9772));
    LocalMux I__1735 (
            .O(N__9772),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2));
    InMux I__1734 (
            .O(N__9769),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1733 (
            .O(N__9766),
            .I(N__9763));
    LocalMux I__1732 (
            .O(N__9763),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__1731 (
            .O(N__9760),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1730 (
            .O(N__9757),
            .I(N__9754));
    LocalMux I__1729 (
            .O(N__9754),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__1728 (
            .O(N__9751),
            .I(N__9743));
    CascadeMux I__1727 (
            .O(N__9750),
            .I(N__9737));
    CascadeMux I__1726 (
            .O(N__9749),
            .I(N__9733));
    CascadeMux I__1725 (
            .O(N__9748),
            .I(N__9729));
    CascadeMux I__1724 (
            .O(N__9747),
            .I(N__9726));
    CascadeMux I__1723 (
            .O(N__9746),
            .I(N__9723));
    InMux I__1722 (
            .O(N__9743),
            .I(N__9718));
    InMux I__1721 (
            .O(N__9742),
            .I(N__9718));
    InMux I__1720 (
            .O(N__9741),
            .I(N__9715));
    InMux I__1719 (
            .O(N__9740),
            .I(N__9712));
    InMux I__1718 (
            .O(N__9737),
            .I(N__9709));
    InMux I__1717 (
            .O(N__9736),
            .I(N__9696));
    InMux I__1716 (
            .O(N__9733),
            .I(N__9696));
    InMux I__1715 (
            .O(N__9732),
            .I(N__9696));
    InMux I__1714 (
            .O(N__9729),
            .I(N__9696));
    InMux I__1713 (
            .O(N__9726),
            .I(N__9696));
    InMux I__1712 (
            .O(N__9723),
            .I(N__9696));
    LocalMux I__1711 (
            .O(N__9718),
            .I(N__9693));
    LocalMux I__1710 (
            .O(N__9715),
            .I(N__9688));
    LocalMux I__1709 (
            .O(N__9712),
            .I(N__9688));
    LocalMux I__1708 (
            .O(N__9709),
            .I(N__9681));
    LocalMux I__1707 (
            .O(N__9696),
            .I(N__9681));
    Span4Mux_h I__1706 (
            .O(N__9693),
            .I(N__9681));
    Span4Mux_s2_v I__1705 (
            .O(N__9688),
            .I(N__9678));
    Odrv4 I__1704 (
            .O(N__9681),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1703 (
            .O(N__9678),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    CascadeMux I__1702 (
            .O(N__9673),
            .I(N__9670));
    InMux I__1701 (
            .O(N__9670),
            .I(N__9667));
    LocalMux I__1700 (
            .O(N__9667),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_0));
    CascadeMux I__1699 (
            .O(N__9664),
            .I(N__9661));
    InMux I__1698 (
            .O(N__9661),
            .I(N__9657));
    InMux I__1697 (
            .O(N__9660),
            .I(N__9653));
    LocalMux I__1696 (
            .O(N__9657),
            .I(N__9649));
    InMux I__1695 (
            .O(N__9656),
            .I(N__9646));
    LocalMux I__1694 (
            .O(N__9653),
            .I(N__9643));
    InMux I__1693 (
            .O(N__9652),
            .I(N__9640));
    Span4Mux_s3_h I__1692 (
            .O(N__9649),
            .I(N__9635));
    LocalMux I__1691 (
            .O(N__9646),
            .I(N__9635));
    Span4Mux_h I__1690 (
            .O(N__9643),
            .I(N__9632));
    LocalMux I__1689 (
            .O(N__9640),
            .I(N__9627));
    Span4Mux_v I__1688 (
            .O(N__9635),
            .I(N__9627));
    Odrv4 I__1687 (
            .O(N__9632),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1686 (
            .O(N__9627),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    InMux I__1685 (
            .O(N__9622),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__1684 (
            .O(N__9619),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__1683 (
            .O(N__9616),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__1682 (
            .O(N__9613),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__1681 (
            .O(N__9610),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__1680 (
            .O(N__9607),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_));
    CascadeMux I__1679 (
            .O(N__9604),
            .I(N__9601));
    InMux I__1678 (
            .O(N__9601),
            .I(N__9598));
    LocalMux I__1677 (
            .O(N__9598),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__1676 (
            .O(N__9595),
            .I(N__9591));
    CascadeMux I__1675 (
            .O(N__9594),
            .I(N__9587));
    LocalMux I__1674 (
            .O(N__9591),
            .I(N__9583));
    InMux I__1673 (
            .O(N__9590),
            .I(N__9578));
    InMux I__1672 (
            .O(N__9587),
            .I(N__9578));
    InMux I__1671 (
            .O(N__9586),
            .I(N__9574));
    Span4Mux_v I__1670 (
            .O(N__9583),
            .I(N__9569));
    LocalMux I__1669 (
            .O(N__9578),
            .I(N__9569));
    InMux I__1668 (
            .O(N__9577),
            .I(N__9566));
    LocalMux I__1667 (
            .O(N__9574),
            .I(N__9561));
    Span4Mux_h I__1666 (
            .O(N__9569),
            .I(N__9556));
    LocalMux I__1665 (
            .O(N__9566),
            .I(N__9556));
    CascadeMux I__1664 (
            .O(N__9565),
            .I(N__9553));
    InMux I__1663 (
            .O(N__9564),
            .I(N__9550));
    Span4Mux_s2_v I__1662 (
            .O(N__9561),
            .I(N__9547));
    Span4Mux_v I__1661 (
            .O(N__9556),
            .I(N__9544));
    InMux I__1660 (
            .O(N__9553),
            .I(N__9541));
    LocalMux I__1659 (
            .O(N__9550),
            .I(N__9538));
    Span4Mux_h I__1658 (
            .O(N__9547),
            .I(N__9535));
    Odrv4 I__1657 (
            .O(N__9544),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    LocalMux I__1656 (
            .O(N__9541),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1655 (
            .O(N__9538),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1654 (
            .O(N__9535),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1653 (
            .O(N__9526),
            .I(N__9523));
    InMux I__1652 (
            .O(N__9523),
            .I(N__9520));
    LocalMux I__1651 (
            .O(N__9520),
            .I(N__9517));
    Odrv4 I__1650 (
            .O(N__9517),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__1649 (
            .O(N__9514),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__1648 (
            .O(N__9511),
            .I(N__9508));
    LocalMux I__1647 (
            .O(N__9508),
            .I(N__9505));
    Odrv4 I__1646 (
            .O(N__9505),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__1645 (
            .O(N__9502),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__1644 (
            .O(N__9499),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__1643 (
            .O(N__9496),
            .I(N__9468));
    InMux I__1642 (
            .O(N__9495),
            .I(N__9468));
    InMux I__1641 (
            .O(N__9494),
            .I(N__9468));
    InMux I__1640 (
            .O(N__9493),
            .I(N__9468));
    InMux I__1639 (
            .O(N__9492),
            .I(N__9465));
    InMux I__1638 (
            .O(N__9491),
            .I(N__9460));
    InMux I__1637 (
            .O(N__9490),
            .I(N__9460));
    InMux I__1636 (
            .O(N__9489),
            .I(N__9447));
    InMux I__1635 (
            .O(N__9488),
            .I(N__9447));
    InMux I__1634 (
            .O(N__9487),
            .I(N__9447));
    InMux I__1633 (
            .O(N__9486),
            .I(N__9447));
    InMux I__1632 (
            .O(N__9485),
            .I(N__9447));
    InMux I__1631 (
            .O(N__9484),
            .I(N__9447));
    InMux I__1630 (
            .O(N__9483),
            .I(N__9434));
    InMux I__1629 (
            .O(N__9482),
            .I(N__9434));
    InMux I__1628 (
            .O(N__9481),
            .I(N__9434));
    InMux I__1627 (
            .O(N__9480),
            .I(N__9434));
    InMux I__1626 (
            .O(N__9479),
            .I(N__9415));
    InMux I__1625 (
            .O(N__9478),
            .I(N__9415));
    InMux I__1624 (
            .O(N__9477),
            .I(N__9415));
    LocalMux I__1623 (
            .O(N__9468),
            .I(N__9412));
    LocalMux I__1622 (
            .O(N__9465),
            .I(N__9403));
    LocalMux I__1621 (
            .O(N__9460),
            .I(N__9400));
    LocalMux I__1620 (
            .O(N__9447),
            .I(N__9397));
    InMux I__1619 (
            .O(N__9446),
            .I(N__9388));
    InMux I__1618 (
            .O(N__9445),
            .I(N__9388));
    InMux I__1617 (
            .O(N__9444),
            .I(N__9388));
    InMux I__1616 (
            .O(N__9443),
            .I(N__9388));
    LocalMux I__1615 (
            .O(N__9434),
            .I(N__9385));
    InMux I__1614 (
            .O(N__9433),
            .I(N__9372));
    InMux I__1613 (
            .O(N__9432),
            .I(N__9372));
    InMux I__1612 (
            .O(N__9431),
            .I(N__9372));
    InMux I__1611 (
            .O(N__9430),
            .I(N__9372));
    InMux I__1610 (
            .O(N__9429),
            .I(N__9372));
    InMux I__1609 (
            .O(N__9428),
            .I(N__9372));
    InMux I__1608 (
            .O(N__9427),
            .I(N__9369));
    InMux I__1607 (
            .O(N__9426),
            .I(N__9361));
    InMux I__1606 (
            .O(N__9425),
            .I(N__9361));
    InMux I__1605 (
            .O(N__9424),
            .I(N__9354));
    InMux I__1604 (
            .O(N__9423),
            .I(N__9354));
    InMux I__1603 (
            .O(N__9422),
            .I(N__9354));
    LocalMux I__1602 (
            .O(N__9415),
            .I(N__9349));
    Span4Mux_v I__1601 (
            .O(N__9412),
            .I(N__9349));
    InMux I__1600 (
            .O(N__9411),
            .I(N__9336));
    InMux I__1599 (
            .O(N__9410),
            .I(N__9336));
    InMux I__1598 (
            .O(N__9409),
            .I(N__9336));
    InMux I__1597 (
            .O(N__9408),
            .I(N__9336));
    InMux I__1596 (
            .O(N__9407),
            .I(N__9336));
    InMux I__1595 (
            .O(N__9406),
            .I(N__9336));
    Span4Mux_v I__1594 (
            .O(N__9403),
            .I(N__9331));
    Span4Mux_h I__1593 (
            .O(N__9400),
            .I(N__9331));
    Span4Mux_h I__1592 (
            .O(N__9397),
            .I(N__9328));
    LocalMux I__1591 (
            .O(N__9388),
            .I(N__9319));
    Span4Mux_h I__1590 (
            .O(N__9385),
            .I(N__9319));
    LocalMux I__1589 (
            .O(N__9372),
            .I(N__9319));
    LocalMux I__1588 (
            .O(N__9369),
            .I(N__9319));
    InMux I__1587 (
            .O(N__9368),
            .I(N__9316));
    InMux I__1586 (
            .O(N__9367),
            .I(N__9311));
    InMux I__1585 (
            .O(N__9366),
            .I(N__9311));
    LocalMux I__1584 (
            .O(N__9361),
            .I(un7_pixel_1_axb3));
    LocalMux I__1583 (
            .O(N__9354),
            .I(un7_pixel_1_axb3));
    Odrv4 I__1582 (
            .O(N__9349),
            .I(un7_pixel_1_axb3));
    LocalMux I__1581 (
            .O(N__9336),
            .I(un7_pixel_1_axb3));
    Odrv4 I__1580 (
            .O(N__9331),
            .I(un7_pixel_1_axb3));
    Odrv4 I__1579 (
            .O(N__9328),
            .I(un7_pixel_1_axb3));
    Odrv4 I__1578 (
            .O(N__9319),
            .I(un7_pixel_1_axb3));
    LocalMux I__1577 (
            .O(N__9316),
            .I(un7_pixel_1_axb3));
    LocalMux I__1576 (
            .O(N__9311),
            .I(un7_pixel_1_axb3));
    CascadeMux I__1575 (
            .O(N__9292),
            .I(un7_pixel_1_axb3_cascade_));
    CascadeMux I__1574 (
            .O(N__9289),
            .I(N__9280));
    CascadeMux I__1573 (
            .O(N__9288),
            .I(N__9273));
    InMux I__1572 (
            .O(N__9287),
            .I(N__9256));
    CascadeMux I__1571 (
            .O(N__9286),
            .I(N__9248));
    InMux I__1570 (
            .O(N__9285),
            .I(N__9238));
    InMux I__1569 (
            .O(N__9284),
            .I(N__9238));
    InMux I__1568 (
            .O(N__9283),
            .I(N__9238));
    InMux I__1567 (
            .O(N__9280),
            .I(N__9238));
    InMux I__1566 (
            .O(N__9279),
            .I(N__9229));
    InMux I__1565 (
            .O(N__9278),
            .I(N__9229));
    InMux I__1564 (
            .O(N__9277),
            .I(N__9229));
    InMux I__1563 (
            .O(N__9276),
            .I(N__9229));
    InMux I__1562 (
            .O(N__9273),
            .I(N__9220));
    InMux I__1561 (
            .O(N__9272),
            .I(N__9220));
    InMux I__1560 (
            .O(N__9271),
            .I(N__9220));
    InMux I__1559 (
            .O(N__9270),
            .I(N__9220));
    CascadeMux I__1558 (
            .O(N__9269),
            .I(N__9213));
    CascadeMux I__1557 (
            .O(N__9268),
            .I(N__9208));
    CascadeMux I__1556 (
            .O(N__9267),
            .I(N__9205));
    CascadeMux I__1555 (
            .O(N__9266),
            .I(N__9201));
    CascadeMux I__1554 (
            .O(N__9265),
            .I(N__9198));
    CascadeMux I__1553 (
            .O(N__9264),
            .I(N__9194));
    InMux I__1552 (
            .O(N__9263),
            .I(N__9189));
    InMux I__1551 (
            .O(N__9262),
            .I(N__9189));
    InMux I__1550 (
            .O(N__9261),
            .I(N__9184));
    InMux I__1549 (
            .O(N__9260),
            .I(N__9184));
    CascadeMux I__1548 (
            .O(N__9259),
            .I(N__9177));
    LocalMux I__1547 (
            .O(N__9256),
            .I(N__9173));
    InMux I__1546 (
            .O(N__9255),
            .I(N__9170));
    InMux I__1545 (
            .O(N__9254),
            .I(N__9157));
    InMux I__1544 (
            .O(N__9253),
            .I(N__9157));
    InMux I__1543 (
            .O(N__9252),
            .I(N__9157));
    InMux I__1542 (
            .O(N__9251),
            .I(N__9157));
    InMux I__1541 (
            .O(N__9248),
            .I(N__9157));
    InMux I__1540 (
            .O(N__9247),
            .I(N__9157));
    LocalMux I__1539 (
            .O(N__9238),
            .I(N__9150));
    LocalMux I__1538 (
            .O(N__9229),
            .I(N__9150));
    LocalMux I__1537 (
            .O(N__9220),
            .I(N__9150));
    InMux I__1536 (
            .O(N__9219),
            .I(N__9137));
    InMux I__1535 (
            .O(N__9218),
            .I(N__9137));
    InMux I__1534 (
            .O(N__9217),
            .I(N__9137));
    InMux I__1533 (
            .O(N__9216),
            .I(N__9137));
    InMux I__1532 (
            .O(N__9213),
            .I(N__9137));
    InMux I__1531 (
            .O(N__9212),
            .I(N__9137));
    InMux I__1530 (
            .O(N__9211),
            .I(N__9134));
    InMux I__1529 (
            .O(N__9208),
            .I(N__9129));
    InMux I__1528 (
            .O(N__9205),
            .I(N__9129));
    InMux I__1527 (
            .O(N__9204),
            .I(N__9118));
    InMux I__1526 (
            .O(N__9201),
            .I(N__9118));
    InMux I__1525 (
            .O(N__9198),
            .I(N__9118));
    InMux I__1524 (
            .O(N__9197),
            .I(N__9118));
    InMux I__1523 (
            .O(N__9194),
            .I(N__9118));
    LocalMux I__1522 (
            .O(N__9189),
            .I(N__9113));
    LocalMux I__1521 (
            .O(N__9184),
            .I(N__9113));
    InMux I__1520 (
            .O(N__9183),
            .I(N__9110));
    InMux I__1519 (
            .O(N__9182),
            .I(N__9105));
    InMux I__1518 (
            .O(N__9181),
            .I(N__9105));
    InMux I__1517 (
            .O(N__9180),
            .I(N__9098));
    InMux I__1516 (
            .O(N__9177),
            .I(N__9098));
    InMux I__1515 (
            .O(N__9176),
            .I(N__9098));
    Odrv4 I__1514 (
            .O(N__9173),
            .I(un7_pixel_1_axb1));
    LocalMux I__1513 (
            .O(N__9170),
            .I(un7_pixel_1_axb1));
    LocalMux I__1512 (
            .O(N__9157),
            .I(un7_pixel_1_axb1));
    Odrv4 I__1511 (
            .O(N__9150),
            .I(un7_pixel_1_axb1));
    LocalMux I__1510 (
            .O(N__9137),
            .I(un7_pixel_1_axb1));
    LocalMux I__1509 (
            .O(N__9134),
            .I(un7_pixel_1_axb1));
    LocalMux I__1508 (
            .O(N__9129),
            .I(un7_pixel_1_axb1));
    LocalMux I__1507 (
            .O(N__9118),
            .I(un7_pixel_1_axb1));
    Odrv4 I__1506 (
            .O(N__9113),
            .I(un7_pixel_1_axb1));
    LocalMux I__1505 (
            .O(N__9110),
            .I(un7_pixel_1_axb1));
    LocalMux I__1504 (
            .O(N__9105),
            .I(un7_pixel_1_axb1));
    LocalMux I__1503 (
            .O(N__9098),
            .I(un7_pixel_1_axb1));
    CascadeMux I__1502 (
            .O(N__9073),
            .I(N__9070));
    InMux I__1501 (
            .O(N__9070),
            .I(N__9067));
    LocalMux I__1500 (
            .O(N__9067),
            .I(N_532_i));
    InMux I__1499 (
            .O(N__9064),
            .I(N__9061));
    LocalMux I__1498 (
            .O(N__9061),
            .I(un117_pixel_2_6_i3_mux));
    CascadeMux I__1497 (
            .O(N__9058),
            .I(N__9047));
    CascadeMux I__1496 (
            .O(N__9057),
            .I(N__9044));
    CascadeMux I__1495 (
            .O(N__9056),
            .I(N__9041));
    CascadeMux I__1494 (
            .O(N__9055),
            .I(N__9036));
    CascadeMux I__1493 (
            .O(N__9054),
            .I(N__9033));
    CascadeMux I__1492 (
            .O(N__9053),
            .I(N__9021));
    CascadeMux I__1491 (
            .O(N__9052),
            .I(N__9013));
    CascadeMux I__1490 (
            .O(N__9051),
            .I(N__9007));
    InMux I__1489 (
            .O(N__9050),
            .I(N__8998));
    InMux I__1488 (
            .O(N__9047),
            .I(N__8998));
    InMux I__1487 (
            .O(N__9044),
            .I(N__8998));
    InMux I__1486 (
            .O(N__9041),
            .I(N__8998));
    CascadeMux I__1485 (
            .O(N__9040),
            .I(N__8992));
    InMux I__1484 (
            .O(N__9039),
            .I(N__8980));
    InMux I__1483 (
            .O(N__9036),
            .I(N__8980));
    InMux I__1482 (
            .O(N__9033),
            .I(N__8980));
    InMux I__1481 (
            .O(N__9032),
            .I(N__8980));
    CascadeMux I__1480 (
            .O(N__9031),
            .I(N__8977));
    CascadeMux I__1479 (
            .O(N__9030),
            .I(N__8973));
    CascadeMux I__1478 (
            .O(N__9029),
            .I(N__8970));
    InMux I__1477 (
            .O(N__9028),
            .I(N__8958));
    InMux I__1476 (
            .O(N__9027),
            .I(N__8958));
    InMux I__1475 (
            .O(N__9026),
            .I(N__8958));
    InMux I__1474 (
            .O(N__9025),
            .I(N__8958));
    InMux I__1473 (
            .O(N__9024),
            .I(N__8953));
    InMux I__1472 (
            .O(N__9021),
            .I(N__8953));
    CascadeMux I__1471 (
            .O(N__9020),
            .I(N__8947));
    CascadeMux I__1470 (
            .O(N__9019),
            .I(N__8944));
    CascadeMux I__1469 (
            .O(N__9018),
            .I(N__8939));
    CascadeMux I__1468 (
            .O(N__9017),
            .I(N__8933));
    InMux I__1467 (
            .O(N__9016),
            .I(N__8928));
    InMux I__1466 (
            .O(N__9013),
            .I(N__8928));
    InMux I__1465 (
            .O(N__9012),
            .I(N__8925));
    InMux I__1464 (
            .O(N__9011),
            .I(N__8918));
    InMux I__1463 (
            .O(N__9010),
            .I(N__8918));
    InMux I__1462 (
            .O(N__9007),
            .I(N__8918));
    LocalMux I__1461 (
            .O(N__8998),
            .I(N__8915));
    InMux I__1460 (
            .O(N__8997),
            .I(N__8902));
    InMux I__1459 (
            .O(N__8996),
            .I(N__8902));
    InMux I__1458 (
            .O(N__8995),
            .I(N__8902));
    InMux I__1457 (
            .O(N__8992),
            .I(N__8902));
    InMux I__1456 (
            .O(N__8991),
            .I(N__8902));
    InMux I__1455 (
            .O(N__8990),
            .I(N__8902));
    InMux I__1454 (
            .O(N__8989),
            .I(N__8899));
    LocalMux I__1453 (
            .O(N__8980),
            .I(N__8896));
    InMux I__1452 (
            .O(N__8977),
            .I(N__8881));
    InMux I__1451 (
            .O(N__8976),
            .I(N__8881));
    InMux I__1450 (
            .O(N__8973),
            .I(N__8881));
    InMux I__1449 (
            .O(N__8970),
            .I(N__8881));
    InMux I__1448 (
            .O(N__8969),
            .I(N__8881));
    InMux I__1447 (
            .O(N__8968),
            .I(N__8881));
    InMux I__1446 (
            .O(N__8967),
            .I(N__8881));
    LocalMux I__1445 (
            .O(N__8958),
            .I(N__8876));
    LocalMux I__1444 (
            .O(N__8953),
            .I(N__8876));
    InMux I__1443 (
            .O(N__8952),
            .I(N__8873));
    CascadeMux I__1442 (
            .O(N__8951),
            .I(N__8869));
    InMux I__1441 (
            .O(N__8950),
            .I(N__8864));
    InMux I__1440 (
            .O(N__8947),
            .I(N__8855));
    InMux I__1439 (
            .O(N__8944),
            .I(N__8855));
    InMux I__1438 (
            .O(N__8943),
            .I(N__8855));
    InMux I__1437 (
            .O(N__8942),
            .I(N__8855));
    InMux I__1436 (
            .O(N__8939),
            .I(N__8844));
    InMux I__1435 (
            .O(N__8938),
            .I(N__8844));
    InMux I__1434 (
            .O(N__8937),
            .I(N__8844));
    InMux I__1433 (
            .O(N__8936),
            .I(N__8844));
    InMux I__1432 (
            .O(N__8933),
            .I(N__8844));
    LocalMux I__1431 (
            .O(N__8928),
            .I(N__8831));
    LocalMux I__1430 (
            .O(N__8925),
            .I(N__8831));
    LocalMux I__1429 (
            .O(N__8918),
            .I(N__8831));
    Span4Mux_h I__1428 (
            .O(N__8915),
            .I(N__8831));
    LocalMux I__1427 (
            .O(N__8902),
            .I(N__8831));
    LocalMux I__1426 (
            .O(N__8899),
            .I(N__8831));
    Span4Mux_v I__1425 (
            .O(N__8896),
            .I(N__8822));
    LocalMux I__1424 (
            .O(N__8881),
            .I(N__8822));
    Span4Mux_v I__1423 (
            .O(N__8876),
            .I(N__8822));
    LocalMux I__1422 (
            .O(N__8873),
            .I(N__8822));
    InMux I__1421 (
            .O(N__8872),
            .I(N__8815));
    InMux I__1420 (
            .O(N__8869),
            .I(N__8815));
    InMux I__1419 (
            .O(N__8868),
            .I(N__8815));
    InMux I__1418 (
            .O(N__8867),
            .I(N__8812));
    LocalMux I__1417 (
            .O(N__8864),
            .I(un7_pixel_1_axb2));
    LocalMux I__1416 (
            .O(N__8855),
            .I(un7_pixel_1_axb2));
    LocalMux I__1415 (
            .O(N__8844),
            .I(un7_pixel_1_axb2));
    Odrv4 I__1414 (
            .O(N__8831),
            .I(un7_pixel_1_axb2));
    Odrv4 I__1413 (
            .O(N__8822),
            .I(un7_pixel_1_axb2));
    LocalMux I__1412 (
            .O(N__8815),
            .I(un7_pixel_1_axb2));
    LocalMux I__1411 (
            .O(N__8812),
            .I(un7_pixel_1_axb2));
    CascadeMux I__1410 (
            .O(N__8797),
            .I(N__8793));
    InMux I__1409 (
            .O(N__8796),
            .I(N__8779));
    InMux I__1408 (
            .O(N__8793),
            .I(N__8776));
    CascadeMux I__1407 (
            .O(N__8792),
            .I(N__8771));
    CascadeMux I__1406 (
            .O(N__8791),
            .I(N__8767));
    InMux I__1405 (
            .O(N__8790),
            .I(N__8755));
    InMux I__1404 (
            .O(N__8789),
            .I(N__8755));
    InMux I__1403 (
            .O(N__8788),
            .I(N__8746));
    InMux I__1402 (
            .O(N__8787),
            .I(N__8746));
    InMux I__1401 (
            .O(N__8786),
            .I(N__8746));
    InMux I__1400 (
            .O(N__8785),
            .I(N__8746));
    CascadeMux I__1399 (
            .O(N__8784),
            .I(N__8743));
    CascadeMux I__1398 (
            .O(N__8783),
            .I(N__8740));
    CascadeMux I__1397 (
            .O(N__8782),
            .I(N__8736));
    LocalMux I__1396 (
            .O(N__8779),
            .I(N__8731));
    LocalMux I__1395 (
            .O(N__8776),
            .I(N__8728));
    CascadeMux I__1394 (
            .O(N__8775),
            .I(N__8723));
    CascadeMux I__1393 (
            .O(N__8774),
            .I(N__8720));
    InMux I__1392 (
            .O(N__8771),
            .I(N__8710));
    InMux I__1391 (
            .O(N__8770),
            .I(N__8710));
    InMux I__1390 (
            .O(N__8767),
            .I(N__8710));
    InMux I__1389 (
            .O(N__8766),
            .I(N__8710));
    InMux I__1388 (
            .O(N__8765),
            .I(N__8701));
    InMux I__1387 (
            .O(N__8764),
            .I(N__8701));
    InMux I__1386 (
            .O(N__8763),
            .I(N__8701));
    InMux I__1385 (
            .O(N__8762),
            .I(N__8701));
    InMux I__1384 (
            .O(N__8761),
            .I(N__8683));
    InMux I__1383 (
            .O(N__8760),
            .I(N__8683));
    LocalMux I__1382 (
            .O(N__8755),
            .I(N__8680));
    LocalMux I__1381 (
            .O(N__8746),
            .I(N__8677));
    InMux I__1380 (
            .O(N__8743),
            .I(N__8668));
    InMux I__1379 (
            .O(N__8740),
            .I(N__8668));
    InMux I__1378 (
            .O(N__8739),
            .I(N__8668));
    InMux I__1377 (
            .O(N__8736),
            .I(N__8668));
    InMux I__1376 (
            .O(N__8735),
            .I(N__8663));
    InMux I__1375 (
            .O(N__8734),
            .I(N__8663));
    Span4Mux_h I__1374 (
            .O(N__8731),
            .I(N__8658));
    Span4Mux_h I__1373 (
            .O(N__8728),
            .I(N__8658));
    InMux I__1372 (
            .O(N__8727),
            .I(N__8647));
    InMux I__1371 (
            .O(N__8726),
            .I(N__8647));
    InMux I__1370 (
            .O(N__8723),
            .I(N__8647));
    InMux I__1369 (
            .O(N__8720),
            .I(N__8647));
    InMux I__1368 (
            .O(N__8719),
            .I(N__8647));
    LocalMux I__1367 (
            .O(N__8710),
            .I(N__8642));
    LocalMux I__1366 (
            .O(N__8701),
            .I(N__8642));
    InMux I__1365 (
            .O(N__8700),
            .I(N__8639));
    InMux I__1364 (
            .O(N__8699),
            .I(N__8624));
    InMux I__1363 (
            .O(N__8698),
            .I(N__8624));
    InMux I__1362 (
            .O(N__8697),
            .I(N__8624));
    InMux I__1361 (
            .O(N__8696),
            .I(N__8624));
    InMux I__1360 (
            .O(N__8695),
            .I(N__8624));
    InMux I__1359 (
            .O(N__8694),
            .I(N__8624));
    InMux I__1358 (
            .O(N__8693),
            .I(N__8624));
    InMux I__1357 (
            .O(N__8692),
            .I(N__8613));
    InMux I__1356 (
            .O(N__8691),
            .I(N__8613));
    InMux I__1355 (
            .O(N__8690),
            .I(N__8613));
    InMux I__1354 (
            .O(N__8689),
            .I(N__8613));
    InMux I__1353 (
            .O(N__8688),
            .I(N__8613));
    LocalMux I__1352 (
            .O(N__8683),
            .I(N__8610));
    Odrv4 I__1351 (
            .O(N__8680),
            .I(un4_pixel_N_3));
    Odrv4 I__1350 (
            .O(N__8677),
            .I(un4_pixel_N_3));
    LocalMux I__1349 (
            .O(N__8668),
            .I(un4_pixel_N_3));
    LocalMux I__1348 (
            .O(N__8663),
            .I(un4_pixel_N_3));
    Odrv4 I__1347 (
            .O(N__8658),
            .I(un4_pixel_N_3));
    LocalMux I__1346 (
            .O(N__8647),
            .I(un4_pixel_N_3));
    Odrv4 I__1345 (
            .O(N__8642),
            .I(un4_pixel_N_3));
    LocalMux I__1344 (
            .O(N__8639),
            .I(un4_pixel_N_3));
    LocalMux I__1343 (
            .O(N__8624),
            .I(un4_pixel_N_3));
    LocalMux I__1342 (
            .O(N__8613),
            .I(un4_pixel_N_3));
    Odrv4 I__1341 (
            .O(N__8610),
            .I(un4_pixel_N_3));
    CascadeMux I__1340 (
            .O(N__8587),
            .I(Pixel_1_RNOZ0Z_73_cascade_));
    InMux I__1339 (
            .O(N__8584),
            .I(N__8581));
    LocalMux I__1338 (
            .O(N__8581),
            .I(Pixel_1_RNOZ0Z_72));
    CascadeMux I__1337 (
            .O(N__8578),
            .I(N__8564));
    InMux I__1336 (
            .O(N__8577),
            .I(N__8556));
    InMux I__1335 (
            .O(N__8576),
            .I(N__8556));
    CascadeMux I__1334 (
            .O(N__8575),
            .I(N__8553));
    InMux I__1333 (
            .O(N__8574),
            .I(N__8549));
    InMux I__1332 (
            .O(N__8573),
            .I(N__8544));
    InMux I__1331 (
            .O(N__8572),
            .I(N__8544));
    InMux I__1330 (
            .O(N__8571),
            .I(N__8541));
    InMux I__1329 (
            .O(N__8570),
            .I(N__8536));
    InMux I__1328 (
            .O(N__8569),
            .I(N__8536));
    InMux I__1327 (
            .O(N__8568),
            .I(N__8533));
    InMux I__1326 (
            .O(N__8567),
            .I(N__8528));
    InMux I__1325 (
            .O(N__8564),
            .I(N__8528));
    InMux I__1324 (
            .O(N__8563),
            .I(N__8523));
    InMux I__1323 (
            .O(N__8562),
            .I(N__8518));
    InMux I__1322 (
            .O(N__8561),
            .I(N__8518));
    LocalMux I__1321 (
            .O(N__8556),
            .I(N__8511));
    InMux I__1320 (
            .O(N__8553),
            .I(N__8505));
    InMux I__1319 (
            .O(N__8552),
            .I(N__8505));
    LocalMux I__1318 (
            .O(N__8549),
            .I(N__8502));
    LocalMux I__1317 (
            .O(N__8544),
            .I(N__8491));
    LocalMux I__1316 (
            .O(N__8541),
            .I(N__8491));
    LocalMux I__1315 (
            .O(N__8536),
            .I(N__8491));
    LocalMux I__1314 (
            .O(N__8533),
            .I(N__8491));
    LocalMux I__1313 (
            .O(N__8528),
            .I(N__8491));
    InMux I__1312 (
            .O(N__8527),
            .I(N__8486));
    InMux I__1311 (
            .O(N__8526),
            .I(N__8486));
    LocalMux I__1310 (
            .O(N__8523),
            .I(N__8481));
    LocalMux I__1309 (
            .O(N__8518),
            .I(N__8481));
    InMux I__1308 (
            .O(N__8517),
            .I(N__8476));
    InMux I__1307 (
            .O(N__8516),
            .I(N__8476));
    InMux I__1306 (
            .O(N__8515),
            .I(N__8471));
    InMux I__1305 (
            .O(N__8514),
            .I(N__8471));
    Span4Mux_v I__1304 (
            .O(N__8511),
            .I(N__8468));
    InMux I__1303 (
            .O(N__8510),
            .I(N__8465));
    LocalMux I__1302 (
            .O(N__8505),
            .I(N__8462));
    Span4Mux_h I__1301 (
            .O(N__8502),
            .I(N__8455));
    Span4Mux_v I__1300 (
            .O(N__8491),
            .I(N__8455));
    LocalMux I__1299 (
            .O(N__8486),
            .I(N__8455));
    Span4Mux_v I__1298 (
            .O(N__8481),
            .I(N__8448));
    LocalMux I__1297 (
            .O(N__8476),
            .I(N__8448));
    LocalMux I__1296 (
            .O(N__8471),
            .I(N__8448));
    Span4Mux_v I__1295 (
            .O(N__8468),
            .I(N__8443));
    LocalMux I__1294 (
            .O(N__8465),
            .I(N__8443));
    Span4Mux_h I__1293 (
            .O(N__8462),
            .I(N__8440));
    Span4Mux_h I__1292 (
            .O(N__8455),
            .I(N__8437));
    Span4Mux_h I__1291 (
            .O(N__8448),
            .I(N__8434));
    Odrv4 I__1290 (
            .O(N__8443),
            .I(font_un36_pixel_23));
    Odrv4 I__1289 (
            .O(N__8440),
            .I(font_un36_pixel_23));
    Odrv4 I__1288 (
            .O(N__8437),
            .I(font_un36_pixel_23));
    Odrv4 I__1287 (
            .O(N__8434),
            .I(font_un36_pixel_23));
    CascadeMux I__1286 (
            .O(N__8425),
            .I(Pixel_1_RNOZ0Z_48_cascade_));
    InMux I__1285 (
            .O(N__8422),
            .I(N__8419));
    LocalMux I__1284 (
            .O(N__8419),
            .I(N_234_0_0));
    InMux I__1283 (
            .O(N__8416),
            .I(N__8413));
    LocalMux I__1282 (
            .O(N__8413),
            .I(N__8410));
    Span4Mux_h I__1281 (
            .O(N__8410),
            .I(N__8407));
    Odrv4 I__1280 (
            .O(N__8407),
            .I(d_N_3_0_0));
    InMux I__1279 (
            .O(N__8404),
            .I(N__8398));
    InMux I__1278 (
            .O(N__8403),
            .I(N__8398));
    LocalMux I__1277 (
            .O(N__8398),
            .I(un7_pixel_0_axb3_i));
    InMux I__1276 (
            .O(N__8395),
            .I(N__8392));
    LocalMux I__1275 (
            .O(N__8392),
            .I(N_326_0_0));
    InMux I__1274 (
            .O(N__8389),
            .I(N__8386));
    LocalMux I__1273 (
            .O(N__8386),
            .I(g0_18_1));
    CascadeMux I__1272 (
            .O(N__8383),
            .I(N_321_0_cascade_));
    InMux I__1271 (
            .O(N__8380),
            .I(N__8377));
    LocalMux I__1270 (
            .O(N__8377),
            .I(N_314_0_0_0));
    InMux I__1269 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__1268 (
            .O(N__8371),
            .I(N__8368));
    Odrv4 I__1267 (
            .O(N__8368),
            .I(N_328_0_0_0));
    CascadeMux I__1266 (
            .O(N__8365),
            .I(g1_2_0_0_cascade_));
    InMux I__1265 (
            .O(N__8362),
            .I(N__8359));
    LocalMux I__1264 (
            .O(N__8359),
            .I(N__8354));
    InMux I__1263 (
            .O(N__8358),
            .I(N__8351));
    InMux I__1262 (
            .O(N__8357),
            .I(N__8348));
    Odrv4 I__1261 (
            .O(N__8354),
            .I(N_192_0_1));
    LocalMux I__1260 (
            .O(N__8351),
            .I(N_192_0_1));
    LocalMux I__1259 (
            .O(N__8348),
            .I(N_192_0_1));
    CascadeMux I__1258 (
            .O(N__8341),
            .I(un117_pixel_6_1_0_1_4_cascade_));
    InMux I__1257 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__1256 (
            .O(N__8335),
            .I(N_219_0_0_1));
    InMux I__1255 (
            .O(N__8332),
            .I(N__8326));
    InMux I__1254 (
            .O(N__8331),
            .I(N__8326));
    LocalMux I__1253 (
            .O(N__8326),
            .I(un7_pixel_1_axb3_i));
    CascadeMux I__1252 (
            .O(N__8323),
            .I(N__8320));
    InMux I__1251 (
            .O(N__8320),
            .I(N__8317));
    LocalMux I__1250 (
            .O(N__8317),
            .I(N__8314));
    Odrv4 I__1249 (
            .O(N__8314),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__1248 (
            .O(N__8311),
            .I(un4_pixel_if_generate_plus_mult1_un61_sum_cry_1));
    CascadeMux I__1247 (
            .O(N__8308),
            .I(N_1482_0_cascade_));
    CascadeMux I__1246 (
            .O(N__8305),
            .I(N__8302));
    InMux I__1245 (
            .O(N__8302),
            .I(N__8299));
    LocalMux I__1244 (
            .O(N__8299),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    InMux I__1243 (
            .O(N__8296),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__1242 (
            .O(N__8293),
            .I(N__8290));
    InMux I__1241 (
            .O(N__8290),
            .I(N__8287));
    LocalMux I__1240 (
            .O(N__8287),
            .I(N__8284));
    Odrv4 I__1239 (
            .O(N__8284),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    InMux I__1238 (
            .O(N__8281),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1237 (
            .O(N__8278),
            .I(N__8275));
    LocalMux I__1236 (
            .O(N__8275),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__1235 (
            .O(N__8272),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__1234 (
            .O(N__8269),
            .I(un4_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1233 (
            .O(N__8266),
            .I(un7_pixel_1_axb2_cascade_));
    InMux I__1232 (
            .O(N__8263),
            .I(N__8257));
    InMux I__1231 (
            .O(N__8262),
            .I(N__8257));
    LocalMux I__1230 (
            .O(N__8257),
            .I(un7_pixel_1_axb2_i));
    InMux I__1229 (
            .O(N__8254),
            .I(N__8251));
    LocalMux I__1228 (
            .O(N__8251),
            .I(Pixel_1_RNOZ0Z_44));
    CascadeMux I__1227 (
            .O(N__8248),
            .I(N_305_0_cascade_));
    CascadeMux I__1226 (
            .O(N__8245),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_));
    InMux I__1225 (
            .O(N__8242),
            .I(N__8239));
    LocalMux I__1224 (
            .O(N__8239),
            .I(Pixel_1_RNOZ0Z_82));
    CascadeMux I__1223 (
            .O(N__8236),
            .I(font_un127_pixel_m_4_1_1_cascade_));
    InMux I__1222 (
            .O(N__8233),
            .I(N__8230));
    LocalMux I__1221 (
            .O(N__8230),
            .I(font_un127_pixel_m_4_1));
    CascadeMux I__1220 (
            .O(N__8227),
            .I(un7_pixel_1_c4_cascade_));
    InMux I__1219 (
            .O(N__8224),
            .I(N__8221));
    LocalMux I__1218 (
            .O(N__8221),
            .I(N__8218));
    Odrv4 I__1217 (
            .O(N__8218),
            .I(font_un127_pixel_m_7_1_0));
    InMux I__1216 (
            .O(N__8215),
            .I(N__8212));
    LocalMux I__1215 (
            .O(N__8212),
            .I(N__8209));
    Odrv4 I__1214 (
            .O(N__8209),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_i));
    InMux I__1213 (
            .O(N__8206),
            .I(N__8202));
    CascadeMux I__1212 (
            .O(N__8205),
            .I(N__8199));
    LocalMux I__1211 (
            .O(N__8202),
            .I(N__8192));
    InMux I__1210 (
            .O(N__8199),
            .I(N__8189));
    InMux I__1209 (
            .O(N__8198),
            .I(N__8186));
    InMux I__1208 (
            .O(N__8197),
            .I(N__8183));
    InMux I__1207 (
            .O(N__8196),
            .I(N__8178));
    InMux I__1206 (
            .O(N__8195),
            .I(N__8178));
    Odrv4 I__1205 (
            .O(N__8192),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2));
    LocalMux I__1204 (
            .O(N__8189),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2));
    LocalMux I__1203 (
            .O(N__8186),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2));
    LocalMux I__1202 (
            .O(N__8183),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2));
    LocalMux I__1201 (
            .O(N__8178),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2));
    InMux I__1200 (
            .O(N__8167),
            .I(N__8164));
    LocalMux I__1199 (
            .O(N__8164),
            .I(N__8161));
    Span4Mux_h I__1198 (
            .O(N__8161),
            .I(N__8158));
    Odrv4 I__1197 (
            .O(N__8158),
            .I(N_307_0_0_1));
    CascadeMux I__1196 (
            .O(N__8155),
            .I(font_un13_pixel_0_1_0_0_22_cascade_));
    InMux I__1195 (
            .O(N__8152),
            .I(N__8148));
    InMux I__1194 (
            .O(N__8151),
            .I(N__8145));
    LocalMux I__1193 (
            .O(N__8148),
            .I(N__8142));
    LocalMux I__1192 (
            .O(N__8145),
            .I(beamY_RNIVV787O2Z0Z_2));
    Odrv4 I__1191 (
            .O(N__8142),
            .I(beamY_RNIVV787O2Z0Z_2));
    InMux I__1190 (
            .O(N__8137),
            .I(N__8134));
    LocalMux I__1189 (
            .O(N__8134),
            .I(N__8131));
    Odrv4 I__1188 (
            .O(N__8131),
            .I(Pixel_1_RNOZ0Z_47));
    CascadeMux I__1187 (
            .O(N__8128),
            .I(N__8125));
    InMux I__1186 (
            .O(N__8125),
            .I(N__8122));
    LocalMux I__1185 (
            .O(N__8122),
            .I(N_338_0_0_0));
    CascadeMux I__1184 (
            .O(N__8119),
            .I(font_un127_pixel_m_cascade_));
    IoInMux I__1183 (
            .O(N__8116),
            .I(N__8113));
    LocalMux I__1182 (
            .O(N__8113),
            .I(N__8110));
    IoSpan4Mux I__1181 (
            .O(N__8110),
            .I(N__8106));
    IoInMux I__1180 (
            .O(N__8109),
            .I(N__8103));
    Span4Mux_s0_v I__1179 (
            .O(N__8106),
            .I(N__8100));
    LocalMux I__1178 (
            .O(N__8103),
            .I(N__8097));
    Span4Mux_v I__1177 (
            .O(N__8100),
            .I(N__8094));
    Span4Mux_s3_v I__1176 (
            .O(N__8097),
            .I(N__8091));
    Span4Mux_v I__1175 (
            .O(N__8094),
            .I(N__8085));
    Span4Mux_v I__1174 (
            .O(N__8091),
            .I(N__8085));
    InMux I__1173 (
            .O(N__8090),
            .I(N__8082));
    Odrv4 I__1172 (
            .O(N__8085),
            .I(Pixel_c));
    LocalMux I__1171 (
            .O(N__8082),
            .I(Pixel_c));
    InMux I__1170 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__1169 (
            .O(N__8074),
            .I(font_un127_pixel_m_4));
    CascadeMux I__1168 (
            .O(N__8071),
            .I(g0_0_1_cascade_));
    InMux I__1167 (
            .O(N__8068),
            .I(N__8065));
    LocalMux I__1166 (
            .O(N__8065),
            .I(N__8062));
    Span4Mux_h I__1165 (
            .O(N__8062),
            .I(N__8059));
    Odrv4 I__1164 (
            .O(N__8059),
            .I(font_un69_pixellto3));
    InMux I__1163 (
            .O(N__8056),
            .I(N__8053));
    LocalMux I__1162 (
            .O(N__8053),
            .I(g0_0_2));
    InMux I__1161 (
            .O(N__8050),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__1160 (
            .O(N__8047),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__1159 (
            .O(N__8044),
            .I(N__8040));
    CascadeMux I__1158 (
            .O(N__8043),
            .I(N__8037));
    InMux I__1157 (
            .O(N__8040),
            .I(N__8032));
    InMux I__1156 (
            .O(N__8037),
            .I(N__8032));
    LocalMux I__1155 (
            .O(N__8032),
            .I(font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5));
    InMux I__1154 (
            .O(N__8029),
            .I(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1153 (
            .O(N__8026),
            .I(N__8023));
    LocalMux I__1152 (
            .O(N__8023),
            .I(N__8019));
    InMux I__1151 (
            .O(N__8022),
            .I(N__8016));
    Odrv12 I__1150 (
            .O(N__8019),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    LocalMux I__1149 (
            .O(N__8016),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    CascadeMux I__1148 (
            .O(N__8011),
            .I(N__8008));
    InMux I__1147 (
            .O(N__8008),
            .I(N__8005));
    LocalMux I__1146 (
            .O(N__8005),
            .I(N__8002));
    Span4Mux_v I__1145 (
            .O(N__8002),
            .I(N__7999));
    Odrv4 I__1144 (
            .O(N__7999),
            .I(beamY_fastZ0Z_8));
    InMux I__1143 (
            .O(N__7996),
            .I(N__7992));
    InMux I__1142 (
            .O(N__7995),
            .I(N__7989));
    LocalMux I__1141 (
            .O(N__7992),
            .I(N__7986));
    LocalMux I__1140 (
            .O(N__7989),
            .I(beamY_fast_RNIG57DZ0Z_8));
    Odrv4 I__1139 (
            .O(N__7986),
            .I(beamY_fast_RNIG57DZ0Z_8));
    CascadeMux I__1138 (
            .O(N__7981),
            .I(beamY_fast_RNIG57DZ0Z_8_cascade_));
    InMux I__1137 (
            .O(N__7978),
            .I(N__7975));
    LocalMux I__1136 (
            .O(N__7975),
            .I(N__7969));
    InMux I__1135 (
            .O(N__7974),
            .I(N__7966));
    InMux I__1134 (
            .O(N__7973),
            .I(N__7961));
    InMux I__1133 (
            .O(N__7972),
            .I(N__7961));
    Odrv4 I__1132 (
            .O(N__7969),
            .I(un5_visibley_c6_0_1));
    LocalMux I__1131 (
            .O(N__7966),
            .I(un5_visibley_c6_0_1));
    LocalMux I__1130 (
            .O(N__7961),
            .I(un5_visibley_c6_0_1));
    InMux I__1129 (
            .O(N__7954),
            .I(N__7950));
    InMux I__1128 (
            .O(N__7953),
            .I(N__7947));
    LocalMux I__1127 (
            .O(N__7950),
            .I(N__7944));
    LocalMux I__1126 (
            .O(N__7947),
            .I(N__7941));
    Odrv12 I__1125 (
            .O(N__7944),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    Odrv4 I__1124 (
            .O(N__7941),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    InMux I__1123 (
            .O(N__7936),
            .I(N__7933));
    LocalMux I__1122 (
            .O(N__7933),
            .I(N__7930));
    Span4Mux_v I__1121 (
            .O(N__7930),
            .I(N__7926));
    InMux I__1120 (
            .O(N__7929),
            .I(N__7923));
    Odrv4 I__1119 (
            .O(N__7926),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    LocalMux I__1118 (
            .O(N__7923),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    InMux I__1117 (
            .O(N__7918),
            .I(N__7914));
    InMux I__1116 (
            .O(N__7917),
            .I(N__7911));
    LocalMux I__1115 (
            .O(N__7914),
            .I(N__7908));
    LocalMux I__1114 (
            .O(N__7911),
            .I(N__7905));
    Odrv12 I__1113 (
            .O(N__7908),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    Odrv4 I__1112 (
            .O(N__7905),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    CascadeMux I__1111 (
            .O(N__7900),
            .I(N__7895));
    CascadeMux I__1110 (
            .O(N__7899),
            .I(N__7892));
    InMux I__1109 (
            .O(N__7898),
            .I(N__7885));
    InMux I__1108 (
            .O(N__7895),
            .I(N__7885));
    InMux I__1107 (
            .O(N__7892),
            .I(N__7882));
    InMux I__1106 (
            .O(N__7891),
            .I(N__7876));
    InMux I__1105 (
            .O(N__7890),
            .I(N__7873));
    LocalMux I__1104 (
            .O(N__7885),
            .I(N__7868));
    LocalMux I__1103 (
            .O(N__7882),
            .I(N__7865));
    InMux I__1102 (
            .O(N__7881),
            .I(N__7860));
    InMux I__1101 (
            .O(N__7880),
            .I(N__7860));
    InMux I__1100 (
            .O(N__7879),
            .I(N__7857));
    LocalMux I__1099 (
            .O(N__7876),
            .I(N__7854));
    LocalMux I__1098 (
            .O(N__7873),
            .I(N__7850));
    InMux I__1097 (
            .O(N__7872),
            .I(N__7845));
    InMux I__1096 (
            .O(N__7871),
            .I(N__7845));
    Span4Mux_v I__1095 (
            .O(N__7868),
            .I(N__7842));
    Span4Mux_v I__1094 (
            .O(N__7865),
            .I(N__7837));
    LocalMux I__1093 (
            .O(N__7860),
            .I(N__7837));
    LocalMux I__1092 (
            .O(N__7857),
            .I(N__7832));
    Span4Mux_h I__1091 (
            .O(N__7854),
            .I(N__7832));
    InMux I__1090 (
            .O(N__7853),
            .I(N__7829));
    Odrv12 I__1089 (
            .O(N__7850),
            .I(beamYZ0Z_4));
    LocalMux I__1088 (
            .O(N__7845),
            .I(beamYZ0Z_4));
    Odrv4 I__1087 (
            .O(N__7842),
            .I(beamYZ0Z_4));
    Odrv4 I__1086 (
            .O(N__7837),
            .I(beamYZ0Z_4));
    Odrv4 I__1085 (
            .O(N__7832),
            .I(beamYZ0Z_4));
    LocalMux I__1084 (
            .O(N__7829),
            .I(beamYZ0Z_4));
    InMux I__1083 (
            .O(N__7816),
            .I(N__7812));
    InMux I__1082 (
            .O(N__7815),
            .I(N__7804));
    LocalMux I__1081 (
            .O(N__7812),
            .I(N__7801));
    InMux I__1080 (
            .O(N__7811),
            .I(N__7798));
    InMux I__1079 (
            .O(N__7810),
            .I(N__7795));
    InMux I__1078 (
            .O(N__7809),
            .I(N__7788));
    InMux I__1077 (
            .O(N__7808),
            .I(N__7788));
    InMux I__1076 (
            .O(N__7807),
            .I(N__7788));
    LocalMux I__1075 (
            .O(N__7804),
            .I(N__7779));
    Span4Mux_h I__1074 (
            .O(N__7801),
            .I(N__7779));
    LocalMux I__1073 (
            .O(N__7798),
            .I(N__7772));
    LocalMux I__1072 (
            .O(N__7795),
            .I(N__7772));
    LocalMux I__1071 (
            .O(N__7788),
            .I(N__7772));
    InMux I__1070 (
            .O(N__7787),
            .I(N__7763));
    InMux I__1069 (
            .O(N__7786),
            .I(N__7763));
    InMux I__1068 (
            .O(N__7785),
            .I(N__7763));
    InMux I__1067 (
            .O(N__7784),
            .I(N__7763));
    Odrv4 I__1066 (
            .O(N__7779),
            .I(beamY_RNI9DLCZ0Z_0));
    Odrv12 I__1065 (
            .O(N__7772),
            .I(beamY_RNI9DLCZ0Z_0));
    LocalMux I__1064 (
            .O(N__7763),
            .I(beamY_RNI9DLCZ0Z_0));
    InMux I__1063 (
            .O(N__7756),
            .I(N__7749));
    InMux I__1062 (
            .O(N__7755),
            .I(N__7749));
    CascadeMux I__1061 (
            .O(N__7754),
            .I(N__7746));
    LocalMux I__1060 (
            .O(N__7749),
            .I(N__7743));
    InMux I__1059 (
            .O(N__7746),
            .I(N__7740));
    Odrv12 I__1058 (
            .O(N__7743),
            .I(un21_beamy_cry_3_c_RNIERZ0Z93));
    LocalMux I__1057 (
            .O(N__7740),
            .I(un21_beamy_cry_3_c_RNIERZ0Z93));
    InMux I__1056 (
            .O(N__7735),
            .I(N__7732));
    LocalMux I__1055 (
            .O(N__7732),
            .I(N__7728));
    InMux I__1054 (
            .O(N__7731),
            .I(N__7725));
    Span4Mux_v I__1053 (
            .O(N__7728),
            .I(N__7720));
    LocalMux I__1052 (
            .O(N__7725),
            .I(N__7720));
    Odrv4 I__1051 (
            .O(N__7720),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    InMux I__1050 (
            .O(N__7717),
            .I(N__7714));
    LocalMux I__1049 (
            .O(N__7714),
            .I(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0));
    InMux I__1048 (
            .O(N__7711),
            .I(N__7707));
    InMux I__1047 (
            .O(N__7710),
            .I(N__7704));
    LocalMux I__1046 (
            .O(N__7707),
            .I(beamY_fastZ0Z_7));
    LocalMux I__1045 (
            .O(N__7704),
            .I(beamY_fastZ0Z_7));
    InMux I__1044 (
            .O(N__7699),
            .I(N__7696));
    LocalMux I__1043 (
            .O(N__7696),
            .I(N__7691));
    InMux I__1042 (
            .O(N__7695),
            .I(N__7687));
    InMux I__1041 (
            .O(N__7694),
            .I(N__7684));
    Span4Mux_v I__1040 (
            .O(N__7691),
            .I(N__7681));
    InMux I__1039 (
            .O(N__7690),
            .I(N__7678));
    LocalMux I__1038 (
            .O(N__7687),
            .I(beamY_fastZ0Z_6));
    LocalMux I__1037 (
            .O(N__7684),
            .I(beamY_fastZ0Z_6));
    Odrv4 I__1036 (
            .O(N__7681),
            .I(beamY_fastZ0Z_6));
    LocalMux I__1035 (
            .O(N__7678),
            .I(beamY_fastZ0Z_6));
    InMux I__1034 (
            .O(N__7669),
            .I(N__7666));
    LocalMux I__1033 (
            .O(N__7666),
            .I(N__7663));
    Span4Mux_h I__1032 (
            .O(N__7663),
            .I(N__7658));
    InMux I__1031 (
            .O(N__7662),
            .I(N__7655));
    InMux I__1030 (
            .O(N__7661),
            .I(N__7652));
    Odrv4 I__1029 (
            .O(N__7658),
            .I(beamY_fastZ0Z_5));
    LocalMux I__1028 (
            .O(N__7655),
            .I(beamY_fastZ0Z_5));
    LocalMux I__1027 (
            .O(N__7652),
            .I(beamY_fastZ0Z_5));
    InMux I__1026 (
            .O(N__7645),
            .I(N__7642));
    LocalMux I__1025 (
            .O(N__7642),
            .I(N__7639));
    Odrv4 I__1024 (
            .O(N__7639),
            .I(un11_visibleylto9_4));
    CascadeMux I__1023 (
            .O(N__7636),
            .I(beamY_fast_RNI198KZ0Z_2_cascade_));
    InMux I__1022 (
            .O(N__7633),
            .I(N__7630));
    LocalMux I__1021 (
            .O(N__7630),
            .I(N__7627));
    Odrv4 I__1020 (
            .O(N__7627),
            .I(font_un127_pixel_m_1));
    InMux I__1019 (
            .O(N__7624),
            .I(un21_beamy_cry_6));
    InMux I__1018 (
            .O(N__7621),
            .I(N__7615));
    InMux I__1017 (
            .O(N__7620),
            .I(N__7615));
    LocalMux I__1016 (
            .O(N__7615),
            .I(un21_beamy_cry_7_c_RNIM7EZ0Z3));
    InMux I__1015 (
            .O(N__7612),
            .I(un21_beamy_cry_7));
    InMux I__1014 (
            .O(N__7609),
            .I(bfn_6_4_0_));
    InMux I__1013 (
            .O(N__7606),
            .I(N__7600));
    InMux I__1012 (
            .O(N__7605),
            .I(N__7600));
    LocalMux I__1011 (
            .O(N__7600),
            .I(un21_beamy_cry_8_c_RNIOAFZ0Z3));
    InMux I__1010 (
            .O(N__7597),
            .I(N__7593));
    CascadeMux I__1009 (
            .O(N__7596),
            .I(N__7589));
    LocalMux I__1008 (
            .O(N__7593),
            .I(N__7582));
    InMux I__1007 (
            .O(N__7592),
            .I(N__7579));
    InMux I__1006 (
            .O(N__7589),
            .I(N__7576));
    InMux I__1005 (
            .O(N__7588),
            .I(N__7573));
    InMux I__1004 (
            .O(N__7587),
            .I(N__7568));
    InMux I__1003 (
            .O(N__7586),
            .I(N__7568));
    InMux I__1002 (
            .O(N__7585),
            .I(N__7563));
    Span4Mux_v I__1001 (
            .O(N__7582),
            .I(N__7558));
    LocalMux I__1000 (
            .O(N__7579),
            .I(N__7558));
    LocalMux I__999 (
            .O(N__7576),
            .I(N__7555));
    LocalMux I__998 (
            .O(N__7573),
            .I(N__7550));
    LocalMux I__997 (
            .O(N__7568),
            .I(N__7550));
    CascadeMux I__996 (
            .O(N__7567),
            .I(N__7546));
    InMux I__995 (
            .O(N__7566),
            .I(N__7543));
    LocalMux I__994 (
            .O(N__7563),
            .I(N__7540));
    Span4Mux_v I__993 (
            .O(N__7558),
            .I(N__7537));
    Span4Mux_h I__992 (
            .O(N__7555),
            .I(N__7532));
    Span4Mux_v I__991 (
            .O(N__7550),
            .I(N__7532));
    InMux I__990 (
            .O(N__7549),
            .I(N__7527));
    InMux I__989 (
            .O(N__7546),
            .I(N__7527));
    LocalMux I__988 (
            .O(N__7543),
            .I(beamYZ0Z_3));
    Odrv4 I__987 (
            .O(N__7540),
            .I(beamYZ0Z_3));
    Odrv4 I__986 (
            .O(N__7537),
            .I(beamYZ0Z_3));
    Odrv4 I__985 (
            .O(N__7532),
            .I(beamYZ0Z_3));
    LocalMux I__984 (
            .O(N__7527),
            .I(beamYZ0Z_3));
    CascadeMux I__983 (
            .O(N__7516),
            .I(N__7512));
    InMux I__982 (
            .O(N__7515),
            .I(N__7505));
    InMux I__981 (
            .O(N__7512),
            .I(N__7505));
    InMux I__980 (
            .O(N__7511),
            .I(N__7498));
    InMux I__979 (
            .O(N__7510),
            .I(N__7498));
    LocalMux I__978 (
            .O(N__7505),
            .I(N__7494));
    InMux I__977 (
            .O(N__7504),
            .I(N__7491));
    InMux I__976 (
            .O(N__7503),
            .I(N__7488));
    LocalMux I__975 (
            .O(N__7498),
            .I(N__7483));
    CascadeMux I__974 (
            .O(N__7497),
            .I(N__7479));
    Span4Mux_v I__973 (
            .O(N__7494),
            .I(N__7472));
    LocalMux I__972 (
            .O(N__7491),
            .I(N__7472));
    LocalMux I__971 (
            .O(N__7488),
            .I(N__7472));
    InMux I__970 (
            .O(N__7487),
            .I(N__7467));
    InMux I__969 (
            .O(N__7486),
            .I(N__7467));
    Span4Mux_h I__968 (
            .O(N__7483),
            .I(N__7463));
    InMux I__967 (
            .O(N__7482),
            .I(N__7458));
    InMux I__966 (
            .O(N__7479),
            .I(N__7458));
    Span4Mux_h I__965 (
            .O(N__7472),
            .I(N__7455));
    LocalMux I__964 (
            .O(N__7467),
            .I(N__7452));
    InMux I__963 (
            .O(N__7466),
            .I(N__7449));
    Span4Mux_v I__962 (
            .O(N__7463),
            .I(N__7446));
    LocalMux I__961 (
            .O(N__7458),
            .I(N__7443));
    Span4Mux_v I__960 (
            .O(N__7455),
            .I(N__7438));
    Span4Mux_h I__959 (
            .O(N__7452),
            .I(N__7438));
    LocalMux I__958 (
            .O(N__7449),
            .I(beamYZ0Z_2));
    Odrv4 I__957 (
            .O(N__7446),
            .I(beamYZ0Z_2));
    Odrv4 I__956 (
            .O(N__7443),
            .I(beamYZ0Z_2));
    Odrv4 I__955 (
            .O(N__7438),
            .I(beamYZ0Z_2));
    CascadeMux I__954 (
            .O(N__7429),
            .I(N__7426));
    InMux I__953 (
            .O(N__7426),
            .I(N__7423));
    LocalMux I__952 (
            .O(N__7423),
            .I(un11_visibleylto9_1));
    CascadeMux I__951 (
            .O(N__7420),
            .I(N_309_0_cascade_));
    InMux I__950 (
            .O(N__7417),
            .I(N__7414));
    LocalMux I__949 (
            .O(N__7414),
            .I(N_316_0));
    CascadeMux I__948 (
            .O(N__7411),
            .I(N_323_0_cascade_));
    InMux I__947 (
            .O(N__7408),
            .I(N__7405));
    LocalMux I__946 (
            .O(N__7405),
            .I(N_302_0_0_0));
    InMux I__945 (
            .O(N__7402),
            .I(N__7399));
    LocalMux I__944 (
            .O(N__7399),
            .I(N__7396));
    Span4Mux_v I__943 (
            .O(N__7396),
            .I(N__7393));
    Odrv4 I__942 (
            .O(N__7393),
            .I(N_5_0_0_0));
    InMux I__941 (
            .O(N__7390),
            .I(un21_beamy_cry_1));
    InMux I__940 (
            .O(N__7387),
            .I(un21_beamy_cry_2));
    InMux I__939 (
            .O(N__7384),
            .I(un21_beamy_cry_3));
    InMux I__938 (
            .O(N__7381),
            .I(un21_beamy_cry_4));
    InMux I__937 (
            .O(N__7378),
            .I(un21_beamy_cry_5));
    InMux I__936 (
            .O(N__7375),
            .I(N__7372));
    LocalMux I__935 (
            .O(N__7372),
            .I(g0_40_1));
    InMux I__934 (
            .O(N__7369),
            .I(N__7366));
    LocalMux I__933 (
            .O(N__7366),
            .I(N__7363));
    Odrv12 I__932 (
            .O(N__7363),
            .I(N_206));
    CascadeMux I__931 (
            .O(N__7360),
            .I(g0_6_1_1_cascade_));
    CascadeMux I__930 (
            .O(N__7357),
            .I(g0_6_1_cascade_));
    InMux I__929 (
            .O(N__7354),
            .I(N__7350));
    InMux I__928 (
            .O(N__7353),
            .I(N__7347));
    LocalMux I__927 (
            .O(N__7350),
            .I(N_192_0_0));
    LocalMux I__926 (
            .O(N__7347),
            .I(N_192_0_0));
    CascadeMux I__925 (
            .O(N__7342),
            .I(g1_3_1_cascade_));
    InMux I__924 (
            .O(N__7339),
            .I(N__7336));
    LocalMux I__923 (
            .O(N__7336),
            .I(N__7333));
    Span4Mux_h I__922 (
            .O(N__7333),
            .I(N__7330));
    Odrv4 I__921 (
            .O(N__7330),
            .I(g1_3));
    CascadeMux I__920 (
            .O(N__7327),
            .I(g0_10_1_cascade_));
    InMux I__919 (
            .O(N__7324),
            .I(N__7321));
    LocalMux I__918 (
            .O(N__7321),
            .I(if_generate_plus_mult1_un75_sum_cry_2_s));
    InMux I__917 (
            .O(N__7318),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_cry_1));
    CascadeMux I__916 (
            .O(N__7315),
            .I(N__7312));
    InMux I__915 (
            .O(N__7312),
            .I(N__7309));
    LocalMux I__914 (
            .O(N__7309),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__913 (
            .O(N__7306),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__912 (
            .O(N__7303),
            .I(N__7300));
    LocalMux I__911 (
            .O(N__7300),
            .I(un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__910 (
            .O(N__7297),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__909 (
            .O(N__7294),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__908 (
            .O(N__7291),
            .I(un7_pixel_1_axb1_cascade_));
    CascadeMux I__907 (
            .O(N__7288),
            .I(N_203_0_cascade_));
    InMux I__906 (
            .O(N__7285),
            .I(N__7282));
    LocalMux I__905 (
            .O(N__7282),
            .I(N_268_0));
    InMux I__904 (
            .O(N__7279),
            .I(N__7276));
    LocalMux I__903 (
            .O(N__7276),
            .I(m3_0));
    CascadeMux I__902 (
            .O(N__7273),
            .I(Pixel_1_RNOZ0Z_69_cascade_));
    InMux I__901 (
            .O(N__7270),
            .I(N__7267));
    LocalMux I__900 (
            .O(N__7267),
            .I(Pixel_1_RNOZ0Z_70));
    CascadeMux I__899 (
            .O(N__7264),
            .I(g0_35_1_cascade_));
    InMux I__898 (
            .O(N__7261),
            .I(N__7258));
    LocalMux I__897 (
            .O(N__7258),
            .I(un115_pixel_13_15___m1_e_0Z0Z_1));
    InMux I__896 (
            .O(N__7255),
            .I(N__7252));
    LocalMux I__895 (
            .O(N__7252),
            .I(un115_pixel_13_15__i2_mux));
    InMux I__894 (
            .O(N__7249),
            .I(N__7246));
    LocalMux I__893 (
            .O(N__7246),
            .I(d_N_6_0));
    CascadeMux I__892 (
            .O(N__7243),
            .I(N__7240));
    InMux I__891 (
            .O(N__7240),
            .I(N__7237));
    LocalMux I__890 (
            .O(N__7237),
            .I(N_6));
    InMux I__889 (
            .O(N__7234),
            .I(N__7231));
    LocalMux I__888 (
            .O(N__7231),
            .I(N_5_i_0));
    CascadeMux I__887 (
            .O(N__7228),
            .I(g1_0_0_cascade_));
    CascadeMux I__886 (
            .O(N__7225),
            .I(N_250_0_cascade_));
    InMux I__885 (
            .O(N__7222),
            .I(N__7219));
    LocalMux I__884 (
            .O(N__7219),
            .I(N_266_0));
    CascadeMux I__883 (
            .O(N__7216),
            .I(N_242_0_cascade_));
    InMux I__882 (
            .O(N__7213),
            .I(N__7210));
    LocalMux I__881 (
            .O(N__7210),
            .I(Pixel_1_RNOZ0Z_61));
    InMux I__880 (
            .O(N__7207),
            .I(N__7204));
    LocalMux I__879 (
            .O(N__7204),
            .I(N_282));
    CascadeMux I__878 (
            .O(N__7201),
            .I(font_un127_pixel_1_1_cascade_));
    InMux I__877 (
            .O(N__7198),
            .I(N__7195));
    LocalMux I__876 (
            .O(N__7195),
            .I(N_336_0));
    InMux I__875 (
            .O(N__7192),
            .I(N__7189));
    LocalMux I__874 (
            .O(N__7189),
            .I(un5_beamx_6));
    CascadeMux I__873 (
            .O(N__7186),
            .I(N__7183));
    InMux I__872 (
            .O(N__7183),
            .I(N__7179));
    InMux I__871 (
            .O(N__7182),
            .I(N__7176));
    LocalMux I__870 (
            .O(N__7179),
            .I(un8_beamy_3));
    LocalMux I__869 (
            .O(N__7176),
            .I(un8_beamy_3));
    InMux I__868 (
            .O(N__7171),
            .I(N__7168));
    LocalMux I__867 (
            .O(N__7168),
            .I(g1_1));
    CascadeMux I__866 (
            .O(N__7165),
            .I(N_283_cascade_));
    InMux I__865 (
            .O(N__7162),
            .I(N__7159));
    LocalMux I__864 (
            .O(N__7159),
            .I(N_285));
    InMux I__863 (
            .O(N__7156),
            .I(N__7153));
    LocalMux I__862 (
            .O(N__7153),
            .I(font_un13_pixel_23));
    InMux I__861 (
            .O(N__7150),
            .I(N__7147));
    LocalMux I__860 (
            .O(N__7147),
            .I(font_un73_pixellt7_0));
    CascadeMux I__859 (
            .O(N__7144),
            .I(font_un13_pixel_23_cascade_));
    InMux I__858 (
            .O(N__7141),
            .I(N__7138));
    LocalMux I__857 (
            .O(N__7138),
            .I(Pixel_1_RNOZ0Z_60));
    CascadeMux I__856 (
            .O(N__7135),
            .I(Pixel_1_RNOZ0Z_39_cascade_));
    CascadeMux I__855 (
            .O(N__7132),
            .I(N__7128));
    InMux I__854 (
            .O(N__7131),
            .I(N__7123));
    InMux I__853 (
            .O(N__7128),
            .I(N__7123));
    LocalMux I__852 (
            .O(N__7123),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0));
    InMux I__851 (
            .O(N__7120),
            .I(N__7117));
    LocalMux I__850 (
            .O(N__7117),
            .I(beamY_RNIF8TM3Z0Z_9));
    CascadeMux I__849 (
            .O(N__7114),
            .I(beamY_RNIVD444Z0Z_9_cascade_));
    InMux I__848 (
            .O(N__7111),
            .I(N__7105));
    CascadeMux I__847 (
            .O(N__7110),
            .I(N__7100));
    CascadeMux I__846 (
            .O(N__7109),
            .I(N__7096));
    CascadeMux I__845 (
            .O(N__7108),
            .I(N__7093));
    LocalMux I__844 (
            .O(N__7105),
            .I(N__7090));
    CascadeMux I__843 (
            .O(N__7104),
            .I(N__7087));
    CascadeMux I__842 (
            .O(N__7103),
            .I(N__7083));
    InMux I__841 (
            .O(N__7100),
            .I(N__7080));
    InMux I__840 (
            .O(N__7099),
            .I(N__7073));
    InMux I__839 (
            .O(N__7096),
            .I(N__7073));
    InMux I__838 (
            .O(N__7093),
            .I(N__7073));
    Span4Mux_h I__837 (
            .O(N__7090),
            .I(N__7070));
    InMux I__836 (
            .O(N__7087),
            .I(N__7063));
    InMux I__835 (
            .O(N__7086),
            .I(N__7063));
    InMux I__834 (
            .O(N__7083),
            .I(N__7063));
    LocalMux I__833 (
            .O(N__7080),
            .I(beamY_RNIGBU92Z0Z_9));
    LocalMux I__832 (
            .O(N__7073),
            .I(beamY_RNIGBU92Z0Z_9));
    Odrv4 I__831 (
            .O(N__7070),
            .I(beamY_RNIGBU92Z0Z_9));
    LocalMux I__830 (
            .O(N__7063),
            .I(beamY_RNIGBU92Z0Z_9));
    CascadeMux I__829 (
            .O(N__7054),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_));
    InMux I__828 (
            .O(N__7051),
            .I(N__7048));
    LocalMux I__827 (
            .O(N__7048),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1));
    CascadeMux I__826 (
            .O(N__7045),
            .I(N_7_0_0_0_cascade_));
    CascadeMux I__825 (
            .O(N__7042),
            .I(un8_beamy_3_cascade_));
    InMux I__824 (
            .O(N__7039),
            .I(N__7036));
    LocalMux I__823 (
            .O(N__7036),
            .I(Pixel_1_RNOZ0Z_43));
    CascadeMux I__822 (
            .O(N__7033),
            .I(N__7030));
    InMux I__821 (
            .O(N__7030),
            .I(N__7027));
    LocalMux I__820 (
            .O(N__7027),
            .I(Pixel_1_RNOZ0Z_42));
    InMux I__819 (
            .O(N__7024),
            .I(N__7021));
    LocalMux I__818 (
            .O(N__7021),
            .I(N__7018));
    Odrv4 I__817 (
            .O(N__7018),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2));
    CascadeMux I__816 (
            .O(N__7015),
            .I(beamY_RNI9I1Q6Z0Z_9_cascade_));
    InMux I__815 (
            .O(N__7012),
            .I(N__7000));
    InMux I__814 (
            .O(N__7011),
            .I(N__7000));
    InMux I__813 (
            .O(N__7010),
            .I(N__7000));
    InMux I__812 (
            .O(N__7009),
            .I(N__7000));
    LocalMux I__811 (
            .O(N__7000),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3));
    InMux I__810 (
            .O(N__6997),
            .I(N__6994));
    LocalMux I__809 (
            .O(N__6994),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0));
    InMux I__808 (
            .O(N__6991),
            .I(N__6982));
    InMux I__807 (
            .O(N__6990),
            .I(N__6982));
    InMux I__806 (
            .O(N__6989),
            .I(N__6982));
    LocalMux I__805 (
            .O(N__6982),
            .I(N__6974));
    InMux I__804 (
            .O(N__6981),
            .I(N__6963));
    InMux I__803 (
            .O(N__6980),
            .I(N__6963));
    InMux I__802 (
            .O(N__6979),
            .I(N__6963));
    InMux I__801 (
            .O(N__6978),
            .I(N__6963));
    InMux I__800 (
            .O(N__6977),
            .I(N__6963));
    Odrv4 I__799 (
            .O(N__6974),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1));
    LocalMux I__798 (
            .O(N__6963),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1));
    InMux I__797 (
            .O(N__6958),
            .I(N__6941));
    InMux I__796 (
            .O(N__6957),
            .I(N__6941));
    InMux I__795 (
            .O(N__6956),
            .I(N__6941));
    InMux I__794 (
            .O(N__6955),
            .I(N__6941));
    InMux I__793 (
            .O(N__6954),
            .I(N__6941));
    InMux I__792 (
            .O(N__6953),
            .I(N__6936));
    InMux I__791 (
            .O(N__6952),
            .I(N__6936));
    LocalMux I__790 (
            .O(N__6941),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3));
    LocalMux I__789 (
            .O(N__6936),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3));
    CascadeMux I__788 (
            .O(N__6931),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_));
    InMux I__787 (
            .O(N__6928),
            .I(N__6925));
    LocalMux I__786 (
            .O(N__6925),
            .I(beamY_RNIQQREO1Z0Z_3));
    InMux I__785 (
            .O(N__6922),
            .I(N__6914));
    InMux I__784 (
            .O(N__6921),
            .I(N__6914));
    InMux I__783 (
            .O(N__6920),
            .I(N__6909));
    InMux I__782 (
            .O(N__6919),
            .I(N__6909));
    LocalMux I__781 (
            .O(N__6914),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_c5));
    LocalMux I__780 (
            .O(N__6909),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_c5));
    CascadeMux I__779 (
            .O(N__6904),
            .I(N__6901));
    InMux I__778 (
            .O(N__6901),
            .I(N__6893));
    InMux I__777 (
            .O(N__6900),
            .I(N__6893));
    InMux I__776 (
            .O(N__6899),
            .I(N__6888));
    InMux I__775 (
            .O(N__6898),
            .I(N__6888));
    LocalMux I__774 (
            .O(N__6893),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2));
    LocalMux I__773 (
            .O(N__6888),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2));
    CascadeMux I__772 (
            .O(N__6883),
            .I(N__6878));
    InMux I__771 (
            .O(N__6882),
            .I(N__6875));
    InMux I__770 (
            .O(N__6881),
            .I(N__6870));
    InMux I__769 (
            .O(N__6878),
            .I(N__6870));
    LocalMux I__768 (
            .O(N__6875),
            .I(N__6867));
    LocalMux I__767 (
            .O(N__6870),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1));
    Odrv4 I__766 (
            .O(N__6867),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1));
    InMux I__765 (
            .O(N__6862),
            .I(N__6858));
    InMux I__764 (
            .O(N__6861),
            .I(N__6855));
    LocalMux I__763 (
            .O(N__6858),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6));
    LocalMux I__762 (
            .O(N__6855),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6));
    InMux I__761 (
            .O(N__6850),
            .I(N__6847));
    LocalMux I__760 (
            .O(N__6847),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0));
    InMux I__759 (
            .O(N__6844),
            .I(N__6841));
    LocalMux I__758 (
            .O(N__6841),
            .I(beamY_4_rep1_RNI9H1FZ0Z1));
    InMux I__757 (
            .O(N__6838),
            .I(N__6835));
    LocalMux I__756 (
            .O(N__6835),
            .I(N__6832));
    Odrv4 I__755 (
            .O(N__6832),
            .I(beamY_RNIHS041Z0Z_6));
    CascadeMux I__754 (
            .O(N__6829),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_));
    InMux I__753 (
            .O(N__6826),
            .I(N__6822));
    InMux I__752 (
            .O(N__6825),
            .I(N__6819));
    LocalMux I__751 (
            .O(N__6822),
            .I(beamY_fastZ0Z_4));
    LocalMux I__750 (
            .O(N__6819),
            .I(beamY_fastZ0Z_4));
    CascadeMux I__749 (
            .O(N__6814),
            .I(N__6809));
    CascadeMux I__748 (
            .O(N__6813),
            .I(N__6806));
    CascadeMux I__747 (
            .O(N__6812),
            .I(N__6803));
    InMux I__746 (
            .O(N__6809),
            .I(N__6800));
    InMux I__745 (
            .O(N__6806),
            .I(N__6796));
    InMux I__744 (
            .O(N__6803),
            .I(N__6793));
    LocalMux I__743 (
            .O(N__6800),
            .I(N__6790));
    InMux I__742 (
            .O(N__6799),
            .I(N__6787));
    LocalMux I__741 (
            .O(N__6796),
            .I(beamY_fastZ0Z_9));
    LocalMux I__740 (
            .O(N__6793),
            .I(beamY_fastZ0Z_9));
    Odrv4 I__739 (
            .O(N__6790),
            .I(beamY_fastZ0Z_9));
    LocalMux I__738 (
            .O(N__6787),
            .I(beamY_fastZ0Z_9));
    InMux I__737 (
            .O(N__6778),
            .I(N__6775));
    LocalMux I__736 (
            .O(N__6775),
            .I(beamY_fast_RNICEGAZ0Z_4));
    CascadeMux I__735 (
            .O(N__6772),
            .I(N__6768));
    InMux I__734 (
            .O(N__6771),
            .I(N__6757));
    InMux I__733 (
            .O(N__6768),
            .I(N__6757));
    InMux I__732 (
            .O(N__6767),
            .I(N__6757));
    InMux I__731 (
            .O(N__6766),
            .I(N__6757));
    LocalMux I__730 (
            .O(N__6757),
            .I(font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5));
    CascadeMux I__729 (
            .O(N__6754),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_));
    InMux I__728 (
            .O(N__6751),
            .I(N__6748));
    LocalMux I__727 (
            .O(N__6748),
            .I(N__6741));
    InMux I__726 (
            .O(N__6747),
            .I(N__6736));
    InMux I__725 (
            .O(N__6746),
            .I(N__6736));
    InMux I__724 (
            .O(N__6745),
            .I(N__6731));
    InMux I__723 (
            .O(N__6744),
            .I(N__6731));
    Odrv4 I__722 (
            .O(N__6741),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i));
    LocalMux I__721 (
            .O(N__6736),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i));
    LocalMux I__720 (
            .O(N__6731),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i));
    InMux I__719 (
            .O(N__6724),
            .I(N__6721));
    LocalMux I__718 (
            .O(N__6721),
            .I(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i));
    CascadeMux I__717 (
            .O(N__6718),
            .I(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_));
    InMux I__716 (
            .O(N__6715),
            .I(N__6712));
    LocalMux I__715 (
            .O(N__6712),
            .I(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1));
    CascadeMux I__714 (
            .O(N__6709),
            .I(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_));
    InMux I__713 (
            .O(N__6706),
            .I(N__6703));
    LocalMux I__712 (
            .O(N__6703),
            .I(N_208_0_0_1));
    CascadeMux I__711 (
            .O(N__6700),
            .I(N_1260_0_0_1_cascade_));
    CascadeMux I__710 (
            .O(N__6697),
            .I(Z_decfrac2_1_0_0_0_cascade_));
    CascadeMux I__709 (
            .O(N__6694),
            .I(un115_pixel_3_0_3__N_8_0_0_0_cascade_));
    InMux I__708 (
            .O(N__6691),
            .I(N__6688));
    LocalMux I__707 (
            .O(N__6688),
            .I(un117_pixel_3_1_0_1_4));
    CascadeMux I__706 (
            .O(N__6685),
            .I(m4_cascade_));
    InMux I__705 (
            .O(N__6682),
            .I(N__6679));
    LocalMux I__704 (
            .O(N__6679),
            .I(N__6676));
    Odrv4 I__703 (
            .O(N__6676),
            .I(Pixel_1_RNOZ0Z_88));
    InMux I__702 (
            .O(N__6673),
            .I(N__6670));
    LocalMux I__701 (
            .O(N__6670),
            .I(Pixel_1_RNOZ0Z_63));
    InMux I__700 (
            .O(N__6667),
            .I(N__6664));
    LocalMux I__699 (
            .O(N__6664),
            .I(un115_pixel_2_0_5__N_14));
    InMux I__698 (
            .O(N__6661),
            .I(N__6655));
    InMux I__697 (
            .O(N__6660),
            .I(N__6655));
    LocalMux I__696 (
            .O(N__6655),
            .I(G_370));
    InMux I__695 (
            .O(N__6652),
            .I(un4_pixel_if_generate_plus_mult1_un82_sum_cry_4));
    CascadeMux I__694 (
            .O(N__6649),
            .I(un4_pixel_N_3_cascade_));
    CascadeMux I__693 (
            .O(N__6646),
            .I(N__6643));
    InMux I__692 (
            .O(N__6643),
            .I(N__6640));
    LocalMux I__691 (
            .O(N__6640),
            .I(un4_pixel_if_generate_plus_mult1_un75_sum_iZ0));
    CascadeMux I__690 (
            .O(N__6637),
            .I(g0_3_1_cascade_));
    CascadeMux I__689 (
            .O(N__6634),
            .I(un115_pixel_0_a2_0_cascade_));
    InMux I__688 (
            .O(N__6631),
            .I(N__6628));
    LocalMux I__687 (
            .O(N__6628),
            .I(N_281));
    InMux I__686 (
            .O(N__6625),
            .I(N__6622));
    LocalMux I__685 (
            .O(N__6622),
            .I(N_231));
    InMux I__684 (
            .O(N__6619),
            .I(N__6616));
    LocalMux I__683 (
            .O(N__6616),
            .I(Pixel_1_RNOZ0Z_62));
    InMux I__682 (
            .O(N__6613),
            .I(N__6610));
    LocalMux I__681 (
            .O(N__6610),
            .I(N_275_0));
    CascadeMux I__680 (
            .O(N__6607),
            .I(N__6604));
    InMux I__679 (
            .O(N__6604),
            .I(N__6601));
    LocalMux I__678 (
            .O(N__6601),
            .I(un115_pixel_13_15__m3_a0Z0Z_0));
    CascadeMux I__677 (
            .O(N__6598),
            .I(un115_pixel_13_15__m3_a0Z0Z_0_cascade_));
    InMux I__676 (
            .O(N__6595),
            .I(N__6592));
    LocalMux I__675 (
            .O(N__6592),
            .I(N_215_0));
    CascadeMux I__674 (
            .O(N__6589),
            .I(Pixel_1_RNOZ0Z_66_cascade_));
    InMux I__673 (
            .O(N__6586),
            .I(N__6583));
    LocalMux I__672 (
            .O(N__6583),
            .I(un117_pixel_3_1_3));
    InMux I__671 (
            .O(N__6580),
            .I(N__6576));
    InMux I__670 (
            .O(N__6579),
            .I(N__6573));
    LocalMux I__669 (
            .O(N__6576),
            .I(N_234_0));
    LocalMux I__668 (
            .O(N__6573),
            .I(N_234_0));
    CascadeMux I__667 (
            .O(N__6568),
            .I(m3_0_cascade_));
    CascadeMux I__666 (
            .O(N__6565),
            .I(un115_pixel_2_0_5__N_9_cascade_));
    CascadeMux I__665 (
            .O(N__6562),
            .I(N__6559));
    InMux I__664 (
            .O(N__6559),
            .I(N__6556));
    LocalMux I__663 (
            .O(N__6556),
            .I(N__6553));
    Span4Mux_h I__662 (
            .O(N__6553),
            .I(N__6549));
    InMux I__661 (
            .O(N__6552),
            .I(N__6546));
    Odrv4 I__660 (
            .O(N__6549),
            .I(un4_beamylt6));
    LocalMux I__659 (
            .O(N__6546),
            .I(un4_beamylt6));
    CascadeMux I__658 (
            .O(N__6541),
            .I(un4_beamylt8_0_cascade_));
    InMux I__657 (
            .O(N__6538),
            .I(N__6535));
    LocalMux I__656 (
            .O(N__6535),
            .I(un1_beamylto9_0));
    CascadeMux I__655 (
            .O(N__6532),
            .I(un1_beamylto9_3_cascade_));
    CascadeMux I__654 (
            .O(N__6529),
            .I(un5_beamx_4_cascade_));
    CascadeMux I__653 (
            .O(N__6526),
            .I(un117_pixel_6_ns_1_3_cascade_));
    InMux I__652 (
            .O(N__6523),
            .I(N__6520));
    LocalMux I__651 (
            .O(N__6520),
            .I(N_192_0));
    CascadeMux I__650 (
            .O(N__6517),
            .I(N_192_0_cascade_));
    CascadeMux I__649 (
            .O(N__6514),
            .I(beamY_RNI1G0FH2_0Z0Z_3_cascade_));
    CascadeMux I__648 (
            .O(N__6511),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cascade_));
    CascadeMux I__647 (
            .O(N__6508),
            .I(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_));
    InMux I__646 (
            .O(N__6505),
            .I(N__6502));
    LocalMux I__645 (
            .O(N__6502),
            .I(N__6499));
    Odrv4 I__644 (
            .O(N__6499),
            .I(beamY_RNICCIKUQ_0Z0Z_3));
    InMux I__643 (
            .O(N__6496),
            .I(N__6493));
    LocalMux I__642 (
            .O(N__6493),
            .I(N__6488));
    InMux I__641 (
            .O(N__6492),
            .I(N__6483));
    InMux I__640 (
            .O(N__6491),
            .I(N__6483));
    Span4Mux_v I__639 (
            .O(N__6488),
            .I(N__6476));
    LocalMux I__638 (
            .O(N__6483),
            .I(N__6476));
    InMux I__637 (
            .O(N__6482),
            .I(N__6473));
    InMux I__636 (
            .O(N__6481),
            .I(N__6470));
    Odrv4 I__635 (
            .O(N__6476),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3));
    LocalMux I__634 (
            .O(N__6473),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3));
    LocalMux I__633 (
            .O(N__6470),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3));
    InMux I__632 (
            .O(N__6463),
            .I(N__6460));
    LocalMux I__631 (
            .O(N__6460),
            .I(N__6456));
    InMux I__630 (
            .O(N__6459),
            .I(N__6453));
    Span4Mux_s3_h I__629 (
            .O(N__6456),
            .I(N__6449));
    LocalMux I__628 (
            .O(N__6453),
            .I(N__6446));
    InMux I__627 (
            .O(N__6452),
            .I(N__6443));
    Odrv4 I__626 (
            .O(N__6449),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    Odrv4 I__625 (
            .O(N__6446),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    LocalMux I__624 (
            .O(N__6443),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    InMux I__623 (
            .O(N__6436),
            .I(N__6430));
    InMux I__622 (
            .O(N__6435),
            .I(N__6430));
    LocalMux I__621 (
            .O(N__6430),
            .I(N__6426));
    InMux I__620 (
            .O(N__6429),
            .I(N__6423));
    Odrv4 I__619 (
            .O(N__6426),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__618 (
            .O(N__6423),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_c5));
    InMux I__617 (
            .O(N__6418),
            .I(N__6414));
    InMux I__616 (
            .O(N__6417),
            .I(N__6411));
    LocalMux I__615 (
            .O(N__6414),
            .I(N__6408));
    LocalMux I__614 (
            .O(N__6411),
            .I(N__6402));
    Span4Mux_s3_h I__613 (
            .O(N__6408),
            .I(N__6399));
    InMux I__612 (
            .O(N__6407),
            .I(N__6392));
    InMux I__611 (
            .O(N__6406),
            .I(N__6392));
    InMux I__610 (
            .O(N__6405),
            .I(N__6392));
    Odrv4 I__609 (
            .O(N__6402),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i));
    Odrv4 I__608 (
            .O(N__6399),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i));
    LocalMux I__607 (
            .O(N__6392),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i));
    InMux I__606 (
            .O(N__6385),
            .I(N__6382));
    LocalMux I__605 (
            .O(N__6382),
            .I(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11));
    CascadeMux I__604 (
            .O(N__6379),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_));
    InMux I__603 (
            .O(N__6376),
            .I(N__6373));
    LocalMux I__602 (
            .O(N__6373),
            .I(N__6368));
    InMux I__601 (
            .O(N__6372),
            .I(N__6363));
    InMux I__600 (
            .O(N__6371),
            .I(N__6363));
    Odrv4 I__599 (
            .O(N__6368),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_c4));
    LocalMux I__598 (
            .O(N__6363),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_c4));
    InMux I__597 (
            .O(N__6358),
            .I(N__6355));
    LocalMux I__596 (
            .O(N__6355),
            .I(N__6352));
    Odrv4 I__595 (
            .O(N__6352),
            .I(beamY_RNICCIKUQZ0Z_3));
    InMux I__594 (
            .O(N__6349),
            .I(N__6346));
    LocalMux I__593 (
            .O(N__6346),
            .I(beamY_RNIIDGN6_0Z0Z_7));
    CascadeMux I__592 (
            .O(N__6343),
            .I(beamY_RNIIDGN6Z0Z_7_cascade_));
    CascadeMux I__591 (
            .O(N__6340),
            .I(beamY_RNIPM0M5Z0Z_9_cascade_));
    InMux I__590 (
            .O(N__6337),
            .I(N__6334));
    LocalMux I__589 (
            .O(N__6334),
            .I(beamY_RNIPM0M5_0Z0Z_9));
    CascadeMux I__588 (
            .O(N__6331),
            .I(N__6328));
    InMux I__587 (
            .O(N__6328),
            .I(N__6319));
    InMux I__586 (
            .O(N__6327),
            .I(N__6319));
    InMux I__585 (
            .O(N__6326),
            .I(N__6319));
    LocalMux I__584 (
            .O(N__6319),
            .I(N__6316));
    Odrv4 I__583 (
            .O(N__6316),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5));
    CascadeMux I__582 (
            .O(N__6313),
            .I(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_));
    InMux I__581 (
            .O(N__6310),
            .I(N__6301));
    InMux I__580 (
            .O(N__6309),
            .I(N__6301));
    InMux I__579 (
            .O(N__6308),
            .I(N__6301));
    LocalMux I__578 (
            .O(N__6301),
            .I(N__6298));
    Odrv4 I__577 (
            .O(N__6298),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0));
    CascadeMux I__576 (
            .O(N__6295),
            .I(beamY_RNI1G0FH2Z0Z_3_cascade_));
    InMux I__575 (
            .O(N__6292),
            .I(N__6286));
    InMux I__574 (
            .O(N__6291),
            .I(N__6286));
    LocalMux I__573 (
            .O(N__6286),
            .I(font_un36_pixel_if_generate_plus_mult1_un68_sum_c4));
    CascadeMux I__572 (
            .O(N__6283),
            .I(N__6279));
    InMux I__571 (
            .O(N__6282),
            .I(N__6271));
    InMux I__570 (
            .O(N__6279),
            .I(N__6271));
    InMux I__569 (
            .O(N__6278),
            .I(N__6271));
    LocalMux I__568 (
            .O(N__6271),
            .I(beamY_RNIUAN5CR1Z0Z_3));
    InMux I__567 (
            .O(N__6268),
            .I(N__6262));
    InMux I__566 (
            .O(N__6267),
            .I(N__6262));
    LocalMux I__565 (
            .O(N__6262),
            .I(font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i));
    InMux I__564 (
            .O(N__6259),
            .I(N__6256));
    LocalMux I__563 (
            .O(N__6256),
            .I(beamY_fast_RNIEGGAZ0Z_6));
    InMux I__562 (
            .O(N__6253),
            .I(N__6250));
    LocalMux I__561 (
            .O(N__6250),
            .I(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0));
    CascadeMux I__560 (
            .O(N__6247),
            .I(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_));
    CascadeMux I__559 (
            .O(N__6244),
            .I(beamY_RNIGBU92Z0Z_9_cascade_));
    CascadeMux I__558 (
            .O(N__6241),
            .I(beamY_RNIQ8RJCCZ0Z_3_cascade_));
    InMux I__557 (
            .O(N__6238),
            .I(N__6235));
    LocalMux I__556 (
            .O(N__6235),
            .I(beamY_RNIQ8RJCC_0Z0Z_3));
    InMux I__555 (
            .O(N__6232),
            .I(N__6229));
    LocalMux I__554 (
            .O(N__6229),
            .I(font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9));
    CascadeMux I__553 (
            .O(N__6226),
            .I(font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_));
    InMux I__552 (
            .O(N__6223),
            .I(N__6220));
    LocalMux I__551 (
            .O(N__6220),
            .I(beamY_RNI03RTE5Z0Z_4));
    InMux I__550 (
            .O(N__6217),
            .I(N__6214));
    LocalMux I__549 (
            .O(N__6214),
            .I(beamY_RNI03RTE5_0Z0Z_4));
    InMux I__548 (
            .O(N__6211),
            .I(N__6208));
    LocalMux I__547 (
            .O(N__6208),
            .I(font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i));
    InMux I__546 (
            .O(N__6205),
            .I(N__6196));
    InMux I__545 (
            .O(N__6204),
            .I(N__6196));
    InMux I__544 (
            .O(N__6203),
            .I(N__6196));
    LocalMux I__543 (
            .O(N__6196),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1));
    CascadeMux I__542 (
            .O(N__6193),
            .I(Pixel_1_RNOZ0Z_34_cascade_));
    IoInMux I__541 (
            .O(N__6190),
            .I(N__6187));
    LocalMux I__540 (
            .O(N__6187),
            .I(N__6184));
    IoSpan4Mux I__539 (
            .O(N__6184),
            .I(N__6181));
    Odrv4 I__538 (
            .O(N__6181),
            .I(Clock12MHz_c));
    IoInMux I__537 (
            .O(N__6178),
            .I(N__6175));
    LocalMux I__536 (
            .O(N__6175),
            .I(N__6172));
    Span4Mux_s1_h I__535 (
            .O(N__6172),
            .I(N__6169));
    Span4Mux_h I__534 (
            .O(N__6169),
            .I(N__6166));
    Span4Mux_v I__533 (
            .O(N__6166),
            .I(N__6163));
    Odrv4 I__532 (
            .O(N__6163),
            .I(\Clock50MHz.PixelClock ));
    CascadeMux I__531 (
            .O(N__6160),
            .I(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_7_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__6178),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    ICE_GB beamX_RNI5457_0_5 (
            .USERSIGNALTOGLOBALBUFFER(N__13333),
            .GLOBALBUFFEROUTPUT(un3_beamx_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam beamY_RNI03RTE5_4_LC_2_6_0.C_ON=1'b0;
    defparam beamY_RNI03RTE5_4_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI03RTE5_4_LC_2_6_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNI03RTE5_4_LC_2_6_0 (
            .in0(N__6990),
            .in1(N__6327),
            .in2(N__7900),
            .in3(N__6309),
            .lcout(beamY_RNI03RTE5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILAPCPC_3_LC_2_6_1.C_ON=1'b0;
    defparam beamY_RNILAPCPC_3_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNILAPCPC_3_LC_2_6_1.LUT_INIT=16'b1111100111110110;
    LogicCell40 beamY_RNILAPCPC_3_LC_2_6_1 (
            .in0(N__6492),
            .in1(N__6376),
            .in2(N__7596),
            .in3(N__6417),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un75_sum_c5_N_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6IISE5_3_LC_2_6_2.C_ON=1'b0;
    defparam beamY_RNI6IISE5_3_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI6IISE5_3_LC_2_6_2.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI6IISE5_3_LC_2_6_2 (
            .in0(N__6989),
            .in1(N__6308),
            .in2(_gnd_net_),
            .in3(N__6326),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ8RJCC_0_3_LC_2_6_3.C_ON=1'b0;
    defparam beamY_RNIQ8RJCC_0_3_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ8RJCC_0_3_LC_2_6_3.LUT_INIT=16'b0110100100011110;
    LogicCell40 beamY_RNIQ8RJCC_0_3_LC_2_6_3 (
            .in0(N__6491),
            .in1(N__9577),
            .in2(N__6160),
            .in3(N__6459),
            .lcout(beamY_RNIQ8RJCC_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI03RTE5_0_4_LC_2_6_7.C_ON=1'b0;
    defparam beamY_RNI03RTE5_0_4_LC_2_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI03RTE5_0_4_LC_2_6_7.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNI03RTE5_0_4_LC_2_6_7 (
            .in0(N__6310),
            .in1(N__7898),
            .in2(N__6331),
            .in3(N__6991),
            .lcout(beamY_RNI03RTE5_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ8RJCC_3_LC_2_7_0.C_ON=1'b0;
    defparam beamY_RNIQ8RJCC_3_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ8RJCC_3_LC_2_7_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIQ8RJCC_3_LC_2_7_0 (
            .in0(N__6496),
            .in1(N__6463),
            .in2(N__9594),
            .in3(N__6203),
            .lcout(),
            .ltout(beamY_RNIQ8RJCCZ0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFVNMRT_3_LC_2_7_1.C_ON=1'b0;
    defparam beamY_RNIFVNMRT_3_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIFVNMRT_3_LC_2_7_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 beamY_RNIFVNMRT_3_LC_2_7_1 (
            .in0(_gnd_net_),
            .in1(N__6418),
            .in2(N__6241),
            .in3(N__6238),
            .lcout(),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_s_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4J28J12_3_LC_2_7_2.C_ON=1'b0;
    defparam beamY_RNI4J28J12_3_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI4J28J12_3_LC_2_7_2.LUT_INIT=16'b0011110001011010;
    LogicCell40 beamY_RNI4J28J12_3_LC_2_7_2 (
            .in0(N__6552),
            .in1(N__6232),
            .in2(N__6226),
            .in3(N__6211),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un75_sum_axbxc5_1_out_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFA02UM_4_LC_2_7_4.C_ON=1'b0;
    defparam beamY_RNIFA02UM_4_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIFA02UM_4_LC_2_7_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 beamY_RNIFA02UM_4_LC_2_7_4 (
            .in0(N__6223),
            .in1(N__6217),
            .in2(_gnd_net_),
            .in3(N__6435),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un75_sum_c5tt_N_2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_2_7_5.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_2_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_2_7_5.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIHUG2_0_3_LC_2_7_5 (
            .in0(N__7504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7592),
            .lcout(un4_beamylt6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIH479FH_3_LC_2_7_6.C_ON=1'b0;
    defparam beamY_RNIH479FH_3_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIH479FH_3_LC_2_7_6.LUT_INIT=16'b0111000111010100;
    LogicCell40 beamY_RNIH479FH_3_LC_2_7_6 (
            .in0(N__9590),
            .in1(N__6436),
            .in2(N__9664),
            .in3(N__6205),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un68_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUAN5CR1_3_LC_2_7_7.C_ON=1'b0;
    defparam beamY_RNIUAN5CR1_3_LC_2_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIUAN5CR1_3_LC_2_7_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 beamY_RNIUAN5CR1_3_LC_2_7_7 (
            .in0(N__6204),
            .in1(N__6358),
            .in2(_gnd_net_),
            .in3(N__6505),
            .lcout(beamY_RNIUAN5CR1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_34_LC_2_8_1.C_ON=1'b0;
    defparam Pixel_1_RNO_34_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_34_LC_2_8_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 Pixel_1_RNO_34_LC_2_8_1 (
            .in0(N__6268),
            .in1(_gnd_net_),
            .in2(N__6283),
            .in3(N__6292),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_34_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_15_LC_2_8_2.C_ON=1'b0;
    defparam Pixel_1_RNO_15_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_15_LC_2_8_2.LUT_INIT=16'b0110001110011100;
    LogicCell40 Pixel_1_RNO_15_LC_2_8_2 (
            .in0(N__7515),
            .in1(N__7597),
            .in2(N__6193),
            .in3(N__6282),
            .lcout(font_un69_pixellto3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBH9OEE_2_LC_2_8_6.C_ON=1'b0;
    defparam beamY_RNIBH9OEE_2_LC_2_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIBH9OEE_2_LC_2_8_6.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIBH9OEE_2_LC_2_8_6 (
            .in0(N__6291),
            .in1(N__6278),
            .in2(N__7516),
            .in3(N__6267),
            .lcout(font_un36_pixel_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_4_3_0.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_4_3_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 beamY_RNIHUG2_3_LC_4_3_0 (
            .in0(N__7487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7549),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_3_LC_4_3_3.C_ON=1'b0;
    defparam beamY_RNI6125_3_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_3_LC_4_3_3.LUT_INIT=16'b1001010101010101;
    LogicCell40 beamY_RNI6125_3_LC_4_3_3 (
            .in0(N__10474),
            .in1(N__7486),
            .in2(N__7567),
            .in3(N__7891),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIEGGA_6_LC_4_4_4.C_ON=1'b0;
    defparam beamY_fast_RNIEGGA_6_LC_4_4_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIEGGA_6_LC_4_4_4.LUT_INIT=16'b0011001100110111;
    LogicCell40 beamY_fast_RNIEGGA_6_LC_4_4_4 (
            .in0(N__10473),
            .in1(N__10781),
            .in2(N__6814),
            .in3(N__7699),
            .lcout(beamY_fast_RNIEGGAZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNITAOJ_5_LC_4_4_7.C_ON=1'b0;
    defparam beamY_fast_RNITAOJ_5_LC_4_4_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNITAOJ_5_LC_4_4_7.LUT_INIT=16'b0000001110101010;
    LogicCell40 beamY_fast_RNITAOJ_5_LC_4_4_7 (
            .in0(N__6778),
            .in1(N__11007),
            .in2(N__6813),
            .in3(N__7669),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4OJ_8_LC_4_5_0.C_ON=1'b0;
    defparam beamY_RNIN4OJ_8_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4OJ_8_LC_4_5_0.LUT_INIT=16'b0101010111001100;
    LogicCell40 beamY_RNIN4OJ_8_LC_4_5_0 (
            .in0(N__10799),
            .in1(N__6259),
            .in2(_gnd_net_),
            .in3(N__10691),
            .lcout(),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGBU92_9_LC_4_5_1.C_ON=1'b0;
    defparam beamY_RNIGBU92_9_LC_4_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIGBU92_9_LC_4_5_1.LUT_INIT=16'b0000000111111110;
    LogicCell40 beamY_RNIGBU92_9_LC_4_5_1 (
            .in0(N__6253),
            .in1(N__6715),
            .in2(N__6247),
            .in3(N__10887),
            .lcout(beamY_RNIGBU92Z0Z_9),
            .ltout(beamY_RNIGBU92Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIDGN6_0_7_LC_4_5_2.C_ON=1'b0;
    defparam beamY_RNIIDGN6_0_7_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIIDGN6_0_7_LC_4_5_2.LUT_INIT=16'b1001100100001001;
    LogicCell40 beamY_RNIIDGN6_0_7_LC_4_5_2 (
            .in0(N__10733),
            .in1(N__6766),
            .in2(N__6244),
            .in3(N__11791),
            .lcout(beamY_RNIIDGN6_0Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPM0M5_0_9_LC_4_5_3.C_ON=1'b0;
    defparam beamY_RNIPM0M5_0_9_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIPM0M5_0_9_LC_4_5_3.LUT_INIT=16'b0100101100101101;
    LogicCell40 beamY_RNIPM0M5_0_9_LC_4_5_3 (
            .in0(N__11793),
            .in1(N__7086),
            .in2(N__6772),
            .in3(N__11918),
            .lcout(beamY_RNIPM0M5_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIDGN6_7_LC_4_5_4.C_ON=1'b0;
    defparam beamY_RNIIDGN6_7_LC_4_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIIDGN6_7_LC_4_5_4.LUT_INIT=16'b1001111110011001;
    LogicCell40 beamY_RNIIDGN6_7_LC_4_5_4 (
            .in0(N__10734),
            .in1(N__6767),
            .in2(N__7103),
            .in3(N__11792),
            .lcout(),
            .ltout(beamY_RNIIDGN6Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIF0K9E_7_LC_4_5_5.C_ON=1'b0;
    defparam beamY_RNIF0K9E_7_LC_4_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIF0K9E_7_LC_4_5_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 beamY_RNIF0K9E_7_LC_4_5_5 (
            .in0(_gnd_net_),
            .in1(N__6349),
            .in2(N__6343),
            .in3(N__11920),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un47_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPM0M5_9_LC_4_5_6.C_ON=1'b0;
    defparam beamY_RNIPM0M5_9_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIPM0M5_9_LC_4_5_6.LUT_INIT=16'b1100100101101100;
    LogicCell40 beamY_RNIPM0M5_9_LC_4_5_6 (
            .in0(N__11919),
            .in1(N__6771),
            .in2(N__7104),
            .in3(N__11794),
            .lcout(),
            .ltout(beamY_RNIPM0M5Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM948D_7_LC_4_5_7.C_ON=1'b0;
    defparam beamY_RNIM948D_7_LC_4_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIM948D_7_LC_4_5_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNIM948D_7_LC_4_5_7 (
            .in0(_gnd_net_),
            .in1(N__10735),
            .in2(N__6340),
            .in3(N__6337),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPTUH72_3_LC_4_6_0.C_ON=1'b0;
    defparam beamY_RNIPTUH72_3_LC_4_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIPTUH72_3_LC_4_6_0.LUT_INIT=16'b1111111101000000;
    LogicCell40 beamY_RNIPTUH72_3_LC_4_6_0 (
            .in0(N__6746),
            .in1(N__6955),
            .in2(N__9746),
            .in3(N__7009),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII319A3_3_LC_4_6_1.C_ON=1'b0;
    defparam beamY_RNII319A3_3_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNII319A3_3_LC_4_6_1.LUT_INIT=16'b0010101110110010;
    LogicCell40 beamY_RNII319A3_3_LC_4_6_1 (
            .in0(N__9564),
            .in1(N__9736),
            .in2(N__6313),
            .in3(N__6981),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQT00H2_3_LC_4_6_2.C_ON=1'b0;
    defparam beamY_RNIQT00H2_3_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIQT00H2_3_LC_4_6_2.LUT_INIT=16'b0010110000011100;
    LogicCell40 beamY_RNIQT00H2_3_LC_4_6_2 (
            .in0(N__6980),
            .in1(N__6958),
            .in2(N__9749),
            .in3(N__7010),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_ac0_7_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5VCS42_3_LC_4_6_3.C_ON=1'b0;
    defparam beamY_RNI5VCS42_3_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI5VCS42_3_LC_4_6_3.LUT_INIT=16'b1100110010010011;
    LogicCell40 beamY_RNI5VCS42_3_LC_4_6_3 (
            .in0(N__6957),
            .in1(N__6747),
            .in2(N__9750),
            .in3(N__6861),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1G0FH2_3_LC_4_6_4.C_ON=1'b0;
    defparam beamY_RNI1G0FH2_3_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI1G0FH2_3_LC_4_6_4.LUT_INIT=16'b1010010101100101;
    LogicCell40 beamY_RNI1G0FH2_3_LC_4_6_4 (
            .in0(N__6978),
            .in1(N__6956),
            .in2(N__9748),
            .in3(N__6745),
            .lcout(),
            .ltout(beamY_RNI1G0FH2Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIF9EJC4_3_LC_4_6_5.C_ON=1'b0;
    defparam beamY_RNIF9EJC4_3_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIF9EJC4_3_LC_4_6_5.LUT_INIT=16'b0111001011011000;
    LogicCell40 beamY_RNIF9EJC4_3_LC_4_6_5 (
            .in0(N__7012),
            .in1(N__9732),
            .in2(N__6295),
            .in3(N__6979),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1G0FH2_0_3_LC_4_6_6.C_ON=1'b0;
    defparam beamY_RNI1G0FH2_0_3_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI1G0FH2_0_3_LC_4_6_6.LUT_INIT=16'b1001011001010110;
    LogicCell40 beamY_RNI1G0FH2_0_3_LC_4_6_6 (
            .in0(N__6977),
            .in1(N__6954),
            .in2(N__9747),
            .in3(N__6744),
            .lcout(),
            .ltout(beamY_RNI1G0FH2_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRD1F25_3_LC_4_6_7.C_ON=1'b0;
    defparam beamY_RNIRD1F25_3_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIRD1F25_3_LC_4_6_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 beamY_RNIRD1F25_3_LC_4_6_7 (
            .in0(N__7011),
            .in1(_gnd_net_),
            .in2(N__6514),
            .in3(N__6928),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM3H2_3_LC_4_7_0.C_ON=1'b0;
    defparam beamY_RNIM3H2_3_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIM3H2_3_LC_4_7_0.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIM3H2_3_LC_4_7_0 (
            .in0(N__11006),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7587),
            .lcout(un1_beamylto9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_3_LC_4_7_1.C_ON=1'b0;
    defparam beamY_RNIBFP3_3_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_3_LC_4_7_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 beamY_RNIBFP3_3_LC_4_7_1 (
            .in0(N__7586),
            .in1(N__7880),
            .in2(_gnd_net_),
            .in3(N__7503),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum),
            .ltout(un1_beamY_if_generate_plus_mult1_un61_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGM5MH6_3_LC_4_7_2.C_ON=1'b0;
    defparam beamY_RNIGM5MH6_3_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIGM5MH6_3_LC_4_7_2.LUT_INIT=16'b1111000001001101;
    LogicCell40 beamY_RNIGM5MH6_3_LC_4_7_2 (
            .in0(N__9656),
            .in1(N__6724),
            .in2(N__6511),
            .in3(N__6481),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICCIKUQ_0_3_LC_4_7_3.C_ON=1'b0;
    defparam beamY_RNICCIKUQ_0_3_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNICCIKUQ_0_3_LC_4_7_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNICCIKUQ_0_3_LC_4_7_3 (
            .in0(N__6407),
            .in1(N__6372),
            .in2(N__6508),
            .in3(N__6429),
            .lcout(beamY_RNICCIKUQ_0Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIF4A60C_3_LC_4_7_4.C_ON=1'b0;
    defparam beamY_RNIF4A60C_3_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIF4A60C_3_LC_4_7_4.LUT_INIT=16'b1111111100100000;
    LogicCell40 beamY_RNIF4A60C_3_LC_4_7_4 (
            .in0(N__6482),
            .in1(N__6405),
            .in2(N__9565),
            .in3(N__6452),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un61_sum_c5),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un61_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICCIKUQ_3_LC_4_7_5.C_ON=1'b0;
    defparam beamY_RNICCIKUQ_3_LC_4_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNICCIKUQ_3_LC_4_7_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNICCIKUQ_3_LC_4_7_5 (
            .in0(N__6406),
            .in1(N__6385),
            .in2(N__6379),
            .in3(N__6371),
            .lcout(beamY_RNICCIKUQZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_4_LC_4_7_6.C_ON=1'b0;
    defparam beamY_RNI2KA6_4_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_4_LC_4_7_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI2KA6_4_LC_4_7_6 (
            .in0(N__7881),
            .in1(N__10557),
            .in2(N__6562),
            .in3(N__10472),
            .lcout(),
            .ltout(un4_beamylt8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_8_LC_4_7_7.C_ON=1'b0;
    defparam beamY_RNISI4A_8_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_8_LC_4_7_7.LUT_INIT=16'b1010101010101000;
    LogicCell40 beamY_RNISI4A_8_LC_4_7_7 (
            .in0(N__10914),
            .in1(N__11005),
            .in2(N__6541),
            .in3(N__10813),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVGA6_2_LC_4_8_1.C_ON=1'b0;
    defparam beamY_RNIVGA6_2_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIVGA6_2_LC_4_8_1.LUT_INIT=16'b0000010000001100;
    LogicCell40 beamY_RNIVGA6_2_LC_4_8_1 (
            .in0(N__10140),
            .in1(N__6538),
            .in2(N__7899),
            .in3(N__7511),
            .lcout(),
            .ltout(un1_beamylto9_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0DB_8_LC_4_8_2.C_ON=1'b0;
    defparam beamY_RNIJ0DB_8_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0DB_8_LC_4_8_2.LUT_INIT=16'b0000000001000000;
    LogicCell40 beamY_RNIJ0DB_8_LC_4_8_2 (
            .in0(N__10818),
            .in1(N__7182),
            .in2(N__6532),
            .in3(N__10927),
            .lcout(beamY_RNIJ0DBZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEIP3_8_LC_4_8_3.C_ON=1'b0;
    defparam beamY_RNIEIP3_8_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIEIP3_8_LC_4_8_3.LUT_INIT=16'b0000000010001000;
    LogicCell40 beamY_RNIEIP3_8_LC_4_8_3 (
            .in0(N__10139),
            .in1(N__7588),
            .in2(_gnd_net_),
            .in3(N__10817),
            .lcout(),
            .ltout(un5_beamx_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2BJ7_2_LC_4_8_4.C_ON=1'b0;
    defparam beamY_RNI2BJ7_2_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI2BJ7_2_LC_4_8_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 beamY_RNI2BJ7_2_LC_4_8_4 (
            .in0(N__7510),
            .in1(N__11008),
            .in2(N__6529),
            .in3(N__10926),
            .lcout(un5_beamx_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_68_LC_4_8_6.C_ON=1'b0;
    defparam Pixel_1_RNO_68_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_68_LC_4_8_6.LUT_INIT=16'b0001000110111011;
    LogicCell40 Pixel_1_RNO_68_LC_4_8_6 (
            .in0(N__10135),
            .in1(N__6579),
            .in2(_gnd_net_),
            .in3(N__6523),
            .lcout(),
            .ltout(un117_pixel_6_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_43_LC_4_8_7.C_ON=1'b0;
    defparam Pixel_1_RNO_43_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_43_LC_4_8_7.LUT_INIT=16'b1100101001010011;
    LogicCell40 Pixel_1_RNO_43_LC_4_8_7 (
            .in0(N__10138),
            .in1(N__8510),
            .in2(N__6526),
            .in3(N__6595),
            .lcout(Pixel_1_RNOZ0Z_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_i_11_LC_4_9_0.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_i_11_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_i_11_LC_4_9_0.LUT_INIT=16'b0100001000000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_i_11_LC_4_9_0 (
            .in0(N__9276),
            .in1(N__8766),
            .in2(N__9054),
            .in3(N__9481),
            .lcout(N_192_0),
            .ltout(N_192_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_67_LC_4_9_1.C_ON=1'b0;
    defparam Pixel_1_RNO_67_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_67_LC_4_9_1.LUT_INIT=16'b0000010110101111;
    LogicCell40 Pixel_1_RNO_67_LC_4_9_1 (
            .in0(N__10064),
            .in1(_gnd_net_),
            .in2(N__6517),
            .in3(N__6682),
            .lcout(un117_pixel_3_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_i_9_LC_4_9_2.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_i_9_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_i_9_LC_4_9_2.LUT_INIT=16'b0000001010000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_i_9_LC_4_9_2 (
            .in0(N__9278),
            .in1(N__8770),
            .in2(N__9055),
            .in3(N__9482),
            .lcout(N_215_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_66_LC_4_9_3.C_ON=1'b0;
    defparam Pixel_1_RNO_66_LC_4_9_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_66_LC_4_9_3.LUT_INIT=16'b0100000000001000;
    LogicCell40 Pixel_1_RNO_66_LC_4_9_3 (
            .in0(N__9483),
            .in1(N__9039),
            .in2(N__8792),
            .in3(N__9279),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_66_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_42_LC_4_9_4.C_ON=1'b0;
    defparam Pixel_1_RNO_42_LC_4_9_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_42_LC_4_9_4.LUT_INIT=16'b1000000011100110;
    LogicCell40 Pixel_1_RNO_42_LC_4_9_4 (
            .in0(N__10136),
            .in1(N__8552),
            .in2(N__6589),
            .in3(N__6586),
            .lcout(Pixel_1_RNOZ0Z_42),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un117_pixel_3_7_LC_4_9_5.C_ON=1'b0;
    defparam un115_pixel_13_15__un117_pixel_3_7_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un117_pixel_3_7_LC_4_9_5.LUT_INIT=16'b0010100011101011;
    LogicCell40 un115_pixel_13_15__un117_pixel_3_7_LC_4_9_5 (
            .in0(N__6631),
            .in1(N__10137),
            .in2(N__8575),
            .in3(N__6580),
            .lcout(N_282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_0_5_LC_4_9_7.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_0_5_LC_4_9_7.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_0_5_LC_4_9_7.LUT_INIT=16'b0100001010001000;
    LogicCell40 un115_pixel_13_15__un115_pixel_0_5_LC_4_9_7 (
            .in0(N__9480),
            .in1(N__9032),
            .in2(N__8791),
            .in3(N__9277),
            .lcout(N_234_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__m3_0_LC_4_10_0.C_ON=1'b0;
    defparam un115_pixel_13_15__m3_0_LC_4_10_0.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__m3_0_LC_4_10_0.LUT_INIT=16'b0010010000000100;
    LogicCell40 un115_pixel_13_15__m3_0_LC_4_10_0 (
            .in0(N__8762),
            .in1(N__9270),
            .in2(N__9056),
            .in3(N__9493),
            .lcout(m3_0),
            .ltout(m3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_60_LC_4_10_1.C_ON=1'b0;
    defparam Pixel_1_RNO_60_LC_4_10_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_60_LC_4_10_1.LUT_INIT=16'b0011000011111100;
    LogicCell40 Pixel_1_RNO_60_LC_4_10_1 (
            .in0(_gnd_net_),
            .in1(N__10083),
            .in2(N__6568),
            .in3(N__6613),
            .lcout(Pixel_1_RNOZ0Z_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_2_0_5__m8_LC_4_10_2.C_ON=1'b0;
    defparam un115_pixel_2_0_5__m8_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam un115_pixel_2_0_5__m8_LC_4_10_2.LUT_INIT=16'b0110011100000111;
    LogicCell40 un115_pixel_2_0_5__m8_LC_4_10_2 (
            .in0(N__8764),
            .in1(N__9272),
            .in2(N__9058),
            .in3(N__9495),
            .lcout(),
            .ltout(un115_pixel_2_0_5__N_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_64_LC_4_10_3.C_ON=1'b0;
    defparam Pixel_1_RNO_64_LC_4_10_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_64_LC_4_10_3.LUT_INIT=16'b0000010110111011;
    LogicCell40 Pixel_1_RNO_64_LC_4_10_3 (
            .in0(N__10085),
            .in1(N__6625),
            .in2(N__6565),
            .in3(N__8514),
            .lcout(),
            .ltout(g0_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_40_LC_4_10_4.C_ON=1'b0;
    defparam Pixel_1_RNO_40_LC_4_10_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_40_LC_4_10_4.LUT_INIT=16'b0111000001111010;
    LogicCell40 Pixel_1_RNO_40_LC_4_10_4 (
            .in0(N__10084),
            .in1(N__6619),
            .in2(N__6637),
            .in3(N__6673),
            .lcout(d_N_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_53_LC_4_10_5.C_ON=1'b0;
    defparam Pixel_1_RNO_53_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_53_LC_4_10_5.LUT_INIT=16'b1001000100010101;
    LogicCell40 Pixel_1_RNO_53_LC_4_10_5 (
            .in0(N__9496),
            .in1(N__9050),
            .in2(N__9288),
            .in3(N__8765),
            .lcout(font_un73_pixellt7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_0_a2_0_LC_4_10_6.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_0_a2_0_LC_4_10_6.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_0_a2_0_LC_4_10_6.LUT_INIT=16'b0000001010000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_0_a2_0_LC_4_10_6 (
            .in0(N__8763),
            .in1(N__9271),
            .in2(N__9057),
            .in3(N__9494),
            .lcout(),
            .ltout(un115_pixel_0_a2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un117_pixel_2_7_LC_4_10_7.C_ON=1'b0;
    defparam un115_pixel_13_15__un117_pixel_2_7_LC_4_10_7.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un117_pixel_2_7_LC_4_10_7.LUT_INIT=16'b0011000011111100;
    LogicCell40 un115_pixel_13_15__un117_pixel_2_7_LC_4_10_7 (
            .in0(_gnd_net_),
            .in1(N__8515),
            .in2(N__6634),
            .in3(N__6667),
            .lcout(N_281),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_1_0_a2_5_LC_4_11_0.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_1_0_a2_5_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_1_0_a2_5_LC_4_11_0.LUT_INIT=16'b0111000010000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_1_0_a2_5_LC_4_11_0 (
            .in0(N__8697),
            .in1(N__9217),
            .in2(N__9030),
            .in3(N__9488),
            .lcout(N_231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_62_LC_4_11_1.C_ON=1'b0;
    defparam Pixel_1_RNO_62_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_62_LC_4_11_1.LUT_INIT=16'b1011011111101101;
    LogicCell40 Pixel_1_RNO_62_LC_4_11_1 (
            .in0(N__9219),
            .in1(N__8976),
            .in2(N__6607),
            .in3(N__8698),
            .lcout(Pixel_1_RNOZ0Z_62),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_86_LC_4_11_2.C_ON=1'b0;
    defparam Pixel_1_RNO_86_LC_4_11_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_86_LC_4_11_2.LUT_INIT=16'b0101101010000000;
    LogicCell40 Pixel_1_RNO_86_LC_4_11_2 (
            .in0(N__8696),
            .in1(N__9216),
            .in2(N__9029),
            .in3(N__9487),
            .lcout(N_275_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_70_LC_4_11_3.C_ON=1'b0;
    defparam Pixel_1_RNO_70_LC_4_11_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_70_LC_4_11_3.LUT_INIT=16'b0000000010001000;
    LogicCell40 Pixel_1_RNO_70_LC_4_11_3 (
            .in0(N__9486),
            .in1(N__8969),
            .in2(_gnd_net_),
            .in3(N__8695),
            .lcout(Pixel_1_RNOZ0Z_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__m3_a0_0_LC_4_11_4.C_ON=1'b0;
    defparam un115_pixel_13_15__m3_a0_0_LC_4_11_4.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__m3_a0_0_LC_4_11_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 un115_pixel_13_15__m3_a0_0_LC_4_11_4 (
            .in0(_gnd_net_),
            .in1(N__8952),
            .in2(_gnd_net_),
            .in3(N__9484),
            .lcout(un115_pixel_13_15__m3_a0Z0Z_0),
            .ltout(un115_pixel_13_15__m3_a0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_88_LC_4_11_5.C_ON=1'b0;
    defparam Pixel_1_RNO_88_LC_4_11_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_88_LC_4_11_5.LUT_INIT=16'b1010111111011101;
    LogicCell40 Pixel_1_RNO_88_LC_4_11_5 (
            .in0(N__9212),
            .in1(N__8967),
            .in2(N__6598),
            .in3(N__8693),
            .lcout(Pixel_1_RNOZ0Z_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_63_LC_4_11_6.C_ON=1'b0;
    defparam Pixel_1_RNO_63_LC_4_11_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_63_LC_4_11_6.LUT_INIT=16'b1101011101111111;
    LogicCell40 Pixel_1_RNO_63_LC_4_11_6 (
            .in0(N__8699),
            .in1(N__9218),
            .in2(N__9031),
            .in3(N__9489),
            .lcout(Pixel_1_RNOZ0Z_63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_2_0_5__m13_LC_4_11_7.C_ON=1'b0;
    defparam un115_pixel_2_0_5__m13_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam un115_pixel_2_0_5__m13_LC_4_11_7.LUT_INIT=16'b0100101000100010;
    LogicCell40 un115_pixel_2_0_5__m13_LC_4_11_7 (
            .in0(N__9485),
            .in1(N__8968),
            .in2(N__9269),
            .in3(N__8694),
            .lcout(un115_pixel_2_0_5__N_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_1_c_LC_4_12_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_1_c_LC_4_12_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_1_c_LC_4_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_cry_1_c_LC_4_12_0 (
            .in0(_gnd_net_),
            .in1(N__13057),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un82_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_4_12_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_4_12_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_4_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_4_12_1 (
            .in0(_gnd_net_),
            .in1(N__6660),
            .in2(N__6646),
            .in3(N__9176),
            .lcout(G_370),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un82_sum_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_3_c_LC_4_12_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_3_c_LC_4_12_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_3_c_LC_4_12_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_cry_3_c_LC_4_12_2 (
            .in0(_gnd_net_),
            .in1(N__7324),
            .in2(N__9259),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_4_c_LC_4_12_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_4_c_LC_4_12_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_cry_4_c_LC_4_12_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_cry_4_c_LC_4_12_3 (
            .in0(_gnd_net_),
            .in1(N__6661),
            .in2(N__7315),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_s_5_LC_4_12_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_s_5_LC_4_12_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_s_5_LC_4_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_s_5_LC_4_12_4 (
            .in0(_gnd_net_),
            .in1(N__7303),
            .in2(_gnd_net_),
            .in3(N__6652),
            .lcout(un4_pixel_N_3),
            .ltout(un4_pixel_N_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_74_LC_4_12_5.C_ON=1'b0;
    defparam Pixel_1_RNO_74_LC_4_12_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_74_LC_4_12_5.LUT_INIT=16'b0000110100001111;
    LogicCell40 Pixel_1_RNO_74_LC_4_12_5 (
            .in0(N__9024),
            .in1(N__9180),
            .in2(N__6649),
            .in3(N__9491),
            .lcout(N_208_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_i_LC_4_12_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_i_LC_4_12_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_i_LC_4_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_i_LC_4_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14092),
            .lcout(un4_pixel_if_generate_plus_mult1_un75_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__g0_0_LC_4_12_7.C_ON=1'b0;
    defparam un115_pixel_13_15__g0_0_LC_4_12_7.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__g0_0_LC_4_12_7.LUT_INIT=16'b0100001000000000;
    LogicCell40 un115_pixel_13_15__g0_0_LC_4_12_7 (
            .in0(N__9211),
            .in1(N__8700),
            .in2(N__9053),
            .in3(N__9490),
            .lcout(N_192_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_75_LC_4_13_0.C_ON=1'b0;
    defparam Pixel_1_RNO_75_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_75_LC_4_13_0.LUT_INIT=16'b1001010111010100;
    LogicCell40 Pixel_1_RNO_75_LC_4_13_0 (
            .in0(N__10124),
            .in1(N__7375),
            .in2(N__8783),
            .in3(N__9027),
            .lcout(),
            .ltout(N_1260_0_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_49_LC_4_13_1.C_ON=1'b0;
    defparam Pixel_1_RNO_49_LC_4_13_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_49_LC_4_13_1.LUT_INIT=16'b1011100011110000;
    LogicCell40 Pixel_1_RNO_49_LC_4_13_1 (
            .in0(N__6706),
            .in1(N__10126),
            .in2(N__6700),
            .in3(N__8576),
            .lcout(N_307_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_78_LC_4_13_2.C_ON=1'b0;
    defparam Pixel_1_RNO_78_LC_4_13_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_78_LC_4_13_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 Pixel_1_RNO_78_LC_4_13_2 (
            .in0(N__9263),
            .in1(N__9028),
            .in2(N__8784),
            .in3(N__9479),
            .lcout(),
            .ltout(Z_decfrac2_1_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_51_LC_4_13_3.C_ON=1'b0;
    defparam Pixel_1_RNO_51_LC_4_13_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_51_LC_4_13_3.LUT_INIT=16'b0111011111010001;
    LogicCell40 Pixel_1_RNO_51_LC_4_13_3 (
            .in0(N__6691),
            .in1(N__8577),
            .in2(N__6697),
            .in3(N__10127),
            .lcout(N_303_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_3_0_3__g0_0_LC_4_13_4.C_ON=1'b0;
    defparam un115_pixel_3_0_3__g0_0_LC_4_13_4.SEQ_MODE=4'b0000;
    defparam un115_pixel_3_0_3__g0_0_LC_4_13_4.LUT_INIT=16'b0100011010000010;
    LogicCell40 un115_pixel_3_0_3__g0_0_LC_4_13_4 (
            .in0(N__9262),
            .in1(N__9025),
            .in2(N__8782),
            .in3(N__9477),
            .lcout(),
            .ltout(un115_pixel_3_0_3__N_8_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_79_LC_4_13_5.C_ON=1'b0;
    defparam Pixel_1_RNO_79_LC_4_13_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_79_LC_4_13_5.LUT_INIT=16'b0000110000111111;
    LogicCell40 Pixel_1_RNO_79_LC_4_13_5 (
            .in0(_gnd_net_),
            .in1(N__10123),
            .in2(N__6694),
            .in3(N__8357),
            .lcout(un117_pixel_3_1_0_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_3_0_3__m4_LC_4_13_6.C_ON=1'b0;
    defparam un115_pixel_3_0_3__m4_LC_4_13_6.SEQ_MODE=4'b0000;
    defparam un115_pixel_3_0_3__m4_LC_4_13_6.LUT_INIT=16'b0100010000000000;
    LogicCell40 un115_pixel_3_0_3__m4_LC_4_13_6 (
            .in0(N__8739),
            .in1(N__9026),
            .in2(_gnd_net_),
            .in3(N__9478),
            .lcout(),
            .ltout(m4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_59_LC_4_13_7.C_ON=1'b0;
    defparam Pixel_1_RNO_59_LC_4_13_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_59_LC_4_13_7.LUT_INIT=16'b1100111100000011;
    LogicCell40 Pixel_1_RNO_59_LC_4_13_7 (
            .in0(_gnd_net_),
            .in1(N__10125),
            .in2(N__6685),
            .in3(N__7353),
            .lcout(N_316_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_8_LC_5_3_0.C_ON=1'b0;
    defparam beamY_8_LC_5_3_0.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_5_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_8_LC_5_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7620),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13221),
            .ce(N__13274),
            .sr(_gnd_net_));
    defparam beamY_fast_8_LC_5_3_1.C_ON=1'b0;
    defparam beamY_fast_8_LC_5_3_1.SEQ_MODE=4'b1000;
    defparam beamY_fast_8_LC_5_3_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_fast_8_LC_5_3_1 (
            .in0(N__7621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13221),
            .ce(N__13274),
            .sr(_gnd_net_));
    defparam beamY_3_LC_5_3_5.C_ON=1'b0;
    defparam beamY_3_LC_5_3_5.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_5_3_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_3_LC_5_3_5 (
            .in0(_gnd_net_),
            .in1(N__7929),
            .in2(_gnd_net_),
            .in3(N__7810),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13221),
            .ce(N__13274),
            .sr(_gnd_net_));
    defparam beamY_fast_4_LC_5_4_0.C_ON=1'b0;
    defparam beamY_fast_4_LC_5_4_0.SEQ_MODE=4'b1000;
    defparam beamY_fast_4_LC_5_4_0.LUT_INIT=16'b0101000001010000;
    LogicCell40 beamY_fast_4_LC_5_4_0 (
            .in0(N__7808),
            .in1(_gnd_net_),
            .in2(N__7754),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13218),
            .ce(N__13272),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIRPUB_4_LC_5_4_1.C_ON=1'b0;
    defparam beamY_fast_RNIRPUB_4_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIRPUB_4_LC_5_4_1.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_fast_RNIRPUB_4_LC_5_4_1 (
            .in0(N__6799),
            .in1(N__6825),
            .in2(_gnd_net_),
            .in3(N__7662),
            .lcout(),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIT5511_6_LC_5_4_2.C_ON=1'b0;
    defparam beamY_fast_RNIT5511_6_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIT5511_6_LC_5_4_2.LUT_INIT=16'b0010001011110010;
    LogicCell40 beamY_fast_RNIT5511_6_LC_5_4_2 (
            .in0(N__7717),
            .in1(N__10692),
            .in2(N__6718),
            .in3(N__7695),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_9_LC_5_4_3.C_ON=1'b0;
    defparam beamY_fast_9_LC_5_4_3.SEQ_MODE=4'b1000;
    defparam beamY_fast_9_LC_5_4_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_fast_9_LC_5_4_3 (
            .in0(_gnd_net_),
            .in1(N__7606),
            .in2(_gnd_net_),
            .in3(N__7809),
            .lcout(beamY_fastZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13218),
            .ce(N__13272),
            .sr(_gnd_net_));
    defparam beamY_9_LC_5_4_7.C_ON=1'b0;
    defparam beamY_9_LC_5_4_7.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_5_4_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_9_LC_5_4_7 (
            .in0(_gnd_net_),
            .in1(N__7605),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13218),
            .ce(N__13272),
            .sr(_gnd_net_));
    defparam beamY_RNIFIHM2_9_LC_5_5_0.C_ON=1'b0;
    defparam beamY_RNIFIHM2_9_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIFIHM2_9_LC_5_5_0.LUT_INIT=16'b0001010100101010;
    LogicCell40 beamY_RNIFIHM2_9_LC_5_5_0 (
            .in0(N__10885),
            .in1(N__12132),
            .in2(N__11926),
            .in3(N__10363),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC4JRL_9_LC_5_5_1.C_ON=1'b0;
    defparam beamY_RNIC4JRL_9_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIC4JRL_9_LC_5_5_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIC4JRL_9_LC_5_5_1 (
            .in0(N__11797),
            .in1(N__6898),
            .in2(N__6709),
            .in3(N__6919),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNICEGA_4_LC_5_5_2.C_ON=1'b0;
    defparam beamY_fast_RNICEGA_4_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNICEGA_4_LC_5_5_2.LUT_INIT=16'b0000001100010011;
    LogicCell40 beamY_fast_RNICEGA_4_LC_5_5_2 (
            .in0(N__6826),
            .in1(N__10992),
            .in2(N__6812),
            .in3(N__10553),
            .lcout(beamY_fast_RNICEGAZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIF1IR4_9_LC_5_5_3.C_ON=1'b0;
    defparam beamY_RNIF1IR4_9_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIF1IR4_9_LC_5_5_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 beamY_RNIF1IR4_9_LC_5_5_3 (
            .in0(N__11795),
            .in1(N__11924),
            .in2(N__7108),
            .in3(N__12135),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4DUR1_9_LC_5_5_4.C_ON=1'b0;
    defparam beamY_RNI4DUR1_9_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI4DUR1_9_LC_5_5_4.LUT_INIT=16'b1000100001000100;
    LogicCell40 beamY_RNI4DUR1_9_LC_5_5_4 (
            .in0(N__10884),
            .in1(N__12131),
            .in2(_gnd_net_),
            .in3(N__10362),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKOS54_9_LC_5_5_5.C_ON=1'b0;
    defparam beamY_RNIKOS54_9_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIKOS54_9_LC_5_5_5.LUT_INIT=16'b1001011000001111;
    LogicCell40 beamY_RNIKOS54_9_LC_5_5_5 (
            .in0(N__10364),
            .in1(N__10886),
            .in2(N__7109),
            .in3(N__12134),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un47_sum_axbxc5_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIL92Q3_9_LC_5_5_6.C_ON=1'b0;
    defparam beamY_RNIL92Q3_9_LC_5_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIL92Q3_9_LC_5_5_6.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNIL92Q3_9_LC_5_5_6 (
            .in0(N__11925),
            .in1(N__7099),
            .in2(_gnd_net_),
            .in3(N__11796),
            .lcout(),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7L40P_9_LC_5_5_7.C_ON=1'b0;
    defparam beamY_RNI7L40P_9_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI7L40P_9_LC_5_5_7.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNI7L40P_9_LC_5_5_7 (
            .in0(N__6882),
            .in1(N__6899),
            .in2(N__6754),
            .in3(N__6920),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5VCS42_0_3_LC_5_6_0.C_ON=1'b0;
    defparam beamY_RNI5VCS42_0_3_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI5VCS42_0_3_LC_5_6_0.LUT_INIT=16'b0110011001011001;
    LogicCell40 beamY_RNI5VCS42_0_3_LC_5_6_0 (
            .in0(N__6751),
            .in1(N__6953),
            .in2(N__9751),
            .in3(N__6862),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un68_sum_ac0_7_0_N_9_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_4_rep1_RNI9H1F1_LC_5_6_1.C_ON=1'b0;
    defparam beamY_4_rep1_RNI9H1F1_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam beamY_4_rep1_RNI9H1F1_LC_5_6_1.LUT_INIT=16'b0101000001000001;
    LogicCell40 beamY_4_rep1_RNI9H1F1_LC_5_6_1 (
            .in0(N__12145),
            .in1(N__10454),
            .in2(N__10554),
            .in3(N__10596),
            .lcout(beamY_4_rep1_RNI9H1FZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9I1Q6_9_LC_5_6_2.C_ON=1'b0;
    defparam beamY_RNI9I1Q6_9_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI9I1Q6_9_LC_5_6_2.LUT_INIT=16'b1000000000100000;
    LogicCell40 beamY_RNI9I1Q6_9_LC_5_6_2 (
            .in0(N__6850),
            .in1(N__10913),
            .in2(N__7110),
            .in3(N__10365),
            .lcout(),
            .ltout(beamY_RNI9I1Q6Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI035HO_9_LC_5_6_3.C_ON=1'b0;
    defparam beamY_RNI035HO_9_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI035HO_9_LC_5_6_3.LUT_INIT=16'b1111111111111000;
    LogicCell40 beamY_RNI035HO_9_LC_5_6_3 (
            .in0(N__10198),
            .in1(N__7024),
            .in2(N__7015),
            .in3(N__7051),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8L6E21_9_LC_5_6_4.C_ON=1'b0;
    defparam beamY_RNI8L6E21_9_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI8L6E21_9_LC_5_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNI8L6E21_9_LC_5_6_4 (
            .in0(N__6997),
            .in1(N__6881),
            .in2(N__6904),
            .in3(N__6922),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQQREO1_3_LC_5_6_5.C_ON=1'b0;
    defparam beamY_RNIQQREO1_3_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIQQREO1_3_LC_5_6_5.LUT_INIT=16'b0101101010100101;
    LogicCell40 beamY_RNIQQREO1_3_LC_5_6_5 (
            .in0(N__6952),
            .in1(_gnd_net_),
            .in2(N__6931),
            .in3(N__9742),
            .lcout(beamY_RNIQQREO1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHS041_6_LC_5_6_6.C_ON=1'b0;
    defparam beamY_RNIHS041_6_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIHS041_6_LC_5_6_6.LUT_INIT=16'b0000000010011001;
    LogicCell40 beamY_RNIHS041_6_LC_5_6_6 (
            .in0(N__10533),
            .in1(N__10453),
            .in2(_gnd_net_),
            .in3(N__12144),
            .lcout(beamY_RNIHS041Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC4JRL_0_9_LC_5_6_7.C_ON=1'b0;
    defparam beamY_RNIC4JRL_0_9_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIC4JRL_0_9_LC_5_6_7.LUT_INIT=16'b0000000010010110;
    LogicCell40 beamY_RNIC4JRL_0_9_LC_5_6_7 (
            .in0(N__6921),
            .in1(N__6900),
            .in2(N__6883),
            .in3(N__11787),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_5_7_0.C_ON=1'b0;
    defparam beamY_0_LC_5_7_0.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_5_7_0.LUT_INIT=16'b0001000111001100;
    LogicCell40 beamY_0_LC_5_7_0 (
            .in0(N__7815),
            .in1(N__11090),
            .in2(_gnd_net_),
            .in3(N__13294),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13214),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFHKL3_7_LC_5_7_1.C_ON=1'b0;
    defparam beamY_RNIFHKL3_7_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIFHKL3_7_LC_5_7_1.LUT_INIT=16'b0010001000101000;
    LogicCell40 beamY_RNIFHKL3_7_LC_5_7_1 (
            .in0(N__7131),
            .in1(N__10986),
            .in2(N__10285),
            .in3(N__10532),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5D1R2_6_LC_5_7_2.C_ON=1'b0;
    defparam beamY_RNI5D1R2_6_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI5D1R2_6_LC_5_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 beamY_RNI5D1R2_6_LC_5_7_2 (
            .in0(N__6844),
            .in1(N__6838),
            .in2(_gnd_net_),
            .in3(N__10681),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIF8TM3_9_LC_5_7_3.C_ON=1'b0;
    defparam beamY_RNIF8TM3_9_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIF8TM3_9_LC_5_7_3.LUT_INIT=16'b1100000000000000;
    LogicCell40 beamY_RNIF8TM3_9_LC_5_7_3 (
            .in0(_gnd_net_),
            .in1(N__11898),
            .in2(N__6829),
            .in3(N__10911),
            .lcout(beamY_RNIF8TM3Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_4_rep1_RNIQOGL_LC_5_7_4.C_ON=1'b0;
    defparam beamY_4_rep1_RNIQOGL_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam beamY_4_rep1_RNIQOGL_LC_5_7_4.LUT_INIT=16'b1110000110100101;
    LogicCell40 beamY_4_rep1_RNIQOGL_LC_5_7_4 (
            .in0(N__10452),
            .in1(N__10680),
            .in2(N__10552),
            .in3(N__10595),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVD444_9_LC_5_7_5.C_ON=1'b0;
    defparam beamY_RNIVD444_9_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIVD444_9_LC_5_7_5.LUT_INIT=16'b1000000000100000;
    LogicCell40 beamY_RNIVD444_9_LC_5_7_5 (
            .in0(N__11900),
            .in1(N__10912),
            .in2(N__7132),
            .in3(N__7995),
            .lcout(),
            .ltout(beamY_RNIVD444Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9G078_9_LC_5_7_6.C_ON=1'b0;
    defparam beamY_RNI9G078_9_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI9G078_9_LC_5_7_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 beamY_RNI9G078_9_LC_5_7_6 (
            .in0(_gnd_net_),
            .in1(N__7120),
            .in2(N__7114),
            .in3(N__7978),
            .lcout(),
            .ltout(font_un36_pixel_if_generate_plus_mult1_un54_sum_c5_0_a1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUP21C_9_LC_5_7_7.C_ON=1'b0;
    defparam beamY_RNIUP21C_9_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIUP21C_9_LC_5_7_7.LUT_INIT=16'b0111001001010001;
    LogicCell40 beamY_RNIUP21C_9_LC_5_7_7 (
            .in0(N__7111),
            .in1(N__11786),
            .in2(N__7054),
            .in3(N__11899),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_10_LC_5_8_0.C_ON=1'b0;
    defparam Pixel_1_RNO_10_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_10_LC_5_8_0.LUT_INIT=16'b1110001010111000;
    LogicCell40 Pixel_1_RNO_10_LC_5_8_0 (
            .in0(N__7402),
            .in1(N__7171),
            .in2(N__7243),
            .in3(N__11437),
            .lcout(),
            .ltout(N_7_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_3_LC_5_8_1.C_ON=1'b0;
    defparam Pixel_1_RNO_3_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_3_LC_5_8_1.LUT_INIT=16'b1111011010010000;
    LogicCell40 Pixel_1_RNO_3_LC_5_8_1 (
            .in0(N__13075),
            .in1(N__8206),
            .in2(N__7045),
            .in3(N__7198),
            .lcout(N_338_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4H2_6_LC_5_8_2.C_ON=1'b0;
    defparam beamY_RNIN4H2_6_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4H2_6_LC_5_8_2.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIN4H2_6_LC_5_8_2 (
            .in0(N__10545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10458),
            .lcout(un8_beamy_3),
            .ltout(un8_beamy_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISKOB_4_LC_5_8_3.C_ON=1'b0;
    defparam beamY_RNISKOB_4_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam beamY_RNISKOB_4_LC_5_8_3.LUT_INIT=16'b0101000011110000;
    LogicCell40 beamY_RNISKOB_4_LC_5_8_3 (
            .in0(N__10693),
            .in1(_gnd_net_),
            .in2(N__7042),
            .in3(N__7871),
            .lcout(un8_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_26_LC_5_8_4.C_ON=1'b0;
    defparam Pixel_1_RNO_26_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_26_LC_5_8_4.LUT_INIT=16'b0010011101010101;
    LogicCell40 Pixel_1_RNO_26_LC_5_8_4 (
            .in0(N__11088),
            .in1(N__7039),
            .in2(N__7033),
            .in3(N__7156),
            .lcout(),
            .ltout(font_un127_pixel_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_11_LC_5_8_5.C_ON=1'b0;
    defparam Pixel_1_RNO_11_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_11_LC_5_8_5.LUT_INIT=16'b0000111110101100;
    LogicCell40 Pixel_1_RNO_11_LC_5_8_5 (
            .in0(N__7207),
            .in1(N__7162),
            .in2(N__7201),
            .in3(N__7234),
            .lcout(N_336_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_0_LC_5_8_6.C_ON=1'b0;
    defparam beamY_RNI9DLC_0_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_0_LC_5_8_6.LUT_INIT=16'b0000000010000000;
    LogicCell40 beamY_RNI9DLC_0_LC_5_8_6 (
            .in0(N__7872),
            .in1(N__7192),
            .in2(N__7186),
            .in3(N__11089),
            .lcout(beamY_RNI9DLCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_23_LC_5_8_7.C_ON=1'b0;
    defparam Pixel_1_RNO_23_LC_5_8_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_23_LC_5_8_7.LUT_INIT=16'b0101000001010000;
    LogicCell40 Pixel_1_RNO_23_LC_5_8_7 (
            .in0(N__13074),
            .in1(_gnd_net_),
            .in2(N__8205),
            .in3(_gnd_net_),
            .lcout(g1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_41_LC_5_9_0.C_ON=1'b0;
    defparam Pixel_1_RNO_41_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_41_LC_5_9_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 Pixel_1_RNO_41_LC_5_9_0 (
            .in0(N__8562),
            .in1(N__7222),
            .in2(_gnd_net_),
            .in3(N__7369),
            .lcout(),
            .ltout(N_283_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_25_LC_5_9_1.C_ON=1'b0;
    defparam Pixel_1_RNO_25_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_25_LC_5_9_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 Pixel_1_RNO_25_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(N__10095),
            .in2(N__7165),
            .in3(N__8151),
            .lcout(N_285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEQIGK2_LC_5_9_3.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEQIGK2_LC_5_9_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEQIGK2_LC_5_9_3.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEQIGK2_LC_5_9_3 (
            .in0(N__13071),
            .in1(N__11434),
            .in2(_gnd_net_),
            .in3(N__8195),
            .lcout(font_un13_pixel_23),
            .ltout(font_un13_pixel_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_35_LC_5_9_4.C_ON=1'b0;
    defparam Pixel_1_RNO_35_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_35_LC_5_9_4.LUT_INIT=16'b0010000000100010;
    LogicCell40 Pixel_1_RNO_35_LC_5_9_4 (
            .in0(N__7633),
            .in1(N__7150),
            .in2(N__7144),
            .in3(N__8233),
            .lcout(font_un127_pixel_m_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_39_LC_5_9_5.C_ON=1'b0;
    defparam Pixel_1_RNO_39_LC_5_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_39_LC_5_9_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 Pixel_1_RNO_39_LC_5_9_5 (
            .in0(N__7141),
            .in1(N__8561),
            .in2(_gnd_net_),
            .in3(N__7213),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_39_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_22_LC_5_9_6.C_ON=1'b0;
    defparam Pixel_1_RNO_22_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_22_LC_5_9_6.LUT_INIT=16'b0000001111001111;
    LogicCell40 Pixel_1_RNO_22_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(N__11112),
            .in2(N__7135),
            .in3(N__7249),
            .lcout(N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_24_LC_5_9_7.C_ON=1'b0;
    defparam Pixel_1_RNO_24_LC_5_9_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_24_LC_5_9_7.LUT_INIT=16'b1001100111001100;
    LogicCell40 Pixel_1_RNO_24_LC_5_9_7 (
            .in0(N__13072),
            .in1(N__11435),
            .in2(_gnd_net_),
            .in3(N__8196),
            .lcout(N_5_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_45_LC_5_10_0.C_ON=1'b0;
    defparam Pixel_1_RNO_45_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_45_LC_5_10_0.LUT_INIT=16'b0100000000001000;
    LogicCell40 Pixel_1_RNO_45_LC_5_10_0 (
            .in0(N__9446),
            .in1(N__9285),
            .in2(N__9020),
            .in3(N__8788),
            .lcout(),
            .ltout(g1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_28_LC_5_10_1.C_ON=1'b0;
    defparam Pixel_1_RNO_28_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_28_LC_5_10_1.LUT_INIT=16'b1101010110000000;
    LogicCell40 Pixel_1_RNO_28_LC_5_10_1 (
            .in0(N__10087),
            .in1(N__8517),
            .in2(N__7228),
            .in3(N__7339),
            .lcout(N_326_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_5_10_2.C_ON=1'b0;
    defparam beamY_1_LC_5_10_2.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_5_10_2.LUT_INIT=16'b0011011101000000;
    LogicCell40 beamY_1_LC_5_10_2 (
            .in0(N__7811),
            .in1(N__13292),
            .in2(N__11131),
            .in3(N__10088),
            .lcout(un43lto1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13215),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_4_0_1_LC_5_10_3.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_4_0_1_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_4_0_1_LC_5_10_3.LUT_INIT=16'b0001101000000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_4_0_1_LC_5_10_3 (
            .in0(N__8785),
            .in1(N__8942),
            .in2(N__9289),
            .in3(N__9443),
            .lcout(),
            .ltout(N_250_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVV787O2_2_LC_5_10_4.C_ON=1'b0;
    defparam beamY_RNIVV787O2_2_LC_5_10_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIVV787O2_2_LC_5_10_4.LUT_INIT=16'b0000010110101111;
    LogicCell40 beamY_RNIVV787O2_2_LC_5_10_4 (
            .in0(N__8516),
            .in1(_gnd_net_),
            .in2(N__7225),
            .in3(N__7255),
            .lcout(beamY_RNIVV787O2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_1_i_1_LC_5_10_5.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_1_i_1_LC_5_10_5.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_1_i_1_LC_5_10_5.LUT_INIT=16'b0100010000000000;
    LogicCell40 un115_pixel_13_15__un115_pixel_1_i_1_LC_5_10_5 (
            .in0(N__9283),
            .in1(N__8943),
            .in2(_gnd_net_),
            .in3(N__9444),
            .lcout(N_266_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_87_LC_5_10_6.C_ON=1'b0;
    defparam Pixel_1_RNO_87_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_87_LC_5_10_6.LUT_INIT=16'b0110100000101000;
    LogicCell40 Pixel_1_RNO_87_LC_5_10_6 (
            .in0(N__9445),
            .in1(N__9284),
            .in2(N__9019),
            .in3(N__8786),
            .lcout(),
            .ltout(N_242_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_61_LC_5_10_7.C_ON=1'b0;
    defparam Pixel_1_RNO_61_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_61_LC_5_10_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 Pixel_1_RNO_61_LC_5_10_7 (
            .in0(N__8787),
            .in1(_gnd_net_),
            .in2(N__7216),
            .in3(N__10086),
            .lcout(Pixel_1_RNOZ0Z_61),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_69_LC_5_11_0.C_ON=1'b0;
    defparam Pixel_1_RNO_69_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_69_LC_5_11_0.LUT_INIT=16'b0000100011111000;
    LogicCell40 Pixel_1_RNO_69_LC_5_11_0 (
            .in0(N__8727),
            .in1(N__7261),
            .in2(N__10134),
            .in3(N__7279),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_69_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_44_LC_5_11_1.C_ON=1'b0;
    defparam Pixel_1_RNO_44_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_44_LC_5_11_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 Pixel_1_RNO_44_LC_5_11_1 (
            .in0(N__8527),
            .in1(_gnd_net_),
            .in2(N__7273),
            .in3(N__7270),
            .lcout(Pixel_1_RNOZ0Z_44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_1_i_0_LC_5_11_2.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_1_i_0_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_1_i_0_LC_5_11_2.LUT_INIT=16'b0000100010001000;
    LogicCell40 un115_pixel_13_15__un115_pixel_1_i_0_LC_5_11_2 (
            .in0(N__9431),
            .in1(N__8938),
            .in2(N__8775),
            .in3(N__9252),
            .lcout(N_268_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_91_LC_5_11_3.C_ON=1'b0;
    defparam Pixel_1_RNO_91_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_91_LC_5_11_3.LUT_INIT=16'b0010010100101111;
    LogicCell40 Pixel_1_RNO_91_LC_5_11_3 (
            .in0(N__9247),
            .in1(N__8719),
            .in2(N__9017),
            .in3(N__9428),
            .lcout(),
            .ltout(g0_35_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_76_LC_5_11_4.C_ON=1'b0;
    defparam Pixel_1_RNO_76_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_76_LC_5_11_4.LUT_INIT=16'b1000000111000010;
    LogicCell40 Pixel_1_RNO_76_LC_5_11_4 (
            .in0(N__9432),
            .in1(N__8526),
            .in2(N__7264),
            .in3(N__9253),
            .lcout(N_314_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15___m1_e_0_1_LC_5_11_5.C_ON=1'b0;
    defparam un115_pixel_13_15___m1_e_0_1_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15___m1_e_0_1_LC_5_11_5.LUT_INIT=16'b0000000010100000;
    LogicCell40 un115_pixel_13_15___m1_e_0_1_LC_5_11_5 (
            .in0(N__8936),
            .in1(_gnd_net_),
            .in2(N__9286),
            .in3(N__9429),
            .lcout(un115_pixel_13_15___m1_e_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__m9_0_LC_5_11_6.C_ON=1'b0;
    defparam un115_pixel_13_15__m9_0_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__m9_0_LC_5_11_6.LUT_INIT=16'b0100000010001000;
    LogicCell40 un115_pixel_13_15__m9_0_LC_5_11_6 (
            .in0(N__9430),
            .in1(N__8937),
            .in2(N__8774),
            .in3(N__9251),
            .lcout(un115_pixel_13_15__i2_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__g0_9_LC_5_11_7.C_ON=1'b0;
    defparam un115_pixel_13_15__g0_9_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__g0_9_LC_5_11_7.LUT_INIT=16'b0001001000000000;
    LogicCell40 un115_pixel_13_15__g0_9_LC_5_11_7 (
            .in0(N__9254),
            .in1(N__8726),
            .in2(N__9018),
            .in3(N__9433),
            .lcout(N_219_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_5_12_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_5_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__14085),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_2_s_LC_5_12_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_2_s_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_2_s_LC_5_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_cry_2_s_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(N__8262),
            .in2(N__11353),
            .in3(N__7318),
            .lcout(if_generate_plus_mult1_un75_sum_cry_2_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_12_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__8868),
            .in2(N__8305),
            .in3(N__7306),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_axb_5_LC_5_12_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_axb_5_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un82_sum_axb_5_LC_5_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un82_sum_axb_5_LC_5_12_3 (
            .in0(N__9181),
            .in1(N__8263),
            .in2(N__8293),
            .in3(N__7297),
            .lcout(un4_pixel_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_s_5_LC_5_12_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_s_5_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_s_5_LC_5_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_s_5_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(N__8278),
            .in2(_gnd_net_),
            .in3(N__7294),
            .lcout(un7_pixel_1_axb1),
            .ltout(un7_pixel_1_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__un115_pixel_1_i_9_LC_5_12_5.C_ON=1'b0;
    defparam un115_pixel_13_15__un115_pixel_1_i_9_LC_5_12_5.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__un115_pixel_1_i_9_LC_5_12_5.LUT_INIT=16'b1110001001001100;
    LogicCell40 un115_pixel_13_15__un115_pixel_1_i_9_LC_5_12_5 (
            .in0(N__8872),
            .in1(N__8735),
            .in2(N__7291),
            .in3(N__9426),
            .lcout(),
            .ltout(N_203_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_47_LC_5_12_6.C_ON=1'b0;
    defparam Pixel_1_RNO_47_LC_5_12_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_47_LC_5_12_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 Pixel_1_RNO_47_LC_5_12_6 (
            .in0(N__8571),
            .in1(_gnd_net_),
            .in2(N__7288),
            .in3(N__7285),
            .lcout(Pixel_1_RNOZ0Z_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_92_LC_5_12_7.C_ON=1'b0;
    defparam Pixel_1_RNO_92_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_92_LC_5_12_7.LUT_INIT=16'b0100010110001101;
    LogicCell40 Pixel_1_RNO_92_LC_5_12_7 (
            .in0(N__9182),
            .in1(N__8734),
            .in2(N__8951),
            .in3(N__9425),
            .lcout(g0_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__g0_7_LC_5_13_0.C_ON=1'b0;
    defparam un115_pixel_13_15__g0_7_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__g0_7_LC_5_13_0.LUT_INIT=16'b0000100000100000;
    LogicCell40 un115_pixel_13_15__g0_7_LC_5_13_0 (
            .in0(N__9406),
            .in1(N__8990),
            .in2(N__9264),
            .in3(N__8688),
            .lcout(N_192_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_72_LC_5_13_1.C_ON=1'b0;
    defparam Pixel_1_RNO_72_LC_5_13_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_72_LC_5_13_1.LUT_INIT=16'b1010010101111111;
    LogicCell40 Pixel_1_RNO_72_LC_5_13_1 (
            .in0(N__8689),
            .in1(N__9197),
            .in2(N__9040),
            .in3(N__9408),
            .lcout(Pixel_1_RNOZ0Z_72),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un115_pixel_13_15__g0_2_LC_5_13_2.C_ON=1'b0;
    defparam un115_pixel_13_15__g0_2_LC_5_13_2.SEQ_MODE=4'b0000;
    defparam un115_pixel_13_15__g0_2_LC_5_13_2.LUT_INIT=16'b0100100000101000;
    LogicCell40 un115_pixel_13_15__g0_2_LC_5_13_2 (
            .in0(N__9409),
            .in1(N__8995),
            .in2(N__9265),
            .in3(N__8691),
            .lcout(N_234_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_90_LC_5_13_3.C_ON=1'b0;
    defparam Pixel_1_RNO_90_LC_5_13_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_90_LC_5_13_3.LUT_INIT=16'b0000011110100001;
    LogicCell40 Pixel_1_RNO_90_LC_5_13_3 (
            .in0(N__8991),
            .in1(N__10146),
            .in2(N__9267),
            .in3(N__9407),
            .lcout(g0_40_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_65_LC_5_13_4.C_ON=1'b0;
    defparam Pixel_1_RNO_65_LC_5_13_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_65_LC_5_13_4.LUT_INIT=16'b1001010110001000;
    LogicCell40 Pixel_1_RNO_65_LC_5_13_4 (
            .in0(N__9410),
            .in1(N__8996),
            .in2(N__9266),
            .in3(N__8692),
            .lcout(N_206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_84_LC_5_13_5.C_ON=1'b0;
    defparam Pixel_1_RNO_84_LC_5_13_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_84_LC_5_13_5.LUT_INIT=16'b0101000101101111;
    LogicCell40 Pixel_1_RNO_84_LC_5_13_5 (
            .in0(N__8690),
            .in1(N__10147),
            .in2(N__9268),
            .in3(N__9411),
            .lcout(),
            .ltout(g0_6_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_57_LC_5_13_6.C_ON=1'b0;
    defparam Pixel_1_RNO_57_LC_5_13_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_57_LC_5_13_6.LUT_INIT=16'b1101101001111111;
    LogicCell40 Pixel_1_RNO_57_LC_5_13_6 (
            .in0(N__9204),
            .in1(N__10128),
            .in2(N__7360),
            .in3(N__8997),
            .lcout(),
            .ltout(g0_6_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_37_LC_5_13_7.C_ON=1'b0;
    defparam Pixel_1_RNO_37_LC_5_13_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_37_LC_5_13_7.LUT_INIT=16'b0011111100101110;
    LogicCell40 Pixel_1_RNO_37_LC_5_13_7 (
            .in0(N__10129),
            .in1(N__8568),
            .in2(N__7357),
            .in3(N__7354),
            .lcout(N_302_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_71_LC_5_14_0.C_ON=1'b0;
    defparam Pixel_1_RNO_71_LC_5_14_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_71_LC_5_14_0.LUT_INIT=16'b0101010001110000;
    LogicCell40 Pixel_1_RNO_71_LC_5_14_0 (
            .in0(N__8760),
            .in1(N__9260),
            .in2(N__9051),
            .in3(N__9422),
            .lcout(),
            .ltout(g1_3_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_46_LC_5_14_1.C_ON=1'b0;
    defparam Pixel_1_RNO_46_LC_5_14_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_46_LC_5_14_1.LUT_INIT=16'b0111101011011111;
    LogicCell40 Pixel_1_RNO_46_LC_5_14_1 (
            .in0(N__9423),
            .in1(N__8569),
            .in2(N__7342),
            .in3(N__9010),
            .lcout(g1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_85_LC_5_14_4.C_ON=1'b0;
    defparam Pixel_1_RNO_85_LC_5_14_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_85_LC_5_14_4.LUT_INIT=16'b0100010011101110;
    LogicCell40 Pixel_1_RNO_85_LC_5_14_4 (
            .in0(N__9011),
            .in1(N__10153),
            .in2(_gnd_net_),
            .in3(N__9424),
            .lcout(),
            .ltout(g0_10_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_58_LC_5_14_5.C_ON=1'b0;
    defparam Pixel_1_RNO_58_LC_5_14_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_58_LC_5_14_5.LUT_INIT=16'b0001011100110011;
    LogicCell40 Pixel_1_RNO_58_LC_5_14_5 (
            .in0(N__9261),
            .in1(N__10133),
            .in2(N__7327),
            .in3(N__8761),
            .lcout(),
            .ltout(N_309_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_38_LC_5_14_6.C_ON=1'b0;
    defparam Pixel_1_RNO_38_LC_5_14_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_38_LC_5_14_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 Pixel_1_RNO_38_LC_5_14_6 (
            .in0(N__8570),
            .in1(_gnd_net_),
            .in2(N__7420),
            .in3(N__7417),
            .lcout(),
            .ltout(N_323_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_21_LC_5_14_7.C_ON=1'b0;
    defparam Pixel_1_RNO_21_LC_5_14_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_21_LC_5_14_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 Pixel_1_RNO_21_LC_5_14_7 (
            .in0(_gnd_net_),
            .in1(N__11091),
            .in2(N__7411),
            .in3(N__7408),
            .lcout(N_5_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_6_2_7.C_ON=1'b0;
    defparam beamY_2_LC_6_2_7.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_6_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_2_LC_6_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8022),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13225),
            .ce(N__13275),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_6_3_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_6_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(N__10160),
            .in2(N__11128),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_RNIAL73_LC_6_3_1.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_6_3_1.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_6_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_1_c_RNIAL73_LC_6_3_1 (
            .in0(_gnd_net_),
            .in1(N__7466),
            .in2(_gnd_net_),
            .in3(N__7390),
            .lcout(un21_beamy_cry_1_c_RNIALZ0Z73),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_2_c_RNICO83_LC_6_3_2.C_ON=1'b1;
    defparam un21_beamy_cry_2_c_RNICO83_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_2_c_RNICO83_LC_6_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_2_c_RNICO83_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(N__7566),
            .in2(_gnd_net_),
            .in3(N__7387),
            .lcout(un21_beamy_cry_2_c_RNICOZ0Z83),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_3_c_RNIER93_LC_6_3_3.C_ON=1'b1;
    defparam un21_beamy_cry_3_c_RNIER93_LC_6_3_3.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_3_c_RNIER93_LC_6_3_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_3_c_RNIER93_LC_6_3_3 (
            .in0(_gnd_net_),
            .in1(N__7890),
            .in2(_gnd_net_),
            .in3(N__7384),
            .lcout(un21_beamy_cry_3_c_RNIERZ0Z93),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_6_3_4.C_ON=1'b1;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_6_3_4.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_6_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_4_c_RNIGUA3_LC_6_3_4 (
            .in0(_gnd_net_),
            .in1(N__10465),
            .in2(_gnd_net_),
            .in3(N__7381),
            .lcout(un21_beamy_cry_4_c_RNIGUAZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_5_c_RNII1C3_LC_6_3_5.C_ON=1'b1;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_6_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_5_c_RNII1C3_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(N__10558),
            .in2(_gnd_net_),
            .in3(N__7378),
            .lcout(un21_beamy_cry_5_c_RNII1CZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_6_3_6.C_ON=1'b1;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_6_3_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_6_c_RNIK4D3_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(N__11004),
            .in2(_gnd_net_),
            .in3(N__7624),
            .lcout(un21_beamy_cry_6_c_RNIK4DZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_6_3_7.C_ON=1'b1;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_6_3_7.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_6_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_7_c_RNIM7E3_LC_6_3_7 (
            .in0(_gnd_net_),
            .in1(N__10793),
            .in2(_gnd_net_),
            .in3(N__7612),
            .lcout(un21_beamy_cry_7_c_RNIM7EZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_6_4_0.C_ON=1'b0;
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_6_4_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 un21_beamy_cry_8_c_RNIOAF3_LC_6_4_0 (
            .in0(N__10880),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7609),
            .lcout(un21_beamy_cry_8_c_RNIOAFZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5NLM2_3_LC_6_4_1.C_ON=1'b0;
    defparam beamY_RNI5NLM2_3_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI5NLM2_3_LC_6_4_1.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNI5NLM2_3_LC_6_4_1 (
            .in0(N__11915),
            .in1(N__11810),
            .in2(N__7429),
            .in3(N__12146),
            .lcout(un11_visibleylto9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_4_2.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_4_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_4_2 (
            .in0(N__12080),
            .in1(N__14592),
            .in2(_gnd_net_),
            .in3(N__7482),
            .lcout(beamY_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_4_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_4_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_4_3 (
            .in0(N__9660),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIALEQ_0_9_LC_6_4_4.C_ON=1'b0;
    defparam beamY_RNIALEQ_0_9_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIALEQ_0_9_LC_6_4_4.LUT_INIT=16'b0101010101100110;
    LogicCell40 beamY_RNIALEQ_0_9_LC_6_4_4 (
            .in0(N__10879),
            .in1(N__7996),
            .in2(_gnd_net_),
            .in3(N__7974),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_s_4_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_0_3_LC_6_4_5.C_ON=1'b0;
    defparam beamY_RNI6125_0_3_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_0_3_LC_6_4_5.LUT_INIT=16'b0100000000100010;
    LogicCell40 beamY_RNI6125_0_3_LC_6_4_5 (
            .in0(N__10464),
            .in1(N__7585),
            .in2(N__7497),
            .in3(N__7879),
            .lcout(un11_visibleylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_6_4_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_6_4_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_6_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_6_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9595),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIEP79_7_LC_6_4_7.C_ON=1'b0;
    defparam beamY_fast_RNIEP79_7_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIEP79_7_LC_6_4_7.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_fast_RNIEP79_7_LC_6_4_7 (
            .in0(N__10463),
            .in1(N__7711),
            .in2(_gnd_net_),
            .in3(N__7694),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un40_sum_axbxc5_m3_a1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_6_LC_6_5_1.C_ON=1'b0;
    defparam beamY_fast_6_LC_6_5_1.SEQ_MODE=4'b1000;
    defparam beamY_fast_6_LC_6_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_6_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7917),
            .lcout(beamY_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13219),
            .ce(N__13273),
            .sr(_gnd_net_));
    defparam beamY_fast_7_LC_6_5_2.C_ON=1'b0;
    defparam beamY_fast_7_LC_6_5_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_7_LC_6_5_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_fast_7_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(N__7953),
            .in2(_gnd_net_),
            .in3(N__7816),
            .lcout(beamY_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13219),
            .ce(N__13273),
            .sr(_gnd_net_));
    defparam beamY_fast_5_LC_6_5_3.C_ON=1'b0;
    defparam beamY_fast_5_LC_6_5_3.SEQ_MODE=4'b1000;
    defparam beamY_fast_5_LC_6_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_5_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7731),
            .lcout(beamY_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13219),
            .ce(N__13273),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIRPUB_7_LC_6_5_4.C_ON=1'b0;
    defparam beamY_fast_RNIRPUB_7_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIRPUB_7_LC_6_5_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamY_fast_RNIRPUB_7_LC_6_5_4 (
            .in0(N__7710),
            .in1(N__7690),
            .in2(_gnd_net_),
            .in3(N__7661),
            .lcout(un5_visibley_c6_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFC4H3_9_LC_6_6_1.C_ON=1'b0;
    defparam beamY_RNIFC4H3_9_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIFC4H3_9_LC_6_6_1.LUT_INIT=16'b0100010010001000;
    LogicCell40 beamY_RNIFC4H3_9_LC_6_6_1 (
            .in0(N__10915),
            .in1(N__7645),
            .in2(_gnd_net_),
            .in3(N__10366),
            .lcout(un11_visibley),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI198K_2_LC_6_6_2.C_ON=1'b0;
    defparam beamY_fast_RNI198K_2_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI198K_2_LC_6_6_2.LUT_INIT=16'b1001001100110011;
    LogicCell40 beamY_fast_RNI198K_2_LC_6_6_2 (
            .in0(N__10712),
            .in1(N__10811),
            .in2(N__10597),
            .in3(N__10613),
            .lcout(),
            .ltout(beamY_fast_RNI198KZ0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQNF11_8_LC_6_6_3.C_ON=1'b0;
    defparam beamY_RNIQNF11_8_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIQNF11_8_LC_6_6_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 beamY_RNIQNF11_8_LC_6_6_3 (
            .in0(N__10812),
            .in1(_gnd_net_),
            .in2(N__7636),
            .in3(N__7973),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_54_LC_6_6_4.C_ON=1'b0;
    defparam Pixel_1_RNO_54_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_54_LC_6_6_4.LUT_INIT=16'b0000000000001000;
    LogicCell40 Pixel_1_RNO_54_LC_6_6_4 (
            .in0(N__10641),
            .in1(N__12691),
            .in2(N__11182),
            .in3(N__14422),
            .lcout(font_un127_pixel_m_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_2_LC_6_6_5.C_ON=1'b0;
    defparam beamY_fast_2_LC_6_6_5.SEQ_MODE=4'b1000;
    defparam beamY_fast_2_LC_6_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_2_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8026),
            .lcout(beamY_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13217),
            .ce(N__13271),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIG57D_8_LC_6_6_6.C_ON=1'b0;
    defparam beamY_fast_RNIG57D_8_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIG57D_8_LC_6_6_6.LUT_INIT=16'b1111100011110000;
    LogicCell40 beamY_fast_RNIG57D_8_LC_6_6_6 (
            .in0(N__10711),
            .in1(N__10612),
            .in2(N__8011),
            .in3(N__7853),
            .lcout(beamY_fast_RNIG57DZ0Z_8),
            .ltout(beamY_fast_RNIG57DZ0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIBV5P_8_LC_6_6_7.C_ON=1'b0;
    defparam beamY_fast_RNIBV5P_8_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIBV5P_8_LC_6_6_7.LUT_INIT=16'b1111111111110000;
    LogicCell40 beamY_fast_RNIBV5P_8_LC_6_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7981),
            .in3(N__7972),
            .lcout(un5_visibley_c7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_7_LC_6_7_0.C_ON=1'b0;
    defparam beamY_7_LC_6_7_0.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_6_7_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_7_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(N__7954),
            .in2(_gnd_net_),
            .in3(N__7786),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam beamY_fast_3_LC_6_7_1.C_ON=1'b0;
    defparam beamY_fast_3_LC_6_7_1.SEQ_MODE=4'b1000;
    defparam beamY_fast_3_LC_6_7_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_fast_3_LC_6_7_1 (
            .in0(N__7787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7936),
            .lcout(beamY_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam beamY_6_LC_6_7_3.C_ON=1'b0;
    defparam beamY_6_LC_6_7_3.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_6_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_6_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7918),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam beamY_4_LC_6_7_4.C_ON=1'b0;
    defparam beamY_4_LC_6_7_4.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_6_7_4.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_4_LC_6_7_4 (
            .in0(N__7755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7784),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam beamY_4_rep1_LC_6_7_5.C_ON=1'b0;
    defparam beamY_4_rep1_LC_6_7_5.SEQ_MODE=4'b1000;
    defparam beamY_4_rep1_LC_6_7_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_4_rep1_LC_6_7_5 (
            .in0(N__7785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7756),
            .lcout(beamY_4_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam beamY_5_LC_6_7_6.C_ON=1'b0;
    defparam beamY_5_LC_6_7_6.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_6_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_5_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7735),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13216),
            .ce(N__13270),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_1_LC_6_8_0.C_ON=1'b0;
    defparam Pixel_1_RNO_1_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_1_LC_6_8_0.LUT_INIT=16'b1110010000000000;
    LogicCell40 Pixel_1_RNO_1_LC_6_8_0 (
            .in0(N__13179),
            .in1(N__11377),
            .in2(N__8128),
            .in3(N__8056),
            .lcout(),
            .ltout(font_un127_pixel_m_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_6_8_1.C_ON=1'b0;
    defparam Pixel_1_LC_6_8_1.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_6_8_1.LUT_INIT=16'b1110111011110000;
    LogicCell40 Pixel_1_LC_6_8_1 (
            .in0(N__8090),
            .in1(N__12787),
            .in2(N__8119),
            .in3(N__10621),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13213),
            .ce(),
            .sr(N__11337));
    defparam Pixel_1_RNO_16_LC_6_8_2.C_ON=1'b0;
    defparam Pixel_1_RNO_16_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_16_LC_6_8_2.LUT_INIT=16'b0100010100000000;
    LogicCell40 Pixel_1_RNO_16_LC_6_8_2 (
            .in0(N__8224),
            .in1(N__12690),
            .in2(N__14421),
            .in3(N__8077),
            .lcout(),
            .ltout(g0_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_5_LC_6_8_3.C_ON=1'b0;
    defparam Pixel_1_RNO_5_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_5_LC_6_8_3.LUT_INIT=16'b0001000011100000;
    LogicCell40 Pixel_1_RNO_5_LC_6_8_3 (
            .in0(N__8563),
            .in1(N__10144),
            .in2(N__8071),
            .in3(N__8068),
            .lcout(g0_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_9_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__13066),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JF_LC_6_9_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JF_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JF_LC_6_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JF_LC_6_9_1 (
            .in0(_gnd_net_),
            .in1(N__8215),
            .in2(N__8043),
            .in3(N__8050),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNIT3JFZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_82_LC_6_9_2.C_ON=1'b1;
    defparam Pixel_1_RNO_82_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_82_LC_6_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_82_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__10750),
            .in2(N__11200),
            .in3(N__8047),
            .lcout(Pixel_1_RNOZ0Z_82),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_6_9_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_6_9_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_6_9_3 (
            .in0(_gnd_net_),
            .in1(N__11248),
            .in2(N__8044),
            .in3(N__11195),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJ2_LC_6_9_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJ2_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJ2_LC_6_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJ2_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__11218),
            .in2(_gnd_net_),
            .in3(N__8029),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2),
            .ltout(font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI022VJZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_31_LC_6_9_5.C_ON=1'b0;
    defparam Pixel_1_RNO_31_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_31_LC_6_9_5.LUT_INIT=16'b0101000001010000;
    LogicCell40 Pixel_1_RNO_31_LC_6_9_5 (
            .in0(N__13069),
            .in1(_gnd_net_),
            .in2(N__8245),
            .in3(_gnd_net_),
            .lcout(g1_0_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_83_LC_6_9_6.C_ON=1'b0;
    defparam Pixel_1_RNO_83_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_83_LC_6_9_6.LUT_INIT=16'b0101010101100110;
    LogicCell40 Pixel_1_RNO_83_LC_6_9_6 (
            .in0(N__13180),
            .in1(N__13067),
            .in2(_gnd_net_),
            .in3(N__11433),
            .lcout(),
            .ltout(font_un127_pixel_m_4_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_55_LC_6_9_7.C_ON=1'b0;
    defparam Pixel_1_RNO_55_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_55_LC_6_9_7.LUT_INIT=16'b0100000110000010;
    LogicCell40 Pixel_1_RNO_55_LC_6_9_7 (
            .in0(N__13068),
            .in1(N__8242),
            .in2(N__8236),
            .in3(N__8197),
            .lcout(font_un127_pixel_m_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_56_LC_6_10_0.C_ON=1'b0;
    defparam Pixel_1_RNO_56_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_56_LC_6_10_0.LUT_INIT=16'b0111011111111111;
    LogicCell40 Pixel_1_RNO_56_LC_6_10_0 (
            .in0(N__8950),
            .in1(N__9287),
            .in2(_gnd_net_),
            .in3(N__9492),
            .lcout(),
            .ltout(un7_pixel_1_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_36_LC_6_10_1.C_ON=1'b0;
    defparam Pixel_1_RNO_36_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_36_LC_6_10_1.LUT_INIT=16'b0101110111110111;
    LogicCell40 Pixel_1_RNO_36_LC_6_10_1 (
            .in0(N__11599),
            .in1(N__8796),
            .in2(N__8227),
            .in3(N__11524),
            .lcout(font_un127_pixel_m_7_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_6_10_2.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_6_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14086),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHMV0K2_LC_6_10_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHMV0K2_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHMV0K2_LC_6_10_4.LUT_INIT=16'b1100110000110011;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHMV0K2_LC_6_10_4 (
            .in0(_gnd_net_),
            .in1(N__13073),
            .in2(_gnd_net_),
            .in3(N__8198),
            .lcout(font_un13_pixel_0_1_0_0_22),
            .ltout(font_un13_pixel_0_1_0_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_32_LC_6_10_5.C_ON=1'b0;
    defparam Pixel_1_RNO_32_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_32_LC_6_10_5.LUT_INIT=16'b1111000111111011;
    LogicCell40 Pixel_1_RNO_32_LC_6_10_5 (
            .in0(N__11123),
            .in1(N__8167),
            .in2(N__8155),
            .in3(N__8374),
            .lcout(g1_4_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_29_LC_6_10_6.C_ON=1'b0;
    defparam Pixel_1_RNO_29_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_29_LC_6_10_6.LUT_INIT=16'b0010000001111111;
    LogicCell40 Pixel_1_RNO_29_LC_6_10_6 (
            .in0(N__10096),
            .in1(N__8152),
            .in2(N__11129),
            .in3(N__8137),
            .lcout(),
            .ltout(N_1482_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_13_LC_6_10_7.C_ON=1'b0;
    defparam Pixel_1_RNO_13_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_13_LC_6_10_7.LUT_INIT=16'b0000110000111111;
    LogicCell40 Pixel_1_RNO_13_LC_6_10_7 (
            .in0(_gnd_net_),
            .in1(N__11119),
            .in2(N__8308),
            .in3(N__8416),
            .lcout(N_1870_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(N__13970),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__8331),
            .in2(N__11284),
            .in3(N__8296),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(N__9427),
            .in2(N__8323),
            .in3(N__8281),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3 (
            .in0(N__8867),
            .in1(N__8332),
            .in2(N__9526),
            .in3(N__8272),
            .lcout(un4_pixel_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(N__9511),
            .in2(_gnd_net_),
            .in3(N__8269),
            .lcout(un7_pixel_1_axb2),
            .ltout(un7_pixel_1_axb2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_pixel_1_axb2_sbtinv_LC_6_11_5.C_ON=1'b0;
    defparam un7_pixel_1_axb2_sbtinv_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam un7_pixel_1_axb2_sbtinv_LC_6_11_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un7_pixel_1_axb2_sbtinv_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8266),
            .in3(_gnd_net_),
            .lcout(un7_pixel_1_axb2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_27_LC_6_11_6.C_ON=1'b0;
    defparam Pixel_1_RNO_27_LC_6_11_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_27_LC_6_11_6.LUT_INIT=16'b1100111011000100;
    LogicCell40 Pixel_1_RNO_27_LC_6_11_6 (
            .in0(N__8574),
            .in1(N__8254),
            .in2(N__10161),
            .in3(N__8362),
            .lcout(),
            .ltout(N_305_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_12_LC_6_11_7.C_ON=1'b0;
    defparam Pixel_1_RNO_12_LC_6_11_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_12_LC_6_11_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 Pixel_1_RNO_12_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(N__11124),
            .in2(N__8248),
            .in3(N__8395),
            .lcout(N_1869_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_77_LC_6_12_0.C_ON=1'b0;
    defparam Pixel_1_RNO_77_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_77_LC_6_12_0.LUT_INIT=16'b0110011111111110;
    LogicCell40 Pixel_1_RNO_77_LC_6_12_0 (
            .in0(N__9016),
            .in1(N__8389),
            .in2(N__8578),
            .in3(N__8790),
            .lcout(),
            .ltout(N_321_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_50_LC_6_12_1.C_ON=1'b0;
    defparam Pixel_1_RNO_50_LC_6_12_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_50_LC_6_12_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 Pixel_1_RNO_50_LC_6_12_1 (
            .in0(N__10151),
            .in1(_gnd_net_),
            .in2(N__8383),
            .in3(N__8380),
            .lcout(N_328_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_93_LC_6_12_2.C_ON=1'b0;
    defparam Pixel_1_RNO_93_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_93_LC_6_12_2.LUT_INIT=16'b1011111111111111;
    LogicCell40 Pixel_1_RNO_93_LC_6_12_2 (
            .in0(N__9367),
            .in1(N__9255),
            .in2(N__9052),
            .in3(N__8789),
            .lcout(),
            .ltout(g1_2_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_80_LC_6_12_3.C_ON=1'b0;
    defparam Pixel_1_RNO_80_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_80_LC_6_12_3.LUT_INIT=16'b0101000011111010;
    LogicCell40 Pixel_1_RNO_80_LC_6_12_3 (
            .in0(N__10150),
            .in1(_gnd_net_),
            .in2(N__8365),
            .in3(N__8358),
            .lcout(),
            .ltout(un117_pixel_6_1_0_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_52_LC_6_12_4.C_ON=1'b0;
    defparam Pixel_1_RNO_52_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_52_LC_6_12_4.LUT_INIT=16'b0001110000111110;
    LogicCell40 Pixel_1_RNO_52_LC_6_12_4 (
            .in0(N__8567),
            .in1(N__10152),
            .in2(N__8341),
            .in3(N__8338),
            .lcout(N_324_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_pixel_1_axb3_sbtinv_LC_6_12_5.C_ON=1'b0;
    defparam un7_pixel_1_axb3_sbtinv_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam un7_pixel_1_axb3_sbtinv_LC_6_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_pixel_1_axb3_sbtinv_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9366),
            .lcout(un7_pixel_1_axb3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_6_13_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_6_13_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_6_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(N__13868),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_2_s_LC_6_13_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_2_s_LC_6_13_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_2_s_LC_6_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_cry_2_s_LC_6_13_1 (
            .in0(_gnd_net_),
            .in1(N__8403),
            .in2(N__9073),
            .in3(N__8311),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_13_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_13_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(N__11517),
            .in2(N__11611),
            .in3(N__9514),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_axb_5_LC_6_13_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_axb_5_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_axb_5_LC_6_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_axb_5_LC_6_13_3 (
            .in0(N__9368),
            .in1(N__8404),
            .in2(N__11569),
            .in3(N__9502),
            .lcout(un4_pixel_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_s_5_LC_6_13_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_s_5_LC_6_13_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_s_5_LC_6_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_s_5_LC_6_13_4 (
            .in0(_gnd_net_),
            .in1(N__11542),
            .in2(_gnd_net_),
            .in3(N__9499),
            .lcout(un7_pixel_1_axb3),
            .ltout(un7_pixel_1_axb3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_89_LC_6_13_5.C_ON=1'b0;
    defparam Pixel_1_RNO_89_LC_6_13_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_89_LC_6_13_5.LUT_INIT=16'b0011101111000000;
    LogicCell40 Pixel_1_RNO_89_LC_6_13_5 (
            .in0(N__10145),
            .in1(N__8989),
            .in2(N__9292),
            .in3(N__9183),
            .lcout(un117_pixel_2_6_i3_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_N_532_i_LC_6_13_6.C_ON=1'b0;
    defparam un4_pixel_N_532_i_LC_6_13_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_N_532_i_LC_6_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_pixel_N_532_i_LC_6_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13763),
            .lcout(N_532_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_73_LC_6_14_0.C_ON=1'b0;
    defparam Pixel_1_RNO_73_LC_6_14_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_73_LC_6_14_0.LUT_INIT=16'b1000001010010011;
    LogicCell40 Pixel_1_RNO_73_LC_6_14_0 (
            .in0(N__9064),
            .in1(N__9012),
            .in2(N__8797),
            .in3(N__10148),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_73_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_48_LC_6_14_1.C_ON=1'b0;
    defparam Pixel_1_RNO_48_LC_6_14_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_48_LC_6_14_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 Pixel_1_RNO_48_LC_6_14_1 (
            .in0(_gnd_net_),
            .in1(N__8572),
            .in2(N__8587),
            .in3(N__8584),
            .lcout(),
            .ltout(Pixel_1_RNOZ0Z_48_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_30_LC_6_14_2.C_ON=1'b0;
    defparam Pixel_1_RNO_30_LC_6_14_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_30_LC_6_14_2.LUT_INIT=16'b1111000111100000;
    LogicCell40 Pixel_1_RNO_30_LC_6_14_2 (
            .in0(N__8573),
            .in1(N__10149),
            .in2(N__8425),
            .in3(N__8422),
            .lcout(d_N_3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_pixel_0_axb3_sbtinv_LC_6_14_5.C_ON=1'b0;
    defparam un7_pixel_0_axb3_sbtinv_LC_6_14_5.SEQ_MODE=4'b0000;
    defparam un7_pixel_0_axb3_sbtinv_LC_6_14_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_pixel_0_axb3_sbtinv_LC_6_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11515),
            .lcout(un7_pixel_0_axb3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_1_0 (
            .in0(_gnd_net_),
            .in1(N__9740),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_1_1 (
            .in0(_gnd_net_),
            .in1(N__11687),
            .in2(N__9604),
            .in3(N__9622),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_1_2 (
            .in0(_gnd_net_),
            .in1(N__11737),
            .in2(N__11692),
            .in3(N__9619),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTA2_LC_7_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTA2_LC_7_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTA2_LC_7_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTA2_LC_7_1_3 (
            .in0(_gnd_net_),
            .in1(N__11691),
            .in2(N__11728),
            .in3(N__9616),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIMBTAZ0Z2),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI809T4_LC_7_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI809T4_LC_7_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI809T4_LC_7_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI809T4_LC_7_1_4 (
            .in0(N__9811),
            .in1(N__9757),
            .in2(N__11716),
            .in3(N__9613),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_LC_7_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_LC_7_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(N__11704),
            .in2(_gnd_net_),
            .in3(N__9610),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2),
            .ltout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KMEZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_0_LC_7_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_0_LC_7_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_0_LC_7_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6KME2_0_LC_7_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9607),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_1_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_1_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11812),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(N__9586),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQO93_LC_7_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQO93_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQO93_LC_7_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQO93_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(N__9812),
            .in2(N__9673),
            .in3(N__9829),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIHQOZ0Z93),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFP3_LC_7_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFP3_LC_7_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFP3_LC_7_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFP3_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(N__9826),
            .in2(N__9817),
            .in3(N__9820),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNI2HFPZ0Z3),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGC94_LC_7_2_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGC94_LC_7_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGC94_LC_7_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGC94_LC_7_2_3 (
            .in0(_gnd_net_),
            .in1(N__9816),
            .in2(N__9796),
            .in3(N__9787),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHGCZ0Z94),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV5NMA_LC_7_2_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV5NMA_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV5NMA_LC_7_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV5NMA_LC_7_2_4 (
            .in0(N__9882),
            .in1(N__9784),
            .in2(N__9778),
            .in3(N__9769),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_LC_7_2_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_LC_7_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_LC_7_2_5 (
            .in0(_gnd_net_),
            .in1(N__9766),
            .in2(_gnd_net_),
            .in3(N__9760),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6DZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_2_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11685),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_7_2_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_7_2_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_7_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_7_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9741),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_3_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__9652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLK5_LC_7_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLK5_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLK5_LC_7_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLK5_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__9877),
            .in2(N__9937),
            .in3(N__9928),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIMPLKZ0Z5),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAP8_LC_7_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAP8_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAP8_LC_7_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAP8_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__9925),
            .in2(N__9883),
            .in3(N__9919),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIPGAPZ0Z8),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIB9299_LC_7_3_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIB9299_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIB9299_LC_7_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIB9299_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(N__9881),
            .in2(N__9916),
            .in3(N__9907),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIBZ0Z9299),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIVO5IK_LC_7_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIVO5IK_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIVO5IK_LC_7_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIVO5IK_LC_7_3_4 (
            .in0(N__10247),
            .in1(N__9859),
            .in2(N__9904),
            .in3(N__9895),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PA_LC_7_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PA_LC_7_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PA_LC_7_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PA_LC_7_3_5 (
            .in0(_gnd_net_),
            .in1(N__9892),
            .in2(_gnd_net_),
            .in3(N__9886),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNI4E5PAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_0_LC_7_3_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_0_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_0_LC_7_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI6K6D5_0_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9876),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_4_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__12072),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5B_LC_7_4_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5B_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5B_LC_7_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5B_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__9853),
            .in2(N__10248),
            .in3(N__9844),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIP9V5BZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMG_LC_7_4_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMG_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMG_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMG_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__10243),
            .in2(N__9841),
            .in3(N__9832),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIQIDMGZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_18_LC_7_4_3.C_ON=1'b1;
    defparam Pixel_1_RNO_18_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_18_LC_7_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_18_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__10270),
            .in2(N__10249),
            .in3(N__10264),
            .lcout(Pixel_1_RNOZ0Z_18),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_4_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_4_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(N__10222),
            .in2(N__10261),
            .in3(N__10239),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQK_LC_7_4_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQK_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQK_LC_7_4_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQK_LC_7_4_5 (
            .in0(N__10216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10210),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2ARQKZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_6_LC_7_4_6.C_ON=1'b0;
    defparam Pixel_1_RNO_6_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_6_LC_7_4_6.LUT_INIT=16'b1010101010011010;
    LogicCell40 Pixel_1_RNO_6_LC_7_4_6 (
            .in0(N__10207),
            .in1(N__12037),
            .in2(N__10201),
            .in3(N__10183),
            .lcout(un1_beamY_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIALEQ_1_9_LC_7_4_7.C_ON=1'b0;
    defparam beamY_RNIALEQ_1_9_LC_7_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIALEQ_1_9_LC_7_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNIALEQ_1_9_LC_7_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10194),
            .lcout(beamY_RNIALEQ_1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_20_LC_7_5_0.C_ON=1'b0;
    defparam Pixel_1_RNO_20_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_20_LC_7_5_0.LUT_INIT=16'b0001100010001000;
    LogicCell40 Pixel_1_RNO_20_LC_7_5_0 (
            .in0(N__12049),
            .in1(N__10182),
            .in2(N__12084),
            .in3(N__10170),
            .lcout(),
            .ltout(un43lto4_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_9_LC_7_5_1.C_ON=1'b0;
    defparam Pixel_1_RNO_9_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_9_LC_7_5_1.LUT_INIT=16'b1000000001000000;
    LogicCell40 Pixel_1_RNO_9_LC_7_5_1 (
            .in0(N__10171),
            .in1(N__10162),
            .in2(N__9949),
            .in3(N__12079),
            .lcout(),
            .ltout(un43lt10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_2_LC_7_5_2.C_ON=1'b0;
    defparam Pixel_1_RNO_2_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_2_LC_7_5_2.LUT_INIT=16'b0001000100011110;
    LogicCell40 Pixel_1_RNO_2_LC_7_5_2 (
            .in0(N__10291),
            .in1(N__10372),
            .in2(N__9946),
            .in3(N__9943),
            .lcout(un44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_8_LC_7_5_4.C_ON=1'b0;
    defparam Pixel_1_RNO_8_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_8_LC_7_5_4.LUT_INIT=16'b1001100011000100;
    LogicCell40 Pixel_1_RNO_8_LC_7_5_4 (
            .in0(N__13882),
            .in1(N__10312),
            .in2(N__13990),
            .in3(N__10318),
            .lcout(un42lt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIALEQ_9_LC_7_5_5.C_ON=1'b0;
    defparam beamY_RNIALEQ_9_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIALEQ_9_LC_7_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIALEQ_9_LC_7_5_5 (
            .in0(_gnd_net_),
            .in1(N__10924),
            .in2(_gnd_net_),
            .in3(N__10361),
            .lcout(beamY_RNIALEQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_6_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(N__13880),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_7_6_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_7_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__10329),
            .in2(N__11368),
            .in3(N__10336),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_19_LC_7_6_2.C_ON=1'b1;
    defparam Pixel_1_RNO_19_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_19_LC_7_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_19_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(N__12031),
            .in2(N__11995),
            .in3(N__10333),
            .lcout(Pixel_1_RNOZ0Z_19),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_6_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_6_3 (
            .in0(_gnd_net_),
            .in1(N__10330),
            .in2(N__12019),
            .in3(N__11990),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5AS_LC_7_6_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5AS_LC_7_6_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5AS_LC_7_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5AS_LC_7_6_4 (
            .in0(_gnd_net_),
            .in1(N__12007),
            .in2(_gnd_net_),
            .in3(N__10321),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0),
            .ltout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIAF5ASZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_7_LC_7_6_5.C_ON=1'b0;
    defparam Pixel_1_RNO_7_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_7_LC_7_6_5.LUT_INIT=16'b0100111110110000;
    LogicCell40 Pixel_1_RNO_7_LC_7_6_5 (
            .in0(N__13881),
            .in1(N__10311),
            .in2(N__10300),
            .in3(N__10297),
            .lcout(un1_visiblex_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIHT1O_3_LC_7_6_6.C_ON=1'b0;
    defparam beamY_fast_RNIHT1O_3_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIHT1O_3_LC_7_6_6.LUT_INIT=16'b1111000001000100;
    LogicCell40 beamY_fast_RNIHT1O_3_LC_7_6_6 (
            .in0(N__10555),
            .in1(N__10451),
            .in2(N__10567),
            .in3(N__10714),
            .lcout(un5_visibley_ac0_7),
            .ltout(un5_visibley_ac0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4S2S1_7_LC_7_6_7.C_ON=1'b0;
    defparam beamY_RNI4S2S1_7_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI4S2S1_7_LC_7_6_7.LUT_INIT=16'b1010100101010110;
    LogicCell40 beamY_RNI4S2S1_7_LC_7_6_7 (
            .in0(N__10985),
            .in1(N__10556),
            .in2(N__10738),
            .in3(N__12133),
            .lcout(font_un36_pixel_if_generate_plus_mult1_un47_sum_axb4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_4_rep1_RNICDQE_LC_7_7_0.C_ON=1'b0;
    defparam beamY_4_rep1_RNICDQE_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam beamY_4_rep1_RNICDQE_LC_7_7_0.LUT_INIT=16'b1111000011100001;
    LogicCell40 beamY_4_rep1_RNICDQE_LC_7_7_0 (
            .in0(N__10439),
            .in1(N__10527),
            .in2(N__10991),
            .in3(N__10593),
            .lcout(),
            .ltout(beamY_4_rep1_RNICDQEZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIB5JQ_7_LC_7_7_1.C_ON=1'b0;
    defparam beamY_RNIB5JQ_7_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIB5JQ_7_LC_7_7_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 beamY_RNIB5JQ_7_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__10378),
            .in2(N__10717),
            .in3(N__10665),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIBVU7_2_LC_7_7_3.C_ON=1'b0;
    defparam beamY_fast_RNIBVU7_2_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIBVU7_2_LC_7_7_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_fast_RNIBVU7_2_LC_7_7_3 (
            .in0(_gnd_net_),
            .in1(N__10713),
            .in2(_gnd_net_),
            .in3(N__10614),
            .lcout(un5_visibley_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_0_LC_7_7_4.C_ON=1'b0;
    defparam Pixel_1_RNO_0_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_0_LC_7_7_4.LUT_INIT=16'b0001101100010001;
    LogicCell40 Pixel_1_RNO_0_LC_7_7_4 (
            .in0(N__12783),
            .in1(N__12762),
            .in2(N__10645),
            .in3(N__10630),
            .lcout(Pixel_1_e_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIK8HH_2_LC_7_7_6.C_ON=1'b0;
    defparam beamY_fast_RNIK8HH_2_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIK8HH_2_LC_7_7_6.LUT_INIT=16'b0011001000110000;
    LogicCell40 beamY_fast_RNIK8HH_2_LC_7_7_6 (
            .in0(N__10615),
            .in1(N__10528),
            .in2(N__10462),
            .in3(N__10594),
            .lcout(beamY_fast_RNIK8HHZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKOP3_7_LC_7_7_7.C_ON=1'b0;
    defparam beamY_RNIKOP3_7_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIKOP3_7_LC_7_7_7.LUT_INIT=16'b1100110010011001;
    LogicCell40 beamY_RNIKOP3_7_LC_7_7_7 (
            .in0(N__10526),
            .in1(N__10969),
            .in2(_gnd_net_),
            .in3(N__10435),
            .lcout(beamY_RNIKOP3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__13982),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKB_LC_7_8_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKB_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKB_LC_7_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKB_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__11014),
            .in2(N__12276),
            .in3(N__11029),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIHANKBZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONH_LC_7_8_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONH_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONH_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONH_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__12295),
            .in2(N__12334),
            .in3(N__11026),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIMUONHZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI0MA3B1_LC_7_8_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI0MA3B1_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI0MA3B1_LC_7_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI0MA3B1_LC_7_8_3 (
            .in0(N__11259),
            .in1(N__12322),
            .in2(N__12277),
            .in3(N__11023),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_LC_7_8_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_LC_7_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__12313),
            .in2(_gnd_net_),
            .in3(N__11020),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0),
            .ltout(font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77MZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_0_LC_7_8_5.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_0_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_0_LC_7_8_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A77M_0_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11017),
            .in3(_gnd_net_),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_8_6.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13870),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMJIF_8_LC_7_8_7.C_ON=1'b0;
    defparam beamY_RNIMJIF_8_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIMJIF_8_LC_7_8_7.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNIMJIF_8_LC_7_8_7 (
            .in0(N__10987),
            .in1(N__10925),
            .in2(N__10831),
            .in3(N__10819),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_9_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_9_0 (
            .in0(_gnd_net_),
            .in1(N__14090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGM_LC_7_9_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGM_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGM_LC_7_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGM_LC_7_9_1 (
            .in0(_gnd_net_),
            .in1(N__12403),
            .in2(N__11232),
            .in3(N__10741),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI18KGMZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPC321_LC_7_9_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPC321_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPC321_LC_7_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPC321_LC_7_9_2 (
            .in0(_gnd_net_),
            .in1(N__11269),
            .in2(N__11263),
            .in3(N__11242),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNIUPCZ0Z321),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJFAHJ2_LC_7_9_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJFAHJ2_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJFAHJ2_LC_7_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJFAHJ2_LC_7_9_3 (
            .in0(N__11199),
            .in1(N__11239),
            .in2(N__11233),
            .in3(N__11212),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQAB1_LC_7_9_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQAB1_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQAB1_LC_7_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQAB1_LC_7_9_4 (
            .in0(_gnd_net_),
            .in1(N__11209),
            .in2(_gnd_net_),
            .in3(N__11203),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIFVQABZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_81_LC_7_9_5.C_ON=1'b0;
    defparam Pixel_1_RNO_81_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_81_LC_7_9_5.LUT_INIT=16'b1010100000000000;
    LogicCell40 Pixel_1_RNO_81_LC_7_9_5 (
            .in0(N__13642),
            .in1(N__13869),
            .in2(N__11167),
            .in3(N__13765),
            .lcout(un14_visibleylt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_94_LC_7_9_6.C_ON=1'b0;
    defparam Pixel_1_RNO_94_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_94_LC_7_9_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 Pixel_1_RNO_94_LC_7_9_6 (
            .in0(N__13070),
            .in1(N__14091),
            .in2(_gnd_net_),
            .in3(N__13983),
            .lcout(un14_visibleylt4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_7_9_7.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_7_9_7.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamX_RNIQCL_1_LC_7_9_7 (
            .in0(N__14123),
            .in1(N__13120),
            .in2(N__14038),
            .in3(N__13178),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_10_LC_7_10_1.C_ON=1'b0;
    defparam beamX_RNICPU5_10_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_10_LC_7_10_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNICPU5_10_LC_7_10_1 (
            .in0(N__13927),
            .in1(N__14128),
            .in2(N__13390),
            .in3(N__13118),
            .lcout(),
            .ltout(un3_beamx_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_3_LC_7_10_2.C_ON=1'b0;
    defparam beamX_RNIKVE6_3_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_3_LC_7_10_2.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNIKVE6_3_LC_7_10_2 (
            .in0(N__13693),
            .in1(N__14037),
            .in2(N__11158),
            .in3(N__13168),
            .lcout(un3_beamx_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_33_LC_7_10_3.C_ON=1'b0;
    defparam Pixel_1_RNO_33_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_33_LC_7_10_3.LUT_INIT=16'b0000000001010011;
    LogicCell40 Pixel_1_RNO_33_LC_7_10_3 (
            .in0(N__11155),
            .in1(N__11143),
            .in2(N__11130),
            .in3(N__11385),
            .lcout(),
            .ltout(g3_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_14_LC_7_10_4.C_ON=1'b0;
    defparam Pixel_1_RNO_14_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_14_LC_7_10_4.LUT_INIT=16'b1111100101100000;
    LogicCell40 Pixel_1_RNO_14_LC_7_10_4 (
            .in0(N__11443),
            .in1(N__11436),
            .in2(N__11410),
            .in3(N__11407),
            .lcout(),
            .ltout(font_un127_pixel_6_ns_1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_4_LC_7_10_5.C_ON=1'b0;
    defparam Pixel_1_RNO_4_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_4_LC_7_10_5.LUT_INIT=16'b1010110000001111;
    LogicCell40 Pixel_1_RNO_4_LC_7_10_5 (
            .in0(N__11401),
            .in1(N__11395),
            .in2(N__11389),
            .in3(N__11386),
            .lcout(N_520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_10_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_7_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13762),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_i_LC_7_11_3.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_i_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un68_sum_i_LC_7_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un68_sum_i_LC_7_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13971),
            .lcout(un4_pixel_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_7_11_5.C_ON=1'b0;
    defparam VSync_1_LC_7_11_5.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_7_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 VSync_1_LC_7_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11338),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13222),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_i_LC_7_11_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_i_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_i_LC_7_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_i_LC_7_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13856),
            .lcout(un4_pixel_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_12_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(N__13641),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_2_LC_7_12_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_2_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_2_LC_7_12_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_m_2_LC_7_12_1 (
            .in0(N__11464),
            .in1(N__14406),
            .in2(N__12523),
            .in3(N__11272),
            .lcout(if_generate_plus_mult1_un47_sum_m_2),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_12_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_12_2 (
            .in0(_gnd_net_),
            .in1(N__12565),
            .in2(N__12544),
            .in3(N__11473),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum1_3),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_12_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_12_3 (
            .in0(_gnd_net_),
            .in1(N__14407),
            .in2(N__12574),
            .in3(N__11470),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum1_4),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_12_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_12_4.LUT_INIT=16'b1000000001111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_12_4 (
            .in0(N__14408),
            .in1(N__13521),
            .in2(N__14707),
            .in3(N__11467),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_13_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_13_0 (
            .in0(_gnd_net_),
            .in1(N__13634),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_13_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_13_1 (
            .in0(_gnd_net_),
            .in1(N__12550),
            .in2(N__12559),
            .in3(N__11458),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum0_2),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_13_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_13_2 (
            .in0(_gnd_net_),
            .in1(N__12724),
            .in2(N__12718),
            .in3(N__11455),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum0_3),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_13_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_13_3 (
            .in0(_gnd_net_),
            .in1(N__12709),
            .in2(N__12619),
            .in3(N__11452),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum0_4),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_13_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_13_4 (
            .in0(_gnd_net_),
            .in1(N__14409),
            .in2(_gnd_net_),
            .in3(N__11449),
            .lcout(un4_pixel_if_generate_plus_mult1_un47_sum0_5),
            .ltout(un4_pixel_if_generate_plus_mult1_un47_sum0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_5_LC_7_13_5.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_5_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_5_LC_7_13_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_m_5_LC_7_13_5 (
            .in0(N__11628),
            .in1(_gnd_net_),
            .in2(N__11446),
            .in3(N__14413),
            .lcout(un7_pixel_0_axb4),
            .ltout(un7_pixel_0_axb4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_axb_5_LC_7_13_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_axb_5_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_axb_5_LC_7_13_6.LUT_INIT=16'b1100001110100101;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un54_sum_axb_5_LC_7_13_6 (
            .in0(N__11644),
            .in1(N__11638),
            .in2(N__11632),
            .in3(N__14411),
            .lcout(un4_pixel_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_un7_pixel_0_axb4_i_LC_7_13_7.C_ON=1'b0;
    defparam un4_pixel_un7_pixel_0_axb4_i_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam un4_pixel_un7_pixel_0_axb4_i_LC_7_13_7.LUT_INIT=16'b0000010110101111;
    LogicCell40 un4_pixel_un7_pixel_0_axb4_i_LC_7_13_7 (
            .in0(N__14410),
            .in1(_gnd_net_),
            .in2(N__11629),
            .in3(N__11617),
            .lcout(un7_pixel_0_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0 (
            .in0(_gnd_net_),
            .in1(N__13760),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(un4_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_14_1.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_14_1 (
            .in0(_gnd_net_),
            .in1(N__12535),
            .in2(N__11556),
            .in3(N__11602),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(un4_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_2.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_14_2 (
            .in0(_gnd_net_),
            .in1(N__11592),
            .in2(N__11581),
            .in3(N__11560),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un4_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_axb_5_LC_7_14_3.C_ON=1'b1;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_axb_5_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un61_sum_axb_5_LC_7_14_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un61_sum_axb_5_LC_7_14_3 (
            .in0(N__11516),
            .in1(N__11479),
            .in2(N__11557),
            .in3(N__11536),
            .lcout(un4_pixel_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(un4_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un4_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_s_5_LC_7_14_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_s_5_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un54_sum_s_5_LC_7_14_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un54_sum_s_5_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(N__11533),
            .in2(_gnd_net_),
            .in3(N__11527),
            .lcout(un7_pixel_0_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_3_LC_7_14_7.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_3_LC_7_14_7.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_3_LC_7_14_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_m_3_LC_7_14_7 (
            .in0(N__11494),
            .in1(N__11485),
            .in2(_gnd_net_),
            .in3(N__14412),
            .lcout(if_generate_plus_mult1_un47_sum_m_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_2_0 (
            .in0(_gnd_net_),
            .in1(N__11811),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_2_1 (
            .in0(_gnd_net_),
            .in1(N__11947),
            .in2(N__11851),
            .in3(N__11731),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689H1_LC_8_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689H1_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689H1_LC_8_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689H1_LC_8_2_2 (
            .in0(_gnd_net_),
            .in1(N__11665),
            .in2(N__11953),
            .in3(N__11719),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNI689HZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_8_2_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_8_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_8_2_3 (
            .in0(_gnd_net_),
            .in1(N__11951),
            .in2(N__11656),
            .in3(N__11707),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI69052_LC_8_2_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI69052_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI69052_LC_8_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI69052_LC_8_2_4 (
            .in0(N__11686),
            .in1(N__11932),
            .in2(N__11977),
            .in3(N__11698),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_2_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_2_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_2_5 (
            .in0(N__11965),
            .in1(N__11952),
            .in2(N__12172),
            .in3(N__11695),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_3_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__11916),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHT921_LC_8_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHT921_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHT921_LC_8_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHT921_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(N__12091),
            .in2(N__14606),
            .in3(N__11659),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHTZ0Z921),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(N__11836),
            .in2(N__14556),
            .in3(N__11647),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_3_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_3_3 (
            .in0(_gnd_net_),
            .in1(N__11821),
            .in2(N__14607),
            .in3(N__11968),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_3_4 (
            .in0(_gnd_net_),
            .in1(N__12164),
            .in2(_gnd_net_),
            .in3(N__11959),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(N__12181),
            .in2(_gnd_net_),
            .in3(N__11956),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_8_3_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_8_3_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11935),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_3_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_3_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_3_7 (
            .in0(N__11917),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_4_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__12147),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_8_4_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_8_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__11842),
            .in2(N__14608),
            .in3(N__11830),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_8_4_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_8_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__11827),
            .in2(N__14609),
            .in3(N__11815),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_4_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12184),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_4_4.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_4_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12175),
            .in3(N__12168),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQNF11_0_8_LC_8_4_7.C_ON=1'b0;
    defparam beamY_RNIQNF11_0_8_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIQNF11_0_8_LC_8_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 beamY_RNIQNF11_0_8_LC_8_4_7 (
            .in0(N__12148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_RNIQNF11_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_17_LC_8_5_5.C_ON=1'b0;
    defparam Pixel_1_RNO_17_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_17_LC_8_5_5.LUT_INIT=16'b1111111100110011;
    LogicCell40 Pixel_1_RNO_17_LC_8_5_5 (
            .in0(_gnd_net_),
            .in1(N__12085),
            .in2(_gnd_net_),
            .in3(N__12048),
            .lcout(un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_8_6_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__13764),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VG6_LC_8_6_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VG6_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VG6_LC_8_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VG6_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__12247),
            .in2(N__12256),
            .in3(N__12022),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK3VGZ0Z6),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6N9_LC_8_6_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6N9_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6N9_LC_8_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6N9_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(N__12241),
            .in2(N__12205),
            .in3(N__12010),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIGU6NZ0Z9),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIE7K6S_LC_8_6_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIE7K6S_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIE7K6S_LC_8_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIE7K6S_LC_8_6_3 (
            .in0(N__11994),
            .in1(N__12262),
            .in2(N__12232),
            .in3(N__12001),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07C_LC_8_6_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07C_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07C_LC_8_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07C_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(N__12217),
            .in2(_gnd_net_),
            .in3(N__11998),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI7L07CZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPA_LC_8_6_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPA_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPA_LC_8_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPA_LC_8_6_5 (
            .in0(N__12231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12200),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI4UVPAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_8_6_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_8_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13637),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_0_LC_8_6_7.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_0_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_0_LC_8_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_0_LC_8_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12199),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_7_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(N__13636),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMS983_LC_8_7_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMS983_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMS983_LC_8_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMS983_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(N__12342),
            .in2(N__12472),
            .in3(N__12235),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMSZ0Z983),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAO4_LC_8_7_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAO4_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAO4_LC_8_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAO4_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__12607),
            .in2(N__12460),
            .in3(N__12220),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI6NAOZ0Z4),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI9MMPB_LC_8_7_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI9MMPB_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI9MMPB_LC_8_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI9MMPB_LC_8_7_3 (
            .in0(N__12204),
            .in1(N__12343),
            .in2(N__12442),
            .in3(N__12211),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_LC_8_7_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_LC_8_7_4.LUT_INIT=16'b0101010110101010;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6L16_LC_8_7_4 (
            .in0(N__12427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12208),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIU6LZ0Z16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI8P51_4_LC_8_7_5.C_ON=1'b0;
    defparam beamX_RNI8P51_4_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam beamX_RNI8P51_4_LC_8_7_5.LUT_INIT=16'b0011000100110011;
    LogicCell40 beamX_RNI8P51_4_LC_8_7_5 (
            .in0(N__13925),
            .in1(N__13686),
            .in2(N__12844),
            .in3(N__13808),
            .lcout(un13_beamylt7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_8_7_6.C_ON=1'b0;
    defparam HSync_1_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_8_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 HSync_1_LC_8_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12763),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13220),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_0_LC_8_7_7.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_0_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_0_LC_8_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_0_LC_8_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12606),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_8_8_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_8_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13879),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRF156_LC_8_8_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRF156_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRF156_LC_8_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRF156_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__12301),
            .in2(N__12903),
            .in3(N__12325),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNIRFZ0Z156),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RA99_LC_8_8_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RA99_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RA99_LC_8_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RA99_LC_8_8_2 (
            .in0(_gnd_net_),
            .in1(N__12919),
            .in2(N__12973),
            .in3(N__12316),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI4RAZ0Z99),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIOK72M_LC_8_8_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIOK72M_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIOK72M_LC_8_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIOK72M_LC_8_8_3 (
            .in0(N__12294),
            .in1(N__12952),
            .in2(N__12904),
            .in3(N__12307),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_LC_8_8_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_LC_8_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_LC_8_8_4 (
            .in0(_gnd_net_),
            .in1(N__12937),
            .in2(_gnd_net_),
            .in3(N__12304),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_8_8_5.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_8_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_8_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13761),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_0_LC_8_8_7.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_0_LC_8_8_7.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_0_LC_8_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNILTPDB_0_LC_8_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12293),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_8_9_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_8_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_8_9_0 (
            .in0(_gnd_net_),
            .in1(N__13635),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3D1_LC_8_9_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3D1_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3D1_LC_8_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3D1_LC_8_9_1 (
            .in0(_gnd_net_),
            .in1(N__13231),
            .in2(N__12486),
            .in3(N__12415),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIOR3DZ0Z1),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UD62_LC_8_9_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UD62_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UD62_LC_8_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UD62_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__12502),
            .in2(N__12394),
            .in3(N__12412),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI8UDZ0Z62),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIF5PB5_LC_8_9_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIF5PB5_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIF5PB5_LC_8_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIF5PB5_LC_8_9_3 (
            .in0(N__12889),
            .in1(N__12382),
            .in2(N__12487),
            .in3(N__12409),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_LC_8_9_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_LC_8_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_LC_8_9_4 (
            .in0(_gnd_net_),
            .in1(N__12514),
            .in2(_gnd_net_),
            .in3(N__12406),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PRZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_9_7.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_9_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_8_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13975),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNISG94_LC_8_10_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNISG94_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNISG94_LC_8_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 un5_visiblex_cry_7_c_RNISG94_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__13499),
            .in2(_gnd_net_),
            .in3(N__14699),
            .lcout(N_32),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DR_LC_8_10_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DR_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DR_LC_8_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DR_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__14449),
            .in2(N__12583),
            .in3(N__12385),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIC7DRZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3U41_LC_8_10_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3U41_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3U41_LC_8_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3U41_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__13314),
            .in2(N__14650),
            .in3(N__12376),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIL3UZ0Z41),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIOPOL2_LC_8_10_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIOPOL2_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIOPOL2_LC_8_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIOPOL2_LC_8_10_3 (
            .in0(N__12501),
            .in1(N__14493),
            .in2(N__13303),
            .in3(N__12508),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_LC_8_10_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_LC_8_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_LC_8_10_4 (
            .in0(N__14467),
            .in1(N__13315),
            .in2(N__14414),
            .in3(N__12505),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251),
            .ltout(font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPBZ0Z251_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_0_LC_8_10_5.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_0_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_0_LC_8_10_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIPB251_0_LC_8_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12490),
            .in3(_gnd_net_),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_10_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_8_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13500),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNISG94_0_LC_8_11_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNISG94_0_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNISG94_0_LC_8_11_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un5_visiblex_cry_7_c_RNISG94_0_LC_8_11_0 (
            .in0(_gnd_net_),
            .in1(N__13501),
            .in2(_gnd_net_),
            .in3(N__14694),
            .lcout(N_20_i),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3I1_LC_8_11_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3I1_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3I1_LC_8_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3I1_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(N__14262),
            .in2(N__14272),
            .in3(N__12445),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNICV3IZ0Z1),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPH2_LC_8_11_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPH2_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPH2_LC_8_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPH2_LC_8_11_2 (
            .in0(_gnd_net_),
            .in1(N__14179),
            .in2(N__14254),
            .in3(N__12430),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIGLPHZ0Z2),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7SRM5_LC_8_11_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7SRM5_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7SRM5_LC_8_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7SRM5_LC_8_11_3 (
            .in0(N__12599),
            .in1(N__14263),
            .in2(N__14224),
            .in3(N__12418),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_LC_8_11_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_LC_8_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFR2_LC_8_11_4 (
            .in0(_gnd_net_),
            .in1(N__14200),
            .in2(_gnd_net_),
            .in3(N__12610),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNI5HFRZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_11_5.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_11_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_8_11_5 (
            .in0(N__14695),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_11_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_11_6.LUT_INIT=16'b0000010110101111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_11_6 (
            .in0(N__14361),
            .in1(_gnd_net_),
            .in2(N__12678),
            .in3(N__12738),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_7.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_7.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_7.LUT_INIT=16'b0001000111101110;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_7 (
            .in0(N__12737),
            .in1(N__12662),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_12_0.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_12_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_2_LC_8_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13502),
            .lcout(un5_visiblex_i_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_12_2.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_12_2.LUT_INIT=16'b0011001111111111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_12_2 (
            .in0(N__13511),
            .in1(N__12656),
            .in2(_gnd_net_),
            .in3(N__14355),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i_LC_8_12_3.C_ON=1'b0;
    defparam un4_pixel_font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam un4_pixel_font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i_LC_8_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_pixel_font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i_LC_8_12_3 (
            .in0(N__14357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_axb_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_1_LC_8_12_4.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_1_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_m_1_LC_8_12_4.LUT_INIT=16'b0011001100001111;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_m_1_LC_8_12_4 (
            .in0(_gnd_net_),
            .in1(N__13607),
            .in2(N__13632),
            .in3(N__14359),
            .lcout(if_generate_plus_mult1_un47_sum_m_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_8_12_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_8_12_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_3_LC_8_12_5 (
            .in0(N__13503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_i_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_12_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_12_6.LUT_INIT=16'b1100011011111010;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_12_6 (
            .in0(N__12742),
            .in1(N__12657),
            .in2(N__12677),
            .in3(N__14358),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_12_7.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_12_7.LUT_INIT=16'b1000100010001000;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_12_7 (
            .in0(N__14356),
            .in1(N__12661),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(if_generate_plus_mult1_un47_sum_0_cry_3_ma),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNITTF6_LC_8_13_0.C_ON=1'b1;
    defparam un5_visiblex_cry_8_c_RNITTF6_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNITTF6_LC_8_13_0.LUT_INIT=16'b0011001111111111;
    LogicCell40 un5_visiblex_cry_8_c_RNITTF6_LC_8_13_0 (
            .in0(_gnd_net_),
            .in1(N__14362),
            .in2(_gnd_net_),
            .in3(N__12679),
            .lcout(N_158_0_i),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMB_LC_8_13_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMB_LC_8_13_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMB_LC_8_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMB_LC_8_13_1 (
            .in0(_gnd_net_),
            .in1(N__14619),
            .in2(_gnd_net_),
            .in3(N__12703),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4_c_RNIHUMBZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OB_LC_8_13_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OB_LC_8_13_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OB_LC_8_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OB_LC_8_13_2 (
            .in0(_gnd_net_),
            .in1(N__14631),
            .in2(N__14630),
            .in3(N__12700),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5_c_RNII0OBZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_8_13_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_8_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_8_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12697),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_8_13_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_8_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_8_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12694),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_13_6.C_ON=1'b0;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_13_6.SEQ_MODE=4'b0000;
    defparam un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_13_6.LUT_INIT=16'b0011001100111100;
    LogicCell40 un4_pixel_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_13_6 (
            .in0(N__12686),
            .in1(N__14363),
            .in2(N__13522),
            .in3(N__14696),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_LC_8_14_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_LC_8_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_LC_8_14_0 (
            .in0(_gnd_net_),
            .in1(N__14632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_LC_8_14_1.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_LC_8_14_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_LC_8_14_1 (
            .in0(_gnd_net_),
            .in1(N__12853),
            .in2(_gnd_net_),
            .in3(N__12847),
            .lcout(un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_2_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_2_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_2_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNII5M_9_LC_9_7_1.C_ON=1'b0;
    defparam beamX_RNII5M_9_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam beamX_RNII5M_9_LC_9_7_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNII5M_9_LC_9_7_1 (
            .in0(N__13556),
            .in1(N__13454),
            .in2(N__13423),
            .in3(N__13688),
            .lcout(),
            .ltout(un18_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_4_LC_9_7_2.C_ON=1'b0;
    defparam beamX_RNIVEM1_4_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_4_LC_9_7_2.LUT_INIT=16'b1101000011000000;
    LogicCell40 beamX_RNIVEM1_4_LC_9_7_2 (
            .in0(N__12840),
            .in1(N__13804),
            .in2(N__12823),
            .in3(N__13923),
            .lcout(),
            .ltout(un18_beamylt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNINAS01_10_LC_9_7_3.C_ON=1'b0;
    defparam beamX_RNINAS01_10_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam beamX_RNINAS01_10_LC_9_7_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNINAS01_10_LC_9_7_3 (
            .in0(N__13388),
            .in1(N__12820),
            .in2(N__12811),
            .in3(N__12808),
            .lcout(),
            .ltout(un15_beamy_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIMPI21_7_LC_9_7_4.C_ON=1'b0;
    defparam beamX_RNIMPI21_7_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam beamX_RNIMPI21_7_LC_9_7_4.LUT_INIT=16'b0111000001010000;
    LogicCell40 beamX_RNIMPI21_7_LC_9_7_4 (
            .in0(N__13347),
            .in1(N__12796),
            .in2(N__12790),
            .in3(N__13557),
            .lcout(un15_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_9_7_5.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_9_7_5.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_RNIR4B_9_LC_9_7_5 (
            .in0(N__13422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13455),
            .lcout(un1_beamx_2),
            .ltout(un1_beamx_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI34L6_10_LC_9_7_6.C_ON=1'b0;
    defparam beamX_RNI34L6_10_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam beamX_RNI34L6_10_LC_9_7_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNI34L6_10_LC_9_7_6 (
            .in0(N__12748),
            .in1(N__13389),
            .in2(N__12766),
            .in3(N__13558),
            .lcout(un1_beamx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI6PL_3_LC_9_7_7.C_ON=1'b0;
    defparam beamX_RNI6PL_3_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam beamX_RNI6PL_3_LC_9_7_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNI6PL_3_LC_9_7_7 (
            .in0(N__13924),
            .in1(N__13687),
            .in2(N__13810),
            .in3(N__14032),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_8_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__13759),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AA63_LC_9_8_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AA63_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AA63_LC_9_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AA63_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__12859),
            .in2(N__12873),
            .in3(N__12964),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1AAZ0Z63),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CH4_LC_9_8_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CH4_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CH4_LC_9_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CH4_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__12888),
            .in2(N__12961),
            .in3(N__12946),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIV3CHZ0Z4),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIBH1VA_LC_9_8_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIBH1VA_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIBH1VA_LC_9_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIBH1VA_LC_9_8_3 (
            .in0(N__12918),
            .in1(N__12943),
            .in2(N__12874),
            .in3(N__12931),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_LC_9_8_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_LC_9_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_LC_9_8_4 (
            .in0(_gnd_net_),
            .in1(N__12928),
            .in2(_gnd_net_),
            .in3(N__12922),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5),
            .ltout(font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AKZ0Z5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_0_LC_9_8_5.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_0_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_0_LC_9_8_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIR8AK5_0_LC_9_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12907),
            .in3(_gnd_net_),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_0_LC_9_8_6.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_0_LC_9_8_6.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_0_LC_9_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIT8PR2_0_LC_9_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12887),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_8_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_8_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_9_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13633),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_9_9_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(N__13164),
            .in2(N__13119),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_9_9_1.C_ON=1'b1;
    defparam beamX_2_LC_9_9_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_9_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(N__14119),
            .in2(_gnd_net_),
            .in3(N__13000),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_9_9_2.C_ON=1'b1;
    defparam beamX_3_LC_9_9_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_9_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__14025),
            .in2(_gnd_net_),
            .in3(N__12997),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_9_9_3.C_ON=1'b1;
    defparam beamX_4_LC_9_9_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_9_9_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_9_9_3 (
            .in0(N__13293),
            .in1(N__13916),
            .in2(_gnd_net_),
            .in3(N__12994),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_9_9_4.C_ON=1'b1;
    defparam beamX_5_LC_9_9_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_9_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(N__13800),
            .in2(_gnd_net_),
            .in3(N__12991),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_9_9_5.C_ON=1'b1;
    defparam beamX_6_LC_9_9_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_9_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(N__13679),
            .in2(_gnd_net_),
            .in3(N__12988),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_9_9_6.C_ON=1'b1;
    defparam beamX_7_LC_9_9_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_9_9_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(N__13554),
            .in2(_gnd_net_),
            .in3(N__12985),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_9_9_7.C_ON=1'b1;
    defparam beamX_8_LC_9_9_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_9_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(N__13450),
            .in2(_gnd_net_),
            .in3(N__12982),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__13223),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_9_10_0.C_ON=1'b1;
    defparam beamX_9_LC_9_10_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_9_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(N__13417),
            .in2(_gnd_net_),
            .in3(N__12979),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__13224),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_9_10_1.C_ON=1'b0;
    defparam beamX_10_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_9_10_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_9_10_1 (
            .in0(N__13384),
            .in1(N__13291),
            .in2(_gnd_net_),
            .in3(N__12976),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13224),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_9_10_2.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_9_10_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNI5457_5_LC_9_10_2 (
            .in0(N__13360),
            .in1(N__13546),
            .in2(N__13351),
            .in3(N__13799),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9TH9_LC_9_10_3.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9TH9_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9TH9_LC_9_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9TH9_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14448),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9),
            .ltout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9THZ0Z9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38L_LC_9_10_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38L_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38L_LC_9_10_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38L_LC_9_10_4 (
            .in0(N__14494),
            .in1(_gnd_net_),
            .in2(N__13306),
            .in3(_gnd_net_),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH38LZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_9_10_5.C_ON=1'b0;
    defparam beamX_0_LC_9_10_5.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_9_10_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_0_LC_9_10_5 (
            .in0(_gnd_net_),
            .in1(N__13290),
            .in2(_gnd_net_),
            .in3(N__13165),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13224),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_9_10_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_9_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13510),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_9_10_7.C_ON=1'b0;
    defparam beamX_1_LC_9_10_7.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_9_10_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_9_10_7 (
            .in0(_gnd_net_),
            .in1(N__13113),
            .in2(_gnd_net_),
            .in3(N__13166),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13224),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_9_11_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_9_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13167),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_9_11_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_9_11_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13114),
            .in3(N__13003),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_9_11_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_9_11_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14127),
            .in3(N__14041),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_9_11_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_9_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(N__14593),
            .in2(N__14036),
            .in3(N__13930),
            .lcout(un1_visiblex_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_9_11_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_9_11_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13926),
            .in3(N__13813),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_9_11_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_9_11_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_9_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13809),
            .in3(N__13696),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_9_11_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_9_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_9_11_6 (
            .in0(_gnd_net_),
            .in1(N__14594),
            .in2(N__13689),
            .in3(N__13561),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_9_11_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_9_11_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_9_11_7 (
            .in0(_gnd_net_),
            .in1(N__13555),
            .in2(_gnd_net_),
            .in3(N__13459),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_9_12_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_9_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_9_12_0 (
            .in0(_gnd_net_),
            .in1(N__14595),
            .in2(N__13456),
            .in3(N__13426),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_9_12_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_9_12_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_9_12_1 (
            .in0(_gnd_net_),
            .in1(N__13418),
            .in2(_gnd_net_),
            .in3(N__13393),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_12_5.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_1_LC_9_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14698),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_0_LC_9_12_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_0_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_0_LC_9_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_0_LC_9_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14174),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_13_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_13_0 (
            .in0(_gnd_net_),
            .in1(N__14697),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UP11_LC_9_13_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UP11_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UP11_LC_9_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UP11_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(N__14136),
            .in2(N__14158),
            .in3(N__14239),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI2UPZ0Z11),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBB1_LC_9_13_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBB1_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBB1_LC_9_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBB1_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(N__14148),
            .in2(N__14236),
            .in3(N__14212),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIJHBBZ0Z1),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_c_RNICFTM2_LC_9_13_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_c_RNICFTM2_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_c_RNICFTM2_LC_9_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_c_RNICFTM2_LC_9_13_3 (
            .in0(N__14175),
            .in1(N__14137),
            .in2(N__14209),
            .in3(N__14191),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_LC_9_13_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_LC_9_13_4.LUT_INIT=16'b0110011010011001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFB1_LC_9_13_4 (
            .in0(N__14188),
            .in1(N__14149),
            .in2(_gnd_net_),
            .in3(N__14182),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNINPFBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_13_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_9_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14370),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_0_LC_9_13_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_0_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_0_LC_9_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un33_sum_cry_6_c_RNI9UBH_0_LC_9_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14147),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_11_12_0.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_11_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_11_12_0 (
            .in0(_gnd_net_),
            .in1(N__14700),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LB_LC_11_12_1.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LB_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LB_LC_11_12_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LB_LC_11_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14281),
            .in3(N__14635),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNI74LBZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MB_LC_11_12_2.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MB_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MB_LC_11_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MB_LC_11_12_2 (
            .in0(_gnd_net_),
            .in1(N__14623),
            .in2(N__14431),
            .in3(N__14470),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNI86MBZ0),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_11_12_3.C_ON=1'b1;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_11_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_11_12_3 (
            .in0(_gnd_net_),
            .in1(N__14376),
            .in2(_gnd_net_),
            .in3(N__14455),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_11_12_4.C_ON=1'b0;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_11_12_4.SEQ_MODE=4'b0000;
    defparam font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_11_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_11_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14452),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_11_12_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_11_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14375),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_12_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_12_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_11_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_2_LC_11_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14374),
            .lcout(font_un13_pixel_if_generate_plus_mult1_un26_sum_s_2_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
