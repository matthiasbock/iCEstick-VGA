-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 24 2015 19:05:04

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSync : out std_logic;
    SCLK1 : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic;
    nCS2 : out std_logic;
    SDATA2 : out std_logic;
    SCLK2 : out std_logic;
    Clock12MHz : in std_logic;
    nCS1 : out std_logic;
    SDATA1 : in std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_1_0_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6 : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \beamY_RNITSR8_0Z0Z_8\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\ : std_logic;
signal \beamY_RNISI4A_0Z0Z_9\ : std_logic;
signal \beamY_RNIE925Z0Z_6_cascade_\ : std_logic;
signal \beamY_RNIKOP3_0Z0Z_6\ : std_logic;
signal \un5_visibley_c2_cascade_\ : std_logic;
signal un5_visibley_c6_0_0_0 : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal un20_beamy_cry_1 : std_logic;
signal un20_beamy_cry_2 : std_logic;
signal un20_beamy_cry_3 : std_logic;
signal un20_beamy_cry_4 : std_logic;
signal un20_beamy_cry_5 : std_logic;
signal un20_beamy_cry_6 : std_logic;
signal un20_beamy_cry_7 : std_logic;
signal un20_beamy_cry_8 : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc5_0_x1 : std_logic;
signal \if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal un1_voltage_0_cry_0 : std_logic;
signal un1_voltage_0_cry_1 : std_logic;
signal un1_voltage_0_cry_2 : std_logic;
signal \N_1503_cascade_\ : std_logic;
signal \SDATA1_ibuf_RNILOUGZ0Z2\ : std_logic;
signal \un1_voltage_1_1_axb_0_cascade_\ : std_logic;
signal \voltage_0_1_sqmuxa_1_cascade_\ : std_logic;
signal \voltage_3_9_iv_0_0_cascade_\ : std_logic;
signal \N_1507\ : std_logic;
signal \N_1507_cascade_\ : std_logic;
signal \voltage_3_RNO_0Z0Z_0\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal un1_voltage_3_1_cry_0 : std_logic;
signal un1_voltage_3_1_cry_1 : std_logic;
signal un1_voltage_3_1_cry_2 : std_logic;
signal \ScreenBuffer_0_0_1_sqmuxa\ : std_logic;
signal \un4_voltage_2_0__N_13_mux_iZ0_cascade_\ : std_logic;
signal \SDATA1_ibuf_RNI098KZ0Z2\ : std_logic;
signal \N_35_0_i_cascade_\ : std_logic;
signal \un4_voltage_10_9__N_4_cascade_\ : std_logic;
signal \un4_voltage_2_0__N_5_iZ0\ : std_logic;
signal \voltage_0_1_sqmuxa_cascade_\ : std_logic;
signal \un1_voltage_0_cry_0_0_c_RNOZ0\ : std_logic;
signal \N_34_0_i\ : std_logic;
signal \N_41_i\ : std_logic;
signal \N_41_i_cascade_\ : std_logic;
signal voltage_0_1_sqmuxa : std_logic;
signal \ScreenBuffer_0_1_1_sqmuxa_2\ : std_logic;
signal \un4_voltage_2_0__i2_mux\ : std_logic;
signal \bfn_2_1_0_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_\ : std_logic;
signal \un5_visibley_axbxc7_1_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un33_sum_axb3_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz : std_logic;
signal \chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_\ : std_logic;
signal \beamY_RNI9425_0Z0Z_6_cascade_\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_\ : std_logic;
signal \beamY_RNI9425Z0Z_6_cascade_\ : std_logic;
signal if_generate_plus_mult1_un61_sum_ac0_x0 : std_logic;
signal if_generate_plus_mult1_un61_sum_ac0_x1 : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_ac0_6 : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_c4_d : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_\ : std_logic;
signal \beamY_RNI75QM4Z0Z_5_cascade_\ : std_logic;
signal if_generate_plus_mult1_un68_sum_axbxc5_x0 : std_logic;
signal \if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8\ : std_logic;
signal if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0 : std_logic;
signal \if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_\ : std_logic;
signal \beamY_RNI75QM4Z0Z_5\ : std_logic;
signal \voltage_0_10_iv_0_2_cascade_\ : std_logic;
signal \voltage_0_RNO_0Z0Z_2\ : std_logic;
signal \voltage_1_9_iv_0_2_cascade_\ : std_logic;
signal \voltage_3_RNO_0Z0Z_2\ : std_logic;
signal \voltage_3_9_iv_0_2_cascade_\ : std_logic;
signal \CO2_3_cascade_\ : std_logic;
signal \N_1155_cascade_\ : std_logic;
signal voltage_0_10_iv_0_3 : std_logic;
signal \N_1519\ : std_logic;
signal \N_1521\ : std_logic;
signal \counter_RNI49LH1_0Z0Z_0\ : std_logic;
signal voltage_1_9_iv_0_0 : std_logic;
signal \CO1_3\ : std_logic;
signal \voltage_2_1_sqmuxa_cascade_\ : std_logic;
signal \N_1155\ : std_logic;
signal voltage_1_1_sqmuxa : std_logic;
signal \voltage_1_1_sqmuxa_cascade_\ : std_logic;
signal voltage_1_9_iv_0_3 : std_logic;
signal \voltage_3_RNO_0Z0Z_3\ : std_logic;
signal voltage_3_9_iv_0_3 : std_logic;
signal \N_1510\ : std_logic;
signal \N_1506_cascade_\ : std_logic;
signal \counter_RNIGLLH1Z0Z_0_cascade_\ : std_logic;
signal \N_2063\ : std_logic;
signal \N_1522\ : std_logic;
signal \un1_voltage_1_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \counter_RNILOUG2Z0Z_3\ : std_logic;
signal un1_voltage_1_1_cry_0 : std_logic;
signal \counter_RNIT58K2Z0Z_2\ : std_logic;
signal \voltage_1_RNO_0Z0Z_2\ : std_logic;
signal un1_voltage_1_1_cry_1 : std_logic;
signal un1_voltage_1_1_cry_2 : std_logic;
signal \voltage_1_RNO_0Z0Z_3\ : std_logic;
signal \un6_slaveselectlto9_1_cascade_\ : std_logic;
signal \un6_slaveselect_0_cascade_\ : std_logic;
signal un3_slaveselectlt9 : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \voltage_2_RNIKG123Z0Z_1\ : std_logic;
signal un1_voltage_2_1_cry_0 : std_logic;
signal \counter_RNI2RBA2Z0Z_3\ : std_logic;
signal un1_voltage_2_1_cry_1 : std_logic;
signal un1_voltage_2_1_axb_3 : std_logic;
signal voltage_2_9_iv_0_3 : std_logic;
signal un1_voltage_2_1_cry_2 : std_logic;
signal \N_46_1\ : std_logic;
signal \un1_sclk17_2_1_cascade_\ : std_logic;
signal \un1_sclk17_1_1_cascade_\ : std_logic;
signal \bfn_4_1_0_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal \bfn_4_2_0_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0 : std_logic;
signal un5_visibley_c2 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_\ : std_logic;
signal \beamY_RNIEDF31Z0Z_6\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c4_3_1 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_6_2 : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0 : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0\ : std_logic;
signal \beamY_RNIFS4TZ0Z_7\ : std_logic;
signal \beamY_RNIFS4TZ0Z_7_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_\ : std_logic;
signal \beamY_RNIQTGS2Z0Z_8_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axb3_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0 : std_logic;
signal \beamY_RNIQTGS2Z0Z_8\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_c4 : std_logic;
signal \beamY_RNI0K169Z0Z_6_cascade_\ : std_logic;
signal un5_visibley_0_29 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_\ : std_logic;
signal \if_m1_x1_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_c5 : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_axb4_i : std_logic;
signal if_m1_x0 : std_logic;
signal \un113_pixel_3_0_11__g1_0\ : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_\ : std_logic;
signal \GB_BUFFER_Clock12MHz_c_g_THRU_CO\ : std_logic;
signal \N_1159_i\ : std_logic;
signal \N_1154\ : std_logic;
signal \N_1159_i_cascade_\ : std_logic;
signal voltage_2_1_sqmuxa : std_logic;
signal voltage_0_0_sqmuxa_1 : std_logic;
signal \slaveselect_RNILOQC2Z0Z_1\ : std_logic;
signal \slaveselect_RNILOQC2Z0Z_1_cascade_\ : std_logic;
signal \counter_RNICHLH1Z0Z_0\ : std_logic;
signal \un1_voltage_012_0_cascade_\ : std_logic;
signal un74_voltage_0 : std_logic;
signal \N_1153\ : std_logic;
signal voltage_0_1_sqmuxa_1 : std_logic;
signal \N_1153_cascade_\ : std_logic;
signal voltage_3_1_sqmuxa : std_logic;
signal \voltage_3_RNO_0Z0Z_1\ : std_logic;
signal \voltage_3_9_iv_0_1_cascade_\ : std_logic;
signal un1_voltage_012_0 : std_logic;
signal voltage_1_9_iv_0_1 : std_logic;
signal \voltage_1_RNO_0Z0Z_1\ : std_logic;
signal \N_1504_cascade_\ : std_logic;
signal \N_1504\ : std_logic;
signal \counter_RNI8DLH1Z0Z_0\ : std_logic;
signal \N_1508\ : std_logic;
signal \slaveselect_RNILOQC2Z0Z_2\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal counter_cry_1 : std_logic;
signal counter_cry_2 : std_logic;
signal counter_cry_3 : std_logic;
signal counter_cry_4 : std_logic;
signal counter_cry_5 : std_logic;
signal counter_cry_6 : std_logic;
signal counter_cry_7 : std_logic;
signal counter_cry_8 : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal un1_counter_i_0 : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_\ : std_logic;
signal chessboardpixel_un173_pixellt10 : std_logic;
signal chessboardpixel_un151_pixel_27 : std_logic;
signal \chessboardpixel_un177_pixel_26_cascade_\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0\ : std_logic;
signal \un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_\ : std_logic;
signal chessboardpixel_un199_pixellt10 : std_logic;
signal \un113_pixel_4_0_15__un1_beamylto9_3\ : std_logic;
signal \VSync_c\ : std_logic;
signal \un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_\ : std_logic;
signal \beamY_RNII8O41Z0Z_9\ : std_logic;
signal \un113_pixel_4_0_15__g0_i_a3_0Z0Z_4\ : std_logic;
signal if_m1_5 : std_logic;
signal \if_generate_plus_mult1_un54_sum_axbxc5_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\ : std_logic;
signal if_generate_plus_mult1_un75_sum_ac0_5_x1 : std_logic;
signal \row_1_if_i2_mux_0_cascade_\ : std_logic;
signal if_generate_plus_mult1_un75_sum_ac0_5_x0 : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_\ : std_logic;
signal un5_visibley_c5 : std_logic;
signal \beamY_RNIJNLCZ0Z_9\ : std_logic;
signal \beamY_RNIJNLCZ0Z_9_cascade_\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal \beamY_RNIVGU01Z0Z_9\ : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0 : std_logic;
signal row_1_if_generate_plus_mult1_un75_sum_ac0_5 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum : std_logic;
signal if_generate_plus_mult1_un75_sum_c5_x0 : std_logic;
signal \if_generate_plus_mult1_un75_sum_c5_x1_cascade_\ : std_logic;
signal \beamY_RNIPNEA3_0Z0Z_6\ : std_logic;
signal \beamY_RNI0K169Z0Z_6\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c4 : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9\ : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_c5_N_9\ : std_logic;
signal \beamY_RNIPLAE31Z0Z_4_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0 : std_logic;
signal \beamY_RNIV42D31_0Z0Z_6\ : std_logic;
signal \un113_pixel_3_0_11__N_4_i_0\ : std_logic;
signal g1_0_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb3 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum : std_logic;
signal \beamY_RNIV42D31Z0Z_6\ : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axbxc5_0 : std_logic;
signal \un113_pixel_3_0_11__g0_0_x2_0Z0Z_0\ : std_logic;
signal \un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0\ : std_logic;
signal \N_1520\ : std_logic;
signal \un1_voltage_2_1_cry_0_c_RNOZ0\ : std_logic;
signal voltage_2_9_iv_0_0 : std_logic;
signal \un1_voltage_2_1_axb_0_cascade_\ : std_logic;
signal voltage_2_9_iv_0_2 : std_logic;
signal \voltage_2_RNO_0Z0Z_2\ : std_logic;
signal un1_voltage_012_3_0 : std_logic;
signal voltage_2_9_iv_0_1 : std_logic;
signal \voltage_2_RNO_0Z0Z_1\ : std_logic;
signal \un42_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal un42_cry_1 : std_logic;
signal \counter_RNIGLLH1Z0Z_0\ : std_logic;
signal un42_cry_2 : std_logic;
signal voltage_011_0 : std_logic;
signal un42_cry_3 : std_logic;
signal voltage_011 : std_logic;
signal \ScreenBuffer_1_122_1_cascade_\ : std_logic;
signal \ScreenBuffer_1_3_1_sqmuxa\ : std_logic;
signal \ScreenBuffer_1_0_1_sqmuxa\ : std_logic;
signal \Z_decfrac4\ : std_logic;
signal \un1_sclk17_0_0_cascade_\ : std_logic;
signal un39_0_3 : std_logic;
signal \un39_0_3_cascade_\ : std_logic;
signal un5_slaveselect_1 : std_logic;
signal \un5_slaveselect_1_cascade_\ : std_logic;
signal \ScreenBuffer_1_122_1\ : std_logic;
signal un39_0_6 : std_logic;
signal \ScreenBuffer_1_2_1_sqmuxa\ : std_logic;
signal \ScreenBuffer_1_2_1_sqmuxa_cascade_\ : std_logic;
signal un10_slaveselect : std_logic;
signal \slaveselect_RNILOQC2Z0Z_0_cascade_\ : std_logic;
signal \Z_decfrac4_2\ : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \un1_counter_1lto9_2_cascade_\ : std_logic;
signal un10_slaveselectlt4 : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal un1_counter_1lt9 : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal slaveselect_1lto9_4 : std_logic;
signal slaveselect_1lto9_3 : std_logic;
signal \SCLK1_0_i\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum : std_logic;
signal \un113_pixel_4_0_15__un5_beamx_2Z0Z_0\ : std_logic;
signal \un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_\ : std_logic;
signal un5_beamx_0 : std_logic;
signal \un5_beamx_0_cascade_\ : std_logic;
signal \un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_\ : std_logic;
signal un13_beamylt6_0 : std_logic;
signal \un13_beamylt6_0_cascade_\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \un113_pixel_4_0_15__un4_rowZ0Z_2\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axbxc5 : std_logic;
signal \r_N_6\ : std_logic;
signal \un113_pixel_4_0_15__un3_beamxZ0Z_7\ : std_logic;
signal \un1_beamxlt10_0_cascade_\ : std_logic;
signal \HSync_c\ : std_logic;
signal un18_beamylt10_0 : std_logic;
signal if_generate_plus_mult1_un82_sum_axbxc5_0_x1 : std_logic;
signal if_generate_plus_mult1_un82_sum_axbxc5_0_x0 : std_logic;
signal un1_beamy_4 : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal \un113_pixel_4_0_15__un4_rowZ0Z_5\ : std_logic;
signal un13_beamy_0 : std_logic;
signal chessboardpixel_un174_pixel : std_logic;
signal \un4_row_cascade_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un4_beamylt8_0 : std_logic;
signal un4_beamy_0 : std_logic;
signal \un113_pixel_4_0_15__un8_beamylto9Z0Z_1\ : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal un8_beamy : std_logic;
signal \N_6_i\ : std_logic;
signal \N_6_i_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un4_beamylt6 : std_logic;
signal if_m1_ns : std_logic;
signal \if_m2_2_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un82_sum_axbxc5_0 : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_i : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\ : std_logic;
signal \voltage_2Z0Z_0\ : std_logic;
signal \voltage_1Z0Z_0\ : std_logic;
signal \voltage_2Z0Z_2\ : std_logic;
signal \voltage_1Z0Z_2\ : std_logic;
signal \voltage_2Z0Z_3\ : std_logic;
signal \voltage_1Z0Z_3\ : std_logic;
signal \voltage_2Z0Z_1\ : std_logic;
signal \voltage_1Z0Z_1\ : std_logic;
signal \un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0\ : std_logic;
signal \N_1505\ : std_logic;
signal \N_1509\ : std_logic;
signal \un42_cry_2_c_RNOZ0\ : std_logic;
signal \un1_sclk17_6_1_cascade_\ : std_logic;
signal \un1_sclk17_3_1_cascade_\ : std_logic;
signal \ScreenBuffer_0_0_1_sqmuxa_0\ : std_logic;
signal \slaveselect_RNILOQCZ0Z2\ : std_logic;
signal \un1_sclk17_8_0_0_cascade_\ : std_logic;
signal \voltage_3Z0Z_2\ : std_logic;
signal \voltage_0Z0Z_2\ : std_logic;
signal un1_sclk17_7_1 : std_logic;
signal un5_slaveselect : std_logic;
signal \SDATA2_c\ : std_logic;
signal \un1_sclk17_9_1_cascade_\ : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal un1_sclk17_4_1 : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_i_5 : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \un113_pixel_4_0_15__un18_beamylto9Z0Z_2\ : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal un1_beamx_2 : std_logic;
signal charx_i_24 : std_logic;
signal \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\ : std_logic;
signal \font_un3_pixel_28_cascade_\ : std_logic;
signal \un113_pixel_4_0_15__un15_beamyZ0Z_2\ : std_logic;
signal un13_beamy : std_logic;
signal \font_un61_pixel_cascade_\ : std_logic;
signal un4_row : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf : std_logic;
signal charx_23 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\ : std_logic;
signal charx_if_generate_plus_mult1_un1_sum_axb1 : std_logic;
signal \N_9_i_cascade_\ : std_logic;
signal \N_13_0\ : std_logic;
signal \ScreenBuffer_0_8Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_0Z0Z_0\ : std_logic;
signal \currentchar_1_9_ns_1_0_cascade_\ : std_logic;
signal \ScreenBuffer_1_1Z0Z_0\ : std_logic;
signal \currentchar_1_6_ns_1_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_1Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_0Z0Z_4\ : std_logic;
signal \ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_\ : std_logic;
signal \ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_cZ0Z4\ : std_logic;
signal row_1_if_generate_plus_mult1_un75_sum_axbxc5_0 : std_logic;
signal \ScreenBuffer_1_2Z0Z_0\ : std_logic;
signal \un3_rowlto1_cascade_\ : std_logic;
signal \ScreenBuffer_0_2Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_1_1_sqmuxa\ : std_logic;
signal \ScreenBuffer_0_0Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_1Z0Z_4\ : std_logic;
signal \ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_\ : std_logic;
signal currentchar_1_11_ns_1_4 : std_logic;
signal \ScreenBuffer_1_2_RNIUP6F2FZ0Z_4\ : std_logic;
signal \ScreenBuffer_1_3Z0Z_4\ : std_logic;
signal \ScreenBuffer_1_3_RNIVS9G2FZ0Z_4\ : std_logic;
signal \g1Z0Z_1_cascade_\ : std_logic;
signal \N_1428_0_cascade_\ : std_logic;
signal \un113_pixel_4_0_15__g1_1_cascade_\ : std_logic;
signal \N_1300_0\ : std_logic;
signal \un112_pixel_0_2_cascade_\ : std_logic;
signal \N_1293_0\ : std_logic;
signal \slaveselect_RNILOQC2Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_2Z0Z_4\ : std_logic;
signal \ScreenBuffer_1_3Z0Z_2\ : std_logic;
signal \ScreenBuffer_1_0Z0Z_2\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_\ : std_logic;
signal m10_0_x1 : std_logic;
signal \un112_pixel_2_2_cascade_\ : std_logic;
signal \un113_pixel_3_0_11__g0_0Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_7_RNIHMH43T2Z0Z_0\ : std_logic;
signal \beamY_RNIDQUNU91Z0Z_0_cascade_\ : std_logic;
signal \un115_pixel_2_sn_5_cascade_\ : std_logic;
signal \un112_pixel_7_cascade_\ : std_logic;
signal \beamY_RNIINK7J73Z0Z_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal un3_beamx_0 : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \CO3_0_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_s_2_sf : std_logic;
signal chary_if_generate_plus_mult1_un33_sum_axb3 : std_logic;
signal chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3 : std_logic;
signal \N_13\ : std_logic;
signal \un113_pixel_4_0_15__un4_rowZ0Z_1\ : std_logic;
signal un1_voltage_0_axb_0 : std_logic;
signal voltage_0_10_iv_0_0 : std_logic;
signal un1_voltage_012_2_0 : std_logic;
signal voltage_0_10_iv_0_1 : std_logic;
signal \voltage_0_RNO_0Z0Z_1\ : std_logic;
signal \nCS1_c\ : std_logic;
signal un1_counter_1_0 : std_logic;
signal voltage_0_0_sqmuxa_1_g : std_logic;
signal \voltage_3Z0Z_0\ : std_logic;
signal \voltage_0Z0Z_0\ : std_logic;
signal \un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal chary_24 : std_logic;
signal \un113_pixel_4_0_15__gZ0Z2\ : std_logic;
signal font_un3_pixel_30 : std_logic;
signal \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1\ : std_logic;
signal \font_un57_pixel_cascade_\ : std_logic;
signal currentchar_1_5 : std_logic;
signal font_un67_pixel_ac0_5 : std_logic;
signal font_un64_pixel_ac0_5 : std_logic;
signal \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_\ : std_logic;
signal \N_12\ : std_logic;
signal \un113_pixel_4_0_15__g0_iZ0Z_2\ : std_logic;
signal \un113_pixel_4_0_15__g0_iZ0Z_5_cascade_\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6\ : std_logic;
signal \beamY_RNIOEPPEK1Z0Z_0_cascade_\ : std_logic;
signal un112_pixel_1_2 : std_logic;
signal \N_3461_0_cascade_\ : std_logic;
signal \N_4568_0_cascade_\ : std_logic;
signal \N_1305_0\ : std_logic;
signal \un113_pixel_4_0_15__g0_0Z0Z_2\ : std_logic;
signal \Pixel_3_sqmuxa_0\ : std_logic;
signal g0_1_1 : std_logic;
signal \N_1_0_cascade_\ : std_logic;
signal \ScreenBuffer_1_3Z0Z_3\ : std_logic;
signal \ScreenBuffer_1_1Z0Z_3\ : std_logic;
signal \ScreenBuffer_1_2Z0Z_3\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_N_13_cascade_\ : std_logic;
signal \voltage_3Z0Z_3\ : std_logic;
signal \voltage_0Z0Z_3\ : std_logic;
signal \ScreenBuffer_1_0Z0Z_3\ : std_logic;
signal \un113_pixel_4_0_15__g0_1Z0Z_0\ : std_logic;
signal \un113_pixel_4_0_15__g0_3_0\ : std_logic;
signal \voltage_3Z0Z_1\ : std_logic;
signal \slaveselectZ0\ : std_logic;
signal \voltage_0Z0Z_1\ : std_logic;
signal \un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0\ : std_logic;
signal \ScreenBuffer_0_12Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_4Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_6Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_\ : std_logic;
signal \currentchar_m7_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_7Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_5Z0Z_0\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_N_13\ : std_logic;
signal un112_pixel_1_2_x1 : std_logic;
signal \un112_pixel_2_8_cascade_\ : std_logic;
signal un115_pixel_4_am_7 : std_logic;
signal \N_1287_cascade_\ : std_logic;
signal \currentchar_1_0_cascade_\ : std_logic;
signal un115_pixel_4_bm_7 : std_logic;
signal \ScreenBuffer_0_7_RNII0GVLQZ0Z_0\ : std_logic;
signal \un113_pixel_1_0_3__N_10_mux_cascade_\ : std_logic;
signal \N_1285_0_0_0_cascade_\ : std_logic;
signal \un113_pixel_3_0_11__g1_0_0_0\ : std_logic;
signal m14 : std_logic;
signal \m14_cascade_\ : std_logic;
signal \beamY_RNI7RM4IFZ0Z_0\ : std_logic;
signal \un113_pixel_3_0_11__g1_1_0\ : std_logic;
signal \beamY_RNIPQEDM42Z0Z_0\ : std_logic;
signal \N_1293\ : std_logic;
signal \N_1306_cascade_\ : std_logic;
signal \N_1327_0\ : std_logic;
signal \m11_cascade_\ : std_logic;
signal \un113_pixel_4_0_15__N_17\ : std_logic;
signal \un115_pixel_6_bm_2_cascade_\ : std_logic;
signal \N_1330\ : std_logic;
signal un115_pixel_6_am_2 : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_1 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx : std_logic;
signal if_generate_plus_mult1_un47_sum_0_cry_3_ma : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_2 : std_logic;
signal \N_1184_0_i\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_4 : std_logic;
signal un5_visiblex_i_25 : std_logic;
signal \N_2110_i_cascade_\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_5 : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_3 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_2 : std_logic;
signal \SDATA1_c\ : std_logic;
signal un1_sclk17_9_0_3 : std_logic;
signal un1_sclk17_5_1_0 : std_logic;
signal \ScreenBuffer_0_9Z0Z_0\ : std_logic;
signal \Clock12MHz_c_g\ : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_4 : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_2_l_fx : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_3_l_fx : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_4_l_fx : std_logic;
signal \N_2110_i\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \if_generate_plus_mult1_un54_sum_s_5_cascade_\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \N_2096_i\ : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal column_1_i_i_3 : std_logic;
signal \N_11\ : std_logic;
signal \un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0\ : std_logic;
signal \un113_pixel_4_0_15__g0_i_a3_2\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \un113_pixel_7_1_7__g0_6Z0Z_0\ : std_logic;
signal \N_3078_0\ : std_logic;
signal \N_1297_0_cascade_\ : std_logic;
signal font_un67_pixel_ac0_5_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c5 : std_logic;
signal chary_if_generate_plus_mult1_un1_sum_axbxc3_2 : std_logic;
signal \un113_pixel_4_0_15__g0_4_0Z0Z_0\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i\ : std_logic;
signal \un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_\ : std_logic;
signal font_un3_pixel_28 : std_logic;
signal \N_1342\ : std_logic;
signal \un113_pixel_4_0_15__g0_5Z0Z_1\ : std_logic;
signal font_un71_pixellt7_0_1 : std_logic;
signal font_un64_pixel_ac0_5_0 : std_logic;
signal \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3\ : std_logic;
signal font_un3_pixel_0_29 : std_logic;
signal \un113_pixel_4_0_15__g0_5Z0Z_4_cascade_\ : std_logic;
signal \N_9\ : std_logic;
signal \un113_pixel_4_0_15__g2Z0Z_0_cascade_\ : std_logic;
signal \N_4566_0\ : std_logic;
signal un115_pixel_4 : std_logic;
signal \N_4564_0\ : std_logic;
signal \N_5_0\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1\ : std_logic;
signal \N_4561_0\ : std_logic;
signal g1_0 : std_logic;
signal \N_2075\ : std_logic;
signal \un115_pixel_2_s_6_cascade_\ : std_logic;
signal \un115_pixel_2_d_0_6_cascade_\ : std_logic;
signal un115_pixel_3_bm_6 : std_logic;
signal \ScreenBuffer_1_2Z0Z_1\ : std_logic;
signal \ScreenBuffer_1_0Z0Z_1\ : std_logic;
signal \N_1_7_0\ : std_logic;
signal \ScreenBuffer_1_3Z0Z_1\ : std_logic;
signal \ScreenBuffer_1_1Z0Z_1\ : std_logic;
signal m8 : std_logic;
signal \ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_\ : std_logic;
signal \un113_pixel_3_0_11__gZ0Z1\ : std_logic;
signal un115_pixel_5_s_7 : std_logic;
signal \un115_pixel_5_am_7_cascade_\ : std_logic;
signal un115_pixel_5_bm_7 : std_logic;
signal \N_1288\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\ : std_logic;
signal \un113_pixel_4_0_15__g1Z0Z_0\ : std_logic;
signal m9 : std_logic;
signal \m9_cascade_\ : std_logic;
signal m6 : std_logic;
signal \m6_cascade_\ : std_logic;
signal \beamY_RNICJUESD2Z0Z_0\ : std_logic;
signal \N_1286_0_0_0\ : std_logic;
signal \N_1289\ : std_logic;
signal font_un3_pixel_29 : std_logic;
signal \N_4562_0_0_0_cascade_\ : std_logic;
signal \N_1340_0\ : std_logic;
signal \beamY_RNICJUESD2_0Z0Z_0\ : std_logic;
signal \beamY_RNI1H36941Z0Z_0\ : std_logic;
signal font_un125_pixel_1_bm : std_logic;
signal \un113_pixel_6_1_5__N_11_cascade_\ : std_logic;
signal \un113_pixel_2_0_3__N_8\ : std_logic;
signal \beamY_RNICJUESD2_2Z0Z_0\ : std_logic;
signal m17 : std_logic;
signal m12 : std_logic;
signal un115_pixel_5_ns_x1_0 : std_logic;
signal un115_pixel_5_ns_x0_0 : std_logic;
signal \N_1325_cascade_\ : std_logic;
signal un115_pixel_7_bm_0 : std_logic;
signal \N_1315_cascade_\ : std_logic;
signal \N_1322\ : std_logic;
signal \N_1329\ : std_logic;
signal \N_1294_cascade_\ : std_logic;
signal \beamY_RNICJUESD2_1Z0Z_0\ : std_logic;
signal \N_1308\ : std_logic;
signal un115_pixel_5_d_2 : std_logic;
signal \un113_pixel_1_0_3__N_10_mux\ : std_logic;
signal \beamY_RNIMR86ES2Z0Z_0\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\ : std_logic;
signal chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_2 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_2 : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_3 : std_logic;
signal \un5_visiblex_cry_7_c_RNIVZ0Z952\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_5 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum : std_logic;
signal un5_visiblex_i_0_25 : std_logic;
signal \N_56\ : std_logic;
signal \N_32_i\ : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx : std_logic;
signal \CO3_0\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_axb_3_i : std_logic;
signal charx_if_generate_plus_mult1_un54_sum : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal column_1_i_i_2 : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un75_sum_axb_4_l_fx : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un6_rowlt7_0 : std_logic;
signal chessboardpixel_un151_pixel_24 : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal un3_rowlto0 : std_logic;
signal \un113_pixel_3_0_11__currentchar_m7_0Z0Z_1\ : std_logic;
signal \d_N_3_mux_cascade_\ : std_logic;
signal \ScreenBuffer_1_2Z0Z_2\ : std_logic;
signal \ScreenBuffer_1_1Z0Z_2\ : std_logic;
signal \un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2\ : std_logic;
signal \ScreenBuffer_0_10Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_11Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_3Z0Z_0\ : std_logic;
signal \currentchar_1_5_ns_1_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_3Z0Z_0\ : std_logic;
signal \beamY_RNIVDIFFI1Z0Z_0\ : std_logic;
signal \beamY_RNI2RNL4M2Z0Z_0\ : std_logic;
signal un3_rowlto1 : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\ : std_logic;
signal \N_52\ : std_logic;
signal un112_pixel_2_8 : std_logic;
signal \N_4581_0_cascade_\ : std_logic;
signal \N_1296_0_cascade_\ : std_logic;
signal \N_1296_0\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \N_1303_0\ : std_logic;
signal \g0_16_x0_cascade_\ : std_logic;
signal g0_16_x1 : std_logic;
signal \N_4560_0\ : std_logic;
signal \N_1309_0\ : std_logic;
signal \un113_pixel_4_0_15__N_2\ : std_logic;
signal \un113_pixel_7_1_7__N_9\ : std_logic;
signal \beamY_RNIJIDRG11Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNIJIDRG11_0Z0Z_0\ : std_logic;
signal \beamY_RNIRG0LHO1Z0Z_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_7_RNIB3R6U63Z0Z_0\ : std_logic;
signal font_un28_pixel_29 : std_logic;
signal \beamY_RNIRG0LHO1Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0\ : std_logic;
signal \g0_2_x1_cascade_\ : std_logic;
signal g0_2_x0 : std_logic;
signal \N_1331_0\ : std_logic;
signal currentchar_1_2 : std_logic;
signal currentchar_m7_0 : std_logic;
signal \un113_pixel_3_0_11__N_16_cascade_\ : std_logic;
signal \un113_pixel_7_1_7__N_11\ : std_logic;
signal \N_4573_0\ : std_logic;
signal un112_pixel_2_2 : std_logic;
signal currentchar_1_1 : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal currentchar_1_0 : std_logic;
signal un115_pixel_3_am_2 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_iZ0\ : std_logic;
signal \G_673\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal \G_674\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal column_1_i_3 : std_logic;
signal \ScreenBuffer_0_10_RNIGDGIE9Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0\ : std_logic;
signal \ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0\ : std_logic;
signal \ScreenBuffer_0_6_RNITJ4B17Z0Z_0\ : std_logic;
signal un6_rowlto1 : std_logic;
signal \ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0\ : std_logic;
signal \ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0\ : std_logic;
signal \ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0\ : std_logic;
signal \ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0\ : std_logic;
signal \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0\ : std_logic;
signal un6_rowlto0 : std_logic;
signal column_1_i_2 : std_logic;
signal \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_\ : std_logic;
signal \ScreenBuffer_0_7_RNIN5F98I1Z0Z_0\ : std_logic;
signal un115_pixel_5_am_sx_1 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \Clock12MHz_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \SDATA2_wire\ : std_logic;
signal \SCLK1_wire\ : std_logic;
signal \nCS2_wire\ : std_logic;
signal \SDATA1_wire\ : std_logic;
signal \nCS1_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \SCLK2_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \Clock12MHz_wire\ <= Clock12MHz;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    SDATA2 <= \SDATA2_wire\;
    SCLK1 <= \SCLK1_wire\;
    nCS2 <= \nCS2_wire\;
    \SDATA1_wire\ <= SDATA1;
    nCS1 <= \nCS1_wire\;
    Pixel <= \Pixel_wire\;
    SCLK2 <= \SCLK2_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__11489\,
            RESETB => \N__21892\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \Clock12MHz_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__26091\,
            GLOBALBUFFEROUTPUT => \Clock12MHz_c_g\
        );

    \Clock12MHz_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26093\,
            DIN => \N__26092\,
            DOUT => \N__26091\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26093\,
            PADOUT => \N__26092\,
            PADIN => \N__26091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26082\,
            DIN => \N__26081\,
            DOUT => \N__26080\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26082\,
            PADOUT => \N__26081\,
            PADIN => \N__26080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26073\,
            DIN => \N__26072\,
            DOUT => \N__26071\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26073\,
            PADOUT => \N__26072\,
            PADIN => \N__26071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDATA2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26064\,
            DIN => \N__26063\,
            DOUT => \N__26062\,
            PACKAGEPIN => \SDATA2_wire\
        );

    \SDATA2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26064\,
            PADOUT => \N__26063\,
            PADIN => \N__26062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26055\,
            DIN => \N__26054\,
            DOUT => \N__26053\,
            PACKAGEPIN => \SCLK1_wire\
        );

    \SCLK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26055\,
            PADOUT => \N__26054\,
            PADIN => \N__26053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13679\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26046\,
            DIN => \N__26045\,
            DOUT => \N__26044\,
            PACKAGEPIN => \nCS2_wire\
        );

    \nCS2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26046\,
            PADOUT => \N__26045\,
            PADIN => \N__26044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDATA1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26037\,
            DIN => \N__26036\,
            DOUT => \N__26035\,
            PACKAGEPIN => \SDATA1_wire\
        );

    \SDATA1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26037\,
            PADOUT => \N__26036\,
            PADIN => \N__26035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SDATA1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26028\,
            DIN => \N__26027\,
            DOUT => \N__26026\,
            PACKAGEPIN => \nCS1_wire\
        );

    \nCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26028\,
            PADOUT => \N__26027\,
            PADIN => \N__26026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26019\,
            DIN => \N__26018\,
            DOUT => \N__26017\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26019\,
            PADOUT => \N__26018\,
            PADIN => \N__26017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26010\,
            DIN => \N__26009\,
            DOUT => \N__26008\,
            PACKAGEPIN => \SCLK2_wire\
        );

    \SCLK2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26010\,
            PADOUT => \N__26009\,
            PADIN => \N__26008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13678\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6199\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25976\
        );

    \I__6198\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25976\
        );

    \I__6197\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25976\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__25988\,
            I => \N__25973\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__25987\,
            I => \N__25963\
        );

    \I__6194\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25953\
        );

    \I__6193\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25953\
        );

    \I__6192\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25950\
        );

    \I__6191\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25947\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__25976\,
            I => \N__25944\
        );

    \I__6189\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25941\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__25972\,
            I => \N__25938\
        );

    \I__6187\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25932\
        );

    \I__6186\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25932\
        );

    \I__6185\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25929\
        );

    \I__6184\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25926\
        );

    \I__6183\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25921\
        );

    \I__6182\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25921\
        );

    \I__6181\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25918\
        );

    \I__6180\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25907\
        );

    \I__6179\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25907\
        );

    \I__6178\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25907\
        );

    \I__6177\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25907\
        );

    \I__6176\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25907\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__25953\,
            I => \N__25902\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25902\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25899\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__25944\,
            I => \N__25896\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__25941\,
            I => \N__25893\
        );

    \I__6170\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25888\
        );

    \I__6169\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25888\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25885\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25882\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__25926\,
            I => \N__25875\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__25921\,
            I => \N__25875\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__25918\,
            I => \N__25875\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25872\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__25902\,
            I => \N__25862\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__25899\,
            I => \N__25862\
        );

    \I__6160\ : Span4Mux_v
    port map (
            O => \N__25896\,
            I => \N__25862\
        );

    \I__6159\ : Span4Mux_h
    port map (
            O => \N__25893\,
            I => \N__25855\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__25888\,
            I => \N__25855\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__25885\,
            I => \N__25855\
        );

    \I__6156\ : Span4Mux_s2_h
    port map (
            O => \N__25882\,
            I => \N__25852\
        );

    \I__6155\ : Span4Mux_s3_h
    port map (
            O => \N__25875\,
            I => \N__25847\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__25872\,
            I => \N__25847\
        );

    \I__6153\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25844\
        );

    \I__6152\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25841\
        );

    \I__6151\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25838\
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__25862\,
            I => column_1_i_3
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__25855\,
            I => column_1_i_3
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__25852\,
            I => column_1_i_3
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__25847\,
            I => column_1_i_3
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__25844\,
            I => column_1_i_3
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__25841\,
            I => column_1_i_3
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__25838\,
            I => column_1_i_3
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__6142\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25814\
        );

    \I__6141\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25814\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__25814\,
            I => \ScreenBuffer_0_10_RNIGDGIE9Z0Z_0\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__6138\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25802\
        );

    \I__6137\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25802\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__6135\ : Span4Mux_s0_h
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__25793\,
            I => \ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0\
        );

    \I__6132\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__6130\ : Odrv12
    port map (
            O => \N__25784\,
            I => \ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__25781\,
            I => \ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_\
        );

    \I__6128\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__25775\,
            I => \ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0\
        );

    \I__6126\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__6124\ : Span4Mux_s3_h
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__6123\ : Odrv4
    port map (
            O => \N__25763\,
            I => \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0\
        );

    \I__6122\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25756\
        );

    \I__6121\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25753\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__25756\,
            I => \N__25750\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__25750\,
            I => \ScreenBuffer_0_6_RNITJ4B17Z0Z_0\
        );

    \I__6117\ : Odrv4
    port map (
            O => \N__25747\,
            I => \ScreenBuffer_0_6_RNITJ4B17Z0Z_0\
        );

    \I__6116\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25729\
        );

    \I__6115\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25729\
        );

    \I__6114\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25726\
        );

    \I__6113\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25723\
        );

    \I__6112\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25720\
        );

    \I__6111\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25715\
        );

    \I__6110\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25715\
        );

    \I__6109\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25710\
        );

    \I__6108\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25710\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25705\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__25726\,
            I => \N__25694\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__25723\,
            I => \N__25694\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__25720\,
            I => \N__25694\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__25715\,
            I => \N__25694\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__25710\,
            I => \N__25694\
        );

    \I__6101\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25683\
        );

    \I__6100\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25680\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__25705\,
            I => \N__25677\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__25694\,
            I => \N__25674\
        );

    \I__6097\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25665\
        );

    \I__6096\ : InMux
    port map (
            O => \N__25692\,
            I => \N__25665\
        );

    \I__6095\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25665\
        );

    \I__6094\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25665\
        );

    \I__6093\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25662\
        );

    \I__6092\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25659\
        );

    \I__6091\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25654\
        );

    \I__6090\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25654\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__25683\,
            I => un6_rowlto1
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__25680\,
            I => un6_rowlto1
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__25677\,
            I => un6_rowlto1
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__25674\,
            I => un6_rowlto1
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__25665\,
            I => un6_rowlto1
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__25662\,
            I => un6_rowlto1
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__25659\,
            I => un6_rowlto1
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__25654\,
            I => un6_rowlto1
        );

    \I__6081\ : CascadeMux
    port map (
            O => \N__25637\,
            I => \N__25634\
        );

    \I__6080\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__6079\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25628\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__25628\,
            I => \ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0\
        );

    \I__6077\ : CascadeMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__6076\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25616\
        );

    \I__6075\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25616\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__6073\ : Span4Mux_s1_h
    port map (
            O => \N__25613\,
            I => \N__25610\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__25610\,
            I => \ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0\
        );

    \I__6071\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__25604\,
            I => \ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__25601\,
            I => \ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_\
        );

    \I__6068\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25595\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__25595\,
            I => \ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0\
        );

    \I__6066\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25587\
        );

    \I__6065\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25580\
        );

    \I__6064\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25580\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25577\
        );

    \I__6062\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25574\
        );

    \I__6061\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25571\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__25580\,
            I => \N__25568\
        );

    \I__6059\ : Span4Mux_v
    port map (
            O => \N__25577\,
            I => \N__25563\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__25574\,
            I => \N__25563\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__25571\,
            I => \N__25560\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__25568\,
            I => \N__25557\
        );

    \I__6055\ : Span4Mux_h
    port map (
            O => \N__25563\,
            I => \N__25554\
        );

    \I__6054\ : Odrv12
    port map (
            O => \N__25560\,
            I => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__25557\,
            I => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__25554\,
            I => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__25547\,
            I => \N__25542\
        );

    \I__6050\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25535\
        );

    \I__6049\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25532\
        );

    \I__6048\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25529\
        );

    \I__6047\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25526\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__25540\,
            I => \N__25522\
        );

    \I__6045\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25519\
        );

    \I__6044\ : CascadeMux
    port map (
            O => \N__25538\,
            I => \N__25514\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__25535\,
            I => \N__25509\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__25532\,
            I => \N__25506\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25501\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__25526\,
            I => \N__25501\
        );

    \I__6039\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25498\
        );

    \I__6038\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25495\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25492\
        );

    \I__6036\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25489\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__25517\,
            I => \N__25486\
        );

    \I__6034\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25483\
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__25513\,
            I => \N__25480\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__25512\,
            I => \N__25474\
        );

    \I__6031\ : Span4Mux_v
    port map (
            O => \N__25509\,
            I => \N__25463\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__25506\,
            I => \N__25463\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__25501\,
            I => \N__25463\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25463\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25463\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__25492\,
            I => \N__25458\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__25489\,
            I => \N__25458\
        );

    \I__6024\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25455\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__25483\,
            I => \N__25452\
        );

    \I__6022\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25443\
        );

    \I__6021\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25443\
        );

    \I__6020\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25443\
        );

    \I__6019\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25443\
        );

    \I__6018\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25440\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__25463\,
            I => \N__25437\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__25458\,
            I => \N__25432\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__25455\,
            I => \N__25432\
        );

    \I__6014\ : Span12Mux_s11_h
    port map (
            O => \N__25452\,
            I => \N__25427\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25427\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__25440\,
            I => un6_rowlto0
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__25437\,
            I => un6_rowlto0
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__25432\,
            I => un6_rowlto0
        );

    \I__6009\ : Odrv12
    port map (
            O => \N__25427\,
            I => un6_rowlto0
        );

    \I__6008\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25410\
        );

    \I__6007\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25410\
        );

    \I__6006\ : CascadeMux
    port map (
            O => \N__25416\,
            I => \N__25407\
        );

    \I__6005\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25391\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__25410\,
            I => \N__25388\
        );

    \I__6003\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25383\
        );

    \I__6002\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25380\
        );

    \I__6001\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25373\
        );

    \I__6000\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25373\
        );

    \I__5999\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25373\
        );

    \I__5998\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25370\
        );

    \I__5997\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25365\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25365\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__25399\,
            I => \N__25361\
        );

    \I__5994\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25357\
        );

    \I__5993\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25354\
        );

    \I__5992\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25351\
        );

    \I__5991\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25348\
        );

    \I__5990\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25345\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__25391\,
            I => \N__25340\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__25388\,
            I => \N__25340\
        );

    \I__5987\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25337\
        );

    \I__5986\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25334\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__25383\,
            I => \N__25327\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__25380\,
            I => \N__25327\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25327\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__25370\,
            I => \N__25322\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__25365\,
            I => \N__25322\
        );

    \I__5980\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25314\
        );

    \I__5979\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25314\
        );

    \I__5978\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25314\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25311\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25307\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25292\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__25348\,
            I => \N__25292\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25292\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__25340\,
            I => \N__25292\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__25337\,
            I => \N__25292\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__25334\,
            I => \N__25292\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__25327\,
            I => \N__25292\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__25322\,
            I => \N__25289\
        );

    \I__5967\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25286\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25280\
        );

    \I__5965\ : Span4Mux_h
    port map (
            O => \N__25311\,
            I => \N__25280\
        );

    \I__5964\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25277\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__25307\,
            I => \N__25268\
        );

    \I__5962\ : Span4Mux_v
    port map (
            O => \N__25292\,
            I => \N__25268\
        );

    \I__5961\ : Span4Mux_s0_h
    port map (
            O => \N__25289\,
            I => \N__25268\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25268\
        );

    \I__5959\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25265\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__25280\,
            I => column_1_i_2
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__25277\,
            I => column_1_i_2
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__25268\,
            I => column_1_i_2
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__25265\,
            I => column_1_i_2
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__25256\,
            I => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_\
        );

    \I__5953\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__5951\ : Span4Mux_s3_h
    port map (
            O => \N__25247\,
            I => \N__25243\
        );

    \I__5950\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25240\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__25243\,
            I => \ScreenBuffer_0_7_RNIN5F98I1Z0Z_0\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__25240\,
            I => \ScreenBuffer_0_7_RNIN5F98I1Z0Z_0\
        );

    \I__5947\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__25232\,
            I => un115_pixel_5_am_sx_1
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__25229\,
            I => \un113_pixel_3_0_11__N_16_cascade_\
        );

    \I__5944\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25221\
        );

    \I__5943\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25218\
        );

    \I__5942\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25215\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N__25208\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__25218\,
            I => \N__25202\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__25215\,
            I => \N__25199\
        );

    \I__5938\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25196\
        );

    \I__5937\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25191\
        );

    \I__5936\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25191\
        );

    \I__5935\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25188\
        );

    \I__5934\ : Span4Mux_s3_h
    port map (
            O => \N__25208\,
            I => \N__25185\
        );

    \I__5933\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25182\
        );

    \I__5932\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25177\
        );

    \I__5931\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25177\
        );

    \I__5930\ : Span4Mux_v
    port map (
            O => \N__25202\,
            I => \N__25168\
        );

    \I__5929\ : Span4Mux_s3_h
    port map (
            O => \N__25199\,
            I => \N__25168\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25168\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__25191\,
            I => \N__25168\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__25188\,
            I => \un113_pixel_7_1_7__N_11\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__25185\,
            I => \un113_pixel_7_1_7__N_11\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__25182\,
            I => \un113_pixel_7_1_7__N_11\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__25177\,
            I => \un113_pixel_7_1_7__N_11\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__25168\,
            I => \un113_pixel_7_1_7__N_11\
        );

    \I__5921\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__25154\,
            I => \N_4573_0\
        );

    \I__5919\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25146\
        );

    \I__5918\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25142\
        );

    \I__5917\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25137\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__25146\,
            I => \N__25130\
        );

    \I__5915\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25127\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__25142\,
            I => \N__25124\
        );

    \I__5913\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25119\
        );

    \I__5912\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25119\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25116\
        );

    \I__5910\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25113\
        );

    \I__5909\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25110\
        );

    \I__5908\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25105\
        );

    \I__5907\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25105\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__25130\,
            I => \N__25098\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__25127\,
            I => \N__25098\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__25124\,
            I => \N__25098\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__25119\,
            I => \N__25095\
        );

    \I__5902\ : Odrv12
    port map (
            O => \N__25116\,
            I => un112_pixel_2_2
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__25113\,
            I => un112_pixel_2_2
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__25110\,
            I => un112_pixel_2_2
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__25105\,
            I => un112_pixel_2_2
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__25098\,
            I => un112_pixel_2_2
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__25095\,
            I => un112_pixel_2_2
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__25082\,
            I => \N__25071\
        );

    \I__5895\ : InMux
    port map (
            O => \N__25081\,
            I => \N__25059\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25059\
        );

    \I__5893\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25053\
        );

    \I__5892\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25050\
        );

    \I__5891\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25043\
        );

    \I__5890\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25043\
        );

    \I__5889\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25043\
        );

    \I__5888\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25037\
        );

    \I__5887\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25037\
        );

    \I__5886\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25032\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__25069\,
            I => \N__25022\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__25068\,
            I => \N__25008\
        );

    \I__5883\ : InMux
    port map (
            O => \N__25067\,
            I => \N__24997\
        );

    \I__5882\ : InMux
    port map (
            O => \N__25066\,
            I => \N__24997\
        );

    \I__5881\ : InMux
    port map (
            O => \N__25065\,
            I => \N__24997\
        );

    \I__5880\ : InMux
    port map (
            O => \N__25064\,
            I => \N__24997\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__24992\
        );

    \I__5878\ : InMux
    port map (
            O => \N__25058\,
            I => \N__24985\
        );

    \I__5877\ : InMux
    port map (
            O => \N__25057\,
            I => \N__24985\
        );

    \I__5876\ : InMux
    port map (
            O => \N__25056\,
            I => \N__24985\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__24978\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__25050\,
            I => \N__24978\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__24978\
        );

    \I__5872\ : InMux
    port map (
            O => \N__25042\,
            I => \N__24975\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__25037\,
            I => \N__24972\
        );

    \I__5870\ : InMux
    port map (
            O => \N__25036\,
            I => \N__24967\
        );

    \I__5869\ : InMux
    port map (
            O => \N__25035\,
            I => \N__24967\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__25032\,
            I => \N__24964\
        );

    \I__5867\ : InMux
    port map (
            O => \N__25031\,
            I => \N__24959\
        );

    \I__5866\ : InMux
    port map (
            O => \N__25030\,
            I => \N__24959\
        );

    \I__5865\ : InMux
    port map (
            O => \N__25029\,
            I => \N__24954\
        );

    \I__5864\ : InMux
    port map (
            O => \N__25028\,
            I => \N__24954\
        );

    \I__5863\ : InMux
    port map (
            O => \N__25027\,
            I => \N__24949\
        );

    \I__5862\ : InMux
    port map (
            O => \N__25026\,
            I => \N__24949\
        );

    \I__5861\ : InMux
    port map (
            O => \N__25025\,
            I => \N__24938\
        );

    \I__5860\ : InMux
    port map (
            O => \N__25022\,
            I => \N__24938\
        );

    \I__5859\ : InMux
    port map (
            O => \N__25021\,
            I => \N__24938\
        );

    \I__5858\ : InMux
    port map (
            O => \N__25020\,
            I => \N__24938\
        );

    \I__5857\ : InMux
    port map (
            O => \N__25019\,
            I => \N__24938\
        );

    \I__5856\ : InMux
    port map (
            O => \N__25018\,
            I => \N__24929\
        );

    \I__5855\ : InMux
    port map (
            O => \N__25017\,
            I => \N__24929\
        );

    \I__5854\ : InMux
    port map (
            O => \N__25016\,
            I => \N__24929\
        );

    \I__5853\ : InMux
    port map (
            O => \N__25015\,
            I => \N__24929\
        );

    \I__5852\ : InMux
    port map (
            O => \N__25014\,
            I => \N__24920\
        );

    \I__5851\ : InMux
    port map (
            O => \N__25013\,
            I => \N__24920\
        );

    \I__5850\ : InMux
    port map (
            O => \N__25012\,
            I => \N__24920\
        );

    \I__5849\ : InMux
    port map (
            O => \N__25011\,
            I => \N__24920\
        );

    \I__5848\ : InMux
    port map (
            O => \N__25008\,
            I => \N__24915\
        );

    \I__5847\ : InMux
    port map (
            O => \N__25007\,
            I => \N__24915\
        );

    \I__5846\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24912\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__24997\,
            I => \N__24909\
        );

    \I__5844\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24904\
        );

    \I__5843\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24904\
        );

    \I__5842\ : Span4Mux_v
    port map (
            O => \N__24992\,
            I => \N__24897\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__24985\,
            I => \N__24897\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__24978\,
            I => \N__24897\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__24975\,
            I => \N__24890\
        );

    \I__5838\ : Span4Mux_s3_v
    port map (
            O => \N__24972\,
            I => \N__24890\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__24967\,
            I => \N__24890\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__24964\,
            I => currentchar_1_1
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__24959\,
            I => currentchar_1_1
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__24954\,
            I => currentchar_1_1
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__24949\,
            I => currentchar_1_1
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__24938\,
            I => currentchar_1_1
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__24929\,
            I => currentchar_1_1
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__24920\,
            I => currentchar_1_1
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__24915\,
            I => currentchar_1_1
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__24912\,
            I => currentchar_1_1
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__24909\,
            I => currentchar_1_1
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__24904\,
            I => currentchar_1_1
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__24897\,
            I => currentchar_1_1
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__24890\,
            I => currentchar_1_1
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__24863\,
            I => \N__24849\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__24862\,
            I => \N__24846\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__24861\,
            I => \N__24843\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__24860\,
            I => \N__24840\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__24859\,
            I => \N__24829\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__24858\,
            I => \N__24822\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__24857\,
            I => \N__24818\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__24856\,
            I => \N__24813\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__24855\,
            I => \N__24810\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__24854\,
            I => \N__24805\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__24853\,
            I => \N__24801\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__24852\,
            I => \N__24797\
        );

    \I__5811\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24794\
        );

    \I__5810\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24791\
        );

    \I__5809\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24786\
        );

    \I__5808\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24786\
        );

    \I__5807\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24781\
        );

    \I__5806\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24781\
        );

    \I__5805\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24778\
        );

    \I__5804\ : InMux
    port map (
            O => \N__24836\,
            I => \N__24773\
        );

    \I__5803\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24770\
        );

    \I__5802\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24767\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__24833\,
            I => \N__24764\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__24832\,
            I => \N__24761\
        );

    \I__5799\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24756\
        );

    \I__5798\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24753\
        );

    \I__5797\ : CascadeMux
    port map (
            O => \N__24827\,
            I => \N__24749\
        );

    \I__5796\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24743\
        );

    \I__5795\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24743\
        );

    \I__5794\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24734\
        );

    \I__5793\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24734\
        );

    \I__5792\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24734\
        );

    \I__5791\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24734\
        );

    \I__5790\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24729\
        );

    \I__5789\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24729\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24726\
        );

    \I__5787\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24718\
        );

    \I__5786\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24718\
        );

    \I__5785\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24718\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__24804\,
            I => \N__24715\
        );

    \I__5783\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24712\
        );

    \I__5782\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24707\
        );

    \I__5781\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24707\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__24794\,
            I => \N__24704\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__24791\,
            I => \N__24695\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24695\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__24781\,
            I => \N__24695\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__24778\,
            I => \N__24695\
        );

    \I__5775\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24690\
        );

    \I__5774\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24690\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24683\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24683\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24683\
        );

    \I__5770\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24678\
        );

    \I__5769\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24678\
        );

    \I__5768\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24673\
        );

    \I__5767\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24673\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24670\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__24753\,
            I => \N__24667\
        );

    \I__5764\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24664\
        );

    \I__5763\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24659\
        );

    \I__5762\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24659\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24656\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__24734\,
            I => \N__24649\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__24729\,
            I => \N__24649\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24649\
        );

    \I__5757\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24646\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__24718\,
            I => \N__24643\
        );

    \I__5755\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24640\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__24712\,
            I => \N__24636\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24629\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__24704\,
            I => \N__24629\
        );

    \I__5751\ : Span4Mux_s3_v
    port map (
            O => \N__24695\,
            I => \N__24629\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24622\
        );

    \I__5749\ : Span4Mux_v
    port map (
            O => \N__24683\,
            I => \N__24622\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24678\,
            I => \N__24622\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24619\
        );

    \I__5746\ : Span4Mux_v
    port map (
            O => \N__24670\,
            I => \N__24616\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__24667\,
            I => \N__24613\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__24664\,
            I => \N__24598\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__24659\,
            I => \N__24598\
        );

    \I__5742\ : Span4Mux_v
    port map (
            O => \N__24656\,
            I => \N__24598\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__24649\,
            I => \N__24598\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24598\
        );

    \I__5739\ : Span4Mux_s2_h
    port map (
            O => \N__24643\,
            I => \N__24598\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24598\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__24639\,
            I => \N__24595\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__24636\,
            I => \N__24588\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__24629\,
            I => \N__24588\
        );

    \I__5734\ : Span4Mux_h
    port map (
            O => \N__24622\,
            I => \N__24583\
        );

    \I__5733\ : Span4Mux_v
    port map (
            O => \N__24619\,
            I => \N__24583\
        );

    \I__5732\ : Span4Mux_s1_h
    port map (
            O => \N__24616\,
            I => \N__24580\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__24613\,
            I => \N__24575\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__24598\,
            I => \N__24575\
        );

    \I__5729\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24572\
        );

    \I__5728\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24567\
        );

    \I__5727\ : InMux
    port map (
            O => \N__24593\,
            I => \N__24567\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__24588\,
            I => \N__24564\
        );

    \I__5725\ : Span4Mux_v
    port map (
            O => \N__24583\,
            I => \N__24561\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__24580\,
            I => \N__24556\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__24575\,
            I => \N__24556\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__24572\,
            I => \beamYZ0Z_0\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__24567\,
            I => \beamYZ0Z_0\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__24564\,
            I => \beamYZ0Z_0\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__24561\,
            I => \beamYZ0Z_0\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__24556\,
            I => \beamYZ0Z_0\
        );

    \I__5717\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24537\
        );

    \I__5716\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24532\
        );

    \I__5715\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24529\
        );

    \I__5714\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24526\
        );

    \I__5713\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24521\
        );

    \I__5712\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24518\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__24537\,
            I => \N__24515\
        );

    \I__5710\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24499\
        );

    \I__5709\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24499\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__24532\,
            I => \N__24496\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__24529\,
            I => \N__24493\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__24526\,
            I => \N__24490\
        );

    \I__5705\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24485\
        );

    \I__5704\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24485\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24468\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24463\
        );

    \I__5701\ : Span4Mux_s3_h
    port map (
            O => \N__24515\,
            I => \N__24463\
        );

    \I__5700\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24458\
        );

    \I__5699\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24458\
        );

    \I__5698\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24451\
        );

    \I__5697\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24451\
        );

    \I__5696\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24451\
        );

    \I__5695\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24440\
        );

    \I__5694\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24440\
        );

    \I__5693\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24440\
        );

    \I__5692\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24440\
        );

    \I__5691\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24440\
        );

    \I__5690\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24437\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__24499\,
            I => \N__24432\
        );

    \I__5688\ : Span4Mux_s3_h
    port map (
            O => \N__24496\,
            I => \N__24432\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__24493\,
            I => \N__24425\
        );

    \I__5686\ : Span4Mux_v
    port map (
            O => \N__24490\,
            I => \N__24425\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__24485\,
            I => \N__24425\
        );

    \I__5684\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24420\
        );

    \I__5683\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24420\
        );

    \I__5682\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24413\
        );

    \I__5681\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24413\
        );

    \I__5680\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24413\
        );

    \I__5679\ : InMux
    port map (
            O => \N__24479\,
            I => \N__24404\
        );

    \I__5678\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24404\
        );

    \I__5677\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24404\
        );

    \I__5676\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24404\
        );

    \I__5675\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24393\
        );

    \I__5674\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24393\
        );

    \I__5673\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24393\
        );

    \I__5672\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24393\
        );

    \I__5671\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24393\
        );

    \I__5670\ : Odrv12
    port map (
            O => \N__24468\,
            I => currentchar_1_0
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__24463\,
            I => currentchar_1_0
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__24458\,
            I => currentchar_1_0
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__24451\,
            I => currentchar_1_0
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__24440\,
            I => currentchar_1_0
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__24437\,
            I => currentchar_1_0
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__24432\,
            I => currentchar_1_0
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__24425\,
            I => currentchar_1_0
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__24420\,
            I => currentchar_1_0
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__24413\,
            I => currentchar_1_0
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__24404\,
            I => currentchar_1_0
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__24393\,
            I => currentchar_1_0
        );

    \I__5658\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__24365\,
            I => un115_pixel_3_am_2
        );

    \I__5656\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24355\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__24358\,
            I => \N__24350\
        );

    \I__5653\ : Span4Mux_s0_h
    port map (
            O => \N__24355\,
            I => \N__24344\
        );

    \I__5652\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24333\
        );

    \I__5651\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24333\
        );

    \I__5650\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24333\
        );

    \I__5649\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24333\
        );

    \I__5648\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24333\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__24347\,
            I => \N__24330\
        );

    \I__5646\ : Span4Mux_h
    port map (
            O => \N__24344\,
            I => \N__24325\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24325\
        );

    \I__5644\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24322\
        );

    \I__5643\ : Sp12to4
    port map (
            O => \N__24325\,
            I => \N__24317\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__24322\,
            I => \N__24317\
        );

    \I__5641\ : Odrv12
    port map (
            O => \N__24317\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__5639\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24308\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__24308\,
            I => \column_1_if_generate_plus_mult1_un75_sum_iZ0\
        );

    \I__5637\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__24302\,
            I => \G_673\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__5634\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__24293\,
            I => if_generate_plus_mult1_un75_sum_cry_2_s
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__5631\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24284\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__24284\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__5629\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24278\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__24278\,
            I => \G_674\
        );

    \I__5627\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__24272\,
            I => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__5625\ : InMux
    port map (
            O => \N__24269\,
            I => column_1_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__5624\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__24263\,
            I => \N_1303_0\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__24260\,
            I => \g0_16_x0_cascade_\
        );

    \I__5621\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__24254\,
            I => g0_16_x1
        );

    \I__5619\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__24245\,
            I => \N_4560_0\
        );

    \I__5616\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__24239\,
            I => \N__24236\
        );

    \I__5614\ : Span4Mux_h
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__24233\,
            I => \N_1309_0\
        );

    \I__5612\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24226\
        );

    \I__5611\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24223\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__24226\,
            I => \N__24220\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__24223\,
            I => \N__24217\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__24220\,
            I => \un113_pixel_4_0_15__N_2\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__24217\,
            I => \un113_pixel_4_0_15__N_2\
        );

    \I__5606\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__5604\ : Span4Mux_s3_h
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__24203\,
            I => \un113_pixel_7_1_7__N_9\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__24200\,
            I => \beamY_RNIJIDRG11Z0Z_0_cascade_\
        );

    \I__5601\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__5599\ : Span4Mux_s2_h
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__24188\,
            I => \beamY_RNIJIDRG11_0Z0Z_0\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__24185\,
            I => \beamY_RNIRG0LHO1Z0Z_0_cascade_\
        );

    \I__5596\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24176\
        );

    \I__5595\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24176\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__24173\,
            I => \ScreenBuffer_0_7_RNIB3R6U63Z0Z_0\
        );

    \I__5592\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24163\
        );

    \I__5591\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24163\
        );

    \I__5590\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24155\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__24163\,
            I => \N__24150\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__24162\,
            I => \N__24147\
        );

    \I__5587\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24139\
        );

    \I__5586\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24139\
        );

    \I__5585\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24139\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__24158\,
            I => \N__24132\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__24155\,
            I => \N__24127\
        );

    \I__5582\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24124\
        );

    \I__5581\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24121\
        );

    \I__5580\ : Span4Mux_s2_v
    port map (
            O => \N__24150\,
            I => \N__24118\
        );

    \I__5579\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24114\
        );

    \I__5578\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24111\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24108\
        );

    \I__5576\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24105\
        );

    \I__5575\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24100\
        );

    \I__5574\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24100\
        );

    \I__5573\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24093\
        );

    \I__5572\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24093\
        );

    \I__5571\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24093\
        );

    \I__5570\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24090\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__24127\,
            I => \N__24081\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__24124\,
            I => \N__24081\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24081\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__24118\,
            I => \N__24081\
        );

    \I__5565\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24078\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__24114\,
            I => \N__24071\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__24111\,
            I => \N__24071\
        );

    \I__5562\ : Span4Mux_s3_v
    port map (
            O => \N__24108\,
            I => \N__24071\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24068\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__24100\,
            I => \N__24063\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__24093\,
            I => \N__24063\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__24090\,
            I => \N__24060\
        );

    \I__5557\ : Span4Mux_v
    port map (
            O => \N__24081\,
            I => \N__24057\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24052\
        );

    \I__5555\ : Span4Mux_v
    port map (
            O => \N__24071\,
            I => \N__24052\
        );

    \I__5554\ : Span4Mux_v
    port map (
            O => \N__24068\,
            I => \N__24049\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__24063\,
            I => \N__24046\
        );

    \I__5552\ : Odrv12
    port map (
            O => \N__24060\,
            I => font_un28_pixel_29
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__24057\,
            I => font_un28_pixel_29
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__24052\,
            I => font_un28_pixel_29
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__24049\,
            I => font_un28_pixel_29
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__24046\,
            I => font_un28_pixel_29
        );

    \I__5547\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24032\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__24032\,
            I => \beamY_RNIRG0LHO1Z0Z_0\
        );

    \I__5545\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__24023\
        );

    \I__5543\ : Odrv12
    port map (
            O => \N__24023\,
            I => \ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__24020\,
            I => \g0_2_x1_cascade_\
        );

    \I__5541\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__24014\,
            I => g0_2_x0
        );

    \I__5539\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24005\
        );

    \I__5538\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24005\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__24005\,
            I => \N_1331_0\
        );

    \I__5536\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23995\
        );

    \I__5535\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23991\
        );

    \I__5534\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23988\
        );

    \I__5533\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23982\
        );

    \I__5532\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23982\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__23995\,
            I => \N__23979\
        );

    \I__5530\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23976\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23973\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23963\
        );

    \I__5527\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23960\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23951\
        );

    \I__5525\ : Span4Mux_s2_v
    port map (
            O => \N__23979\,
            I => \N__23944\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__23976\,
            I => \N__23944\
        );

    \I__5523\ : Span4Mux_s3_h
    port map (
            O => \N__23973\,
            I => \N__23944\
        );

    \I__5522\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23941\
        );

    \I__5521\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23936\
        );

    \I__5520\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23936\
        );

    \I__5519\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23927\
        );

    \I__5518\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23927\
        );

    \I__5517\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23927\
        );

    \I__5516\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23927\
        );

    \I__5515\ : Span12Mux_s4_h
    port map (
            O => \N__23963\,
            I => \N__23922\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23922\
        );

    \I__5513\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23917\
        );

    \I__5512\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23917\
        );

    \I__5511\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23908\
        );

    \I__5510\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23908\
        );

    \I__5509\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23908\
        );

    \I__5508\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23908\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__23951\,
            I => currentchar_1_2
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__23944\,
            I => currentchar_1_2
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__23941\,
            I => currentchar_1_2
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__23936\,
            I => currentchar_1_2
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__23927\,
            I => currentchar_1_2
        );

    \I__5502\ : Odrv12
    port map (
            O => \N__23922\,
            I => currentchar_1_2
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__23917\,
            I => currentchar_1_2
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__23908\,
            I => currentchar_1_2
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__5498\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23874\
        );

    \I__5497\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23871\
        );

    \I__5496\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23867\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__23885\,
            I => \N__23861\
        );

    \I__5494\ : CascadeMux
    port map (
            O => \N__23884\,
            I => \N__23856\
        );

    \I__5493\ : CascadeMux
    port map (
            O => \N__23883\,
            I => \N__23853\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__23882\,
            I => \N__23849\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__23881\,
            I => \N__23846\
        );

    \I__5490\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23839\
        );

    \I__5489\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23839\
        );

    \I__5488\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23836\
        );

    \I__5487\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23833\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23830\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23827\
        );

    \I__5484\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23824\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__23867\,
            I => \N__23821\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__23866\,
            I => \N__23818\
        );

    \I__5481\ : CascadeMux
    port map (
            O => \N__23865\,
            I => \N__23815\
        );

    \I__5480\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23810\
        );

    \I__5479\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23810\
        );

    \I__5478\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23807\
        );

    \I__5477\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23802\
        );

    \I__5476\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23802\
        );

    \I__5475\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23799\
        );

    \I__5474\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23792\
        );

    \I__5473\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23792\
        );

    \I__5472\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23792\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__23845\,
            I => \N__23785\
        );

    \I__5470\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23782\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23779\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__23836\,
            I => \N__23774\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23774\
        );

    \I__5466\ : Span4Mux_s1_h
    port map (
            O => \N__23830\,
            I => \N__23765\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__23827\,
            I => \N__23765\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23765\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__23821\,
            I => \N__23765\
        );

    \I__5462\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23760\
        );

    \I__5461\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23760\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23753\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23753\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__23802\,
            I => \N__23753\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__23799\,
            I => \N__23748\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23748\
        );

    \I__5455\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23745\
        );

    \I__5454\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23736\
        );

    \I__5453\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23736\
        );

    \I__5452\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23736\
        );

    \I__5451\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23736\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__23782\,
            I => currentchar_m7_0
        );

    \I__5449\ : Odrv12
    port map (
            O => \N__23779\,
            I => currentchar_m7_0
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__23774\,
            I => currentchar_m7_0
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__23765\,
            I => currentchar_m7_0
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__23760\,
            I => currentchar_m7_0
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__23753\,
            I => currentchar_m7_0
        );

    \I__5444\ : Odrv12
    port map (
            O => \N__23748\,
            I => currentchar_m7_0
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__23745\,
            I => currentchar_m7_0
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__23736\,
            I => currentchar_m7_0
        );

    \I__5441\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__23708\,
            I => \N__23704\
        );

    \I__5437\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23701\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__23701\,
            I => \ScreenBuffer_0_10Z0Z_0\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__23698\,
            I => \ScreenBuffer_0_10Z0Z_0\
        );

    \I__5433\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__5431\ : Span4Mux_s1_h
    port map (
            O => \N__23687\,
            I => \N__23683\
        );

    \I__5430\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23680\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__23683\,
            I => \N__23677\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__23680\,
            I => \ScreenBuffer_0_11Z0Z_0\
        );

    \I__5427\ : Odrv4
    port map (
            O => \N__23677\,
            I => \ScreenBuffer_0_11Z0Z_0\
        );

    \I__5426\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__23663\,
            I => \ScreenBuffer_1_3Z0Z_0\
        );

    \I__5422\ : CascadeMux
    port map (
            O => \N__23660\,
            I => \currentchar_1_5_ns_1_0_cascade_\
        );

    \I__5421\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__23648\,
            I => \N__23644\
        );

    \I__5417\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23641\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__23644\,
            I => \N__23638\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__23641\,
            I => \ScreenBuffer_0_3Z0Z_0\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__23638\,
            I => \ScreenBuffer_0_3Z0Z_0\
        );

    \I__5413\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__5411\ : Span4Mux_s2_h
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__23624\,
            I => \beamY_RNIVDIFFI1Z0Z_0\
        );

    \I__5409\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__23618\,
            I => \beamY_RNI2RNL4M2Z0Z_0\
        );

    \I__5407\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23609\
        );

    \I__5406\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23600\
        );

    \I__5405\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23595\
        );

    \I__5404\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23595\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23592\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__23608\,
            I => \N__23589\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__23607\,
            I => \N__23586\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23582\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__23605\,
            I => \N__23579\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__23604\,
            I => \N__23576\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__23603\,
            I => \N__23573\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23568\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23568\
        );

    \I__5394\ : Span4Mux_h
    port map (
            O => \N__23592\,
            I => \N__23565\
        );

    \I__5393\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23560\
        );

    \I__5392\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23560\
        );

    \I__5391\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23555\
        );

    \I__5390\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23555\
        );

    \I__5389\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23548\
        );

    \I__5388\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23548\
        );

    \I__5387\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23548\
        );

    \I__5386\ : Span4Mux_v
    port map (
            O => \N__23568\,
            I => \N__23545\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__23565\,
            I => un3_rowlto1
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__23560\,
            I => un3_rowlto1
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__23555\,
            I => un3_rowlto1
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__23548\,
            I => un3_rowlto1
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__23545\,
            I => un3_rowlto1
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__5379\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23524\
        );

    \I__5378\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23519\
        );

    \I__5377\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23519\
        );

    \I__5376\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23514\
        );

    \I__5375\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23514\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__23524\,
            I => \N__23505\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__23519\,
            I => \N__23505\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23499\
        );

    \I__5371\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23496\
        );

    \I__5370\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23489\
        );

    \I__5369\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23489\
        );

    \I__5368\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23489\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__23505\,
            I => \N__23486\
        );

    \I__5366\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23479\
        );

    \I__5365\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23479\
        );

    \I__5364\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23479\
        );

    \I__5363\ : Span4Mux_v
    port map (
            O => \N__23499\,
            I => \N__23468\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23468\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23468\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__23486\,
            I => \N__23468\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23468\
        );

    \I__5358\ : Odrv4
    port map (
            O => \N__23468\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__23465\,
            I => \N__23461\
        );

    \I__5356\ : CascadeMux
    port map (
            O => \N__23464\,
            I => \N__23458\
        );

    \I__5355\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23453\
        );

    \I__5354\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23453\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__23450\,
            I => \N_52\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__5350\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23440\
        );

    \I__5349\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23436\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__23440\,
            I => \N__23430\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__23439\,
            I => \N__23426\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23418\
        );

    \I__5345\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23413\
        );

    \I__5344\ : InMux
    port map (
            O => \N__23434\,
            I => \N__23413\
        );

    \I__5343\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23410\
        );

    \I__5342\ : Span4Mux_s3_h
    port map (
            O => \N__23430\,
            I => \N__23407\
        );

    \I__5341\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23404\
        );

    \I__5340\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23399\
        );

    \I__5339\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23399\
        );

    \I__5338\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23390\
        );

    \I__5337\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23390\
        );

    \I__5336\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23390\
        );

    \I__5335\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23390\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__23418\,
            I => un112_pixel_2_8
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__23413\,
            I => un112_pixel_2_8
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__23410\,
            I => un112_pixel_2_8
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__23407\,
            I => un112_pixel_2_8
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__23404\,
            I => un112_pixel_2_8
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__23399\,
            I => un112_pixel_2_8
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__23390\,
            I => un112_pixel_2_8
        );

    \I__5327\ : CascadeMux
    port map (
            O => \N__23375\,
            I => \N_4581_0_cascade_\
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \N_1296_0_cascade_\
        );

    \I__5325\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N_1296_0\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__5322\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__5321\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23354\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23350\
        );

    \I__5319\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23340\
        );

    \I__5318\ : Span4Mux_v
    port map (
            O => \N__23350\,
            I => \N__23337\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N__23332\
        );

    \I__5316\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23329\
        );

    \I__5315\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23326\
        );

    \I__5314\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23323\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \N__23319\
        );

    \I__5312\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23314\
        );

    \I__5311\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23314\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__23340\,
            I => \N__23311\
        );

    \I__5309\ : IoSpan4Mux
    port map (
            O => \N__23337\,
            I => \N__23308\
        );

    \I__5308\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23303\
        );

    \I__5307\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23303\
        );

    \I__5306\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23297\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__23329\,
            I => \N__23294\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__23326\,
            I => \N__23289\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__23323\,
            I => \N__23289\
        );

    \I__5302\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23286\
        );

    \I__5301\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23281\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__23314\,
            I => \N__23272\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__23311\,
            I => \N__23272\
        );

    \I__5298\ : Span4Mux_s2_h
    port map (
            O => \N__23308\,
            I => \N__23272\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23272\
        );

    \I__5296\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23269\
        );

    \I__5295\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23266\
        );

    \I__5294\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23261\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__23297\,
            I => \N__23254\
        );

    \I__5292\ : Span4Mux_h
    port map (
            O => \N__23294\,
            I => \N__23254\
        );

    \I__5291\ : Span4Mux_s3_v
    port map (
            O => \N__23289\,
            I => \N__23254\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23251\
        );

    \I__5289\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23248\
        );

    \I__5288\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23245\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23236\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__23272\,
            I => \N__23236\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__23269\,
            I => \N__23236\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__23266\,
            I => \N__23233\
        );

    \I__5283\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23226\
        );

    \I__5282\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23226\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23217\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23217\
        );

    \I__5279\ : Span4Mux_v
    port map (
            O => \N__23251\,
            I => \N__23217\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__23248\,
            I => \N__23217\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23214\
        );

    \I__5276\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23209\
        );

    \I__5275\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23209\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__23236\,
            I => \N__23206\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__23233\,
            I => \N__23203\
        );

    \I__5272\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23200\
        );

    \I__5271\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23197\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23192\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__23217\,
            I => \N__23192\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__23214\,
            I => \N__23185\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__23209\,
            I => \N__23185\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__23206\,
            I => \N__23185\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__23203\,
            I => \beamYZ0Z_1\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__23200\,
            I => \beamYZ0Z_1\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__23197\,
            I => \beamYZ0Z_1\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__23192\,
            I => \beamYZ0Z_1\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__23185\,
            I => \beamYZ0Z_1\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__5259\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__23162\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__5255\ : InMux
    port map (
            O => \N__23159\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__5254\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__23153\,
            I => if_generate_plus_mult1_un75_sum_axb_4_l_fx
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__5251\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23143\
        );

    \I__5250\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23140\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23137\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__23140\,
            I => \N__23134\
        );

    \I__5247\ : Span4Mux_s3_h
    port map (
            O => \N__23137\,
            I => \N__23131\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__23134\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__23131\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__5244\ : InMux
    port map (
            O => \N__23126\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__5243\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__5241\ : Span4Mux_s3_h
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__23114\,
            I => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__5239\ : InMux
    port map (
            O => \N__23111\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__5238\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__23102\,
            I => \N__23099\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__23096\,
            I => un6_rowlt7_0
        );

    \I__5233\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23090\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__23090\,
            I => \N__23085\
        );

    \I__5231\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23082\
        );

    \I__5230\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23077\
        );

    \I__5229\ : Span4Mux_v
    port map (
            O => \N__23085\,
            I => \N__23074\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__23082\,
            I => \N__23071\
        );

    \I__5227\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23068\
        );

    \I__5226\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23065\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23062\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__23074\,
            I => \N__23059\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__23071\,
            I => \N__23054\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23054\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23051\
        );

    \I__5220\ : Odrv12
    port map (
            O => \N__23062\,
            I => chessboardpixel_un151_pixel_24
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__23059\,
            I => chessboardpixel_un151_pixel_24
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__23054\,
            I => chessboardpixel_un151_pixel_24
        );

    \I__5217\ : Odrv12
    port map (
            O => \N__23051\,
            I => chessboardpixel_un151_pixel_24
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__23036\,
            I => \column_1_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__23033\,
            I => \N__23027\
        );

    \I__5212\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23024\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__23031\,
            I => \N__23021\
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__23030\,
            I => \N__23012\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23009\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23024\,
            I => \N__23006\
        );

    \I__5207\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23003\
        );

    \I__5206\ : InMux
    port map (
            O => \N__23020\,
            I => \N__22998\
        );

    \I__5205\ : InMux
    port map (
            O => \N__23019\,
            I => \N__22998\
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__23018\,
            I => \N__22995\
        );

    \I__5203\ : InMux
    port map (
            O => \N__23017\,
            I => \N__22991\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__23016\,
            I => \N__22987\
        );

    \I__5201\ : InMux
    port map (
            O => \N__23015\,
            I => \N__22979\
        );

    \I__5200\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22979\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__22970\
        );

    \I__5198\ : Span4Mux_v
    port map (
            O => \N__23006\,
            I => \N__22970\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__23003\,
            I => \N__22970\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__22998\,
            I => \N__22970\
        );

    \I__5195\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22965\
        );

    \I__5194\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22965\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22962\
        );

    \I__5192\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22957\
        );

    \I__5191\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22957\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__22986\,
            I => \N__22954\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__22985\,
            I => \N__22951\
        );

    \I__5188\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22948\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22945\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__22970\,
            I => \N__22940\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22940\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__22962\,
            I => \N__22935\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22935\
        );

    \I__5182\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22930\
        );

    \I__5181\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22930\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__22948\,
            I => un3_rowlto0
        );

    \I__5179\ : Odrv12
    port map (
            O => \N__22945\,
            I => un3_rowlto0
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__22940\,
            I => un3_rowlto0
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__22935\,
            I => un3_rowlto0
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__22930\,
            I => un3_rowlto0
        );

    \I__5175\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__22910\,
            I => \un113_pixel_3_0_11__currentchar_m7_0Z0Z_1\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__22907\,
            I => \d_N_3_mux_cascade_\
        );

    \I__5170\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22898\
        );

    \I__5168\ : Span4Mux_v
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__22892\,
            I => \ScreenBuffer_1_2Z0Z_2\
        );

    \I__5165\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22886\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__5163\ : Span4Mux_s2_h
    port map (
            O => \N__22883\,
            I => \N__22880\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__22880\,
            I => \N__22877\
        );

    \I__5161\ : Odrv4
    port map (
            O => \N__22877\,
            I => \ScreenBuffer_1_1Z0Z_2\
        );

    \I__5160\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__22865\,
            I => \un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__5155\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__5153\ : Odrv12
    port map (
            O => \N__22853\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__5151\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22844\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22844\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\
        );

    \I__5149\ : InMux
    port map (
            O => \N__22841\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__5148\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__22835\,
            I => charx_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__5146\ : InMux
    port map (
            O => \N__22832\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__5145\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__22823\,
            I => charx_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__5142\ : InMux
    port map (
            O => \N__22820\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__5141\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__22814\,
            I => \N__22809\
        );

    \I__5139\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22806\
        );

    \I__5138\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22803\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__22809\,
            I => \N__22800\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__22806\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__22803\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__22800\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__22793\,
            I => \N__22789\
        );

    \I__5132\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22784\
        );

    \I__5131\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22784\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__5129\ : Odrv12
    port map (
            O => \N__22781\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\
        );

    \I__5128\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22773\
        );

    \I__5127\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22770\
        );

    \I__5126\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22766\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22761\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__22770\,
            I => \N__22761\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22758\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__22766\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__5121\ : Odrv12
    port map (
            O => \N__22761\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__22758\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__5119\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__22748\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__22745\,
            I => \N__22740\
        );

    \I__5116\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22737\
        );

    \I__5115\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22733\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22727\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22724\
        );

    \I__5112\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22721\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22717\
        );

    \I__5110\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22712\
        );

    \I__5109\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22712\
        );

    \I__5108\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22709\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22704\
        );

    \I__5106\ : Span4Mux_v
    port map (
            O => \N__22724\,
            I => \N__22704\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__22721\,
            I => \N__22701\
        );

    \I__5104\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22698\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__22717\,
            I => \N__22695\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__22712\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__22709\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__22704\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5099\ : Odrv12
    port map (
            O => \N__22701\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__22698\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__22695\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__5095\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__22676\,
            I => charx_if_generate_plus_mult1_un40_sum_i
        );

    \I__5093\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22669\
        );

    \I__5092\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22666\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__22669\,
            I => \N__22659\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22659\
        );

    \I__5089\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22656\
        );

    \I__5088\ : InMux
    port map (
            O => \N__22664\,
            I => \N__22653\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__22659\,
            I => \N__22650\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22645\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22645\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__22650\,
            I => \N__22642\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__22645\,
            I => \N__22639\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__22642\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__22639\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__5080\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__5078\ : Odrv12
    port map (
            O => \N__22628\,
            I => column_1_i_i_2
        );

    \I__5077\ : InMux
    port map (
            O => \N__22625\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__22622\,
            I => \N__22615\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__22621\,
            I => \N__22612\
        );

    \I__5074\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22608\
        );

    \I__5073\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22604\
        );

    \I__5072\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22601\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22598\
        );

    \I__5070\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22593\
        );

    \I__5069\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22593\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__22608\,
            I => \N__22590\
        );

    \I__5067\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22587\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__22604\,
            I => \N__22582\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22582\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22577\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__22593\,
            I => \N__22577\
        );

    \I__5062\ : Span4Mux_s3_h
    port map (
            O => \N__22590\,
            I => \N__22574\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22569\
        );

    \I__5060\ : Span4Mux_v
    port map (
            O => \N__22582\,
            I => \N__22569\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__22577\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__22574\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__22569\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__5055\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__22550\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\
        );

    \I__5051\ : InMux
    port map (
            O => \N__22547\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__5049\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__22532\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\
        );

    \I__5045\ : InMux
    port map (
            O => \N__22529\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__5044\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22520\
        );

    \I__5043\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22520\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22517\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__22517\,
            I => charx_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__5040\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__22505\,
            I => charx_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__5036\ : InMux
    port map (
            O => \N__22502\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__5035\ : InMux
    port map (
            O => \N__22499\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__5034\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22488\
        );

    \I__5032\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22485\
        );

    \I__5031\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22482\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__22488\,
            I => \N__22477\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__22485\,
            I => \N__22477\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__22482\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__22477\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__5025\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__22466\,
            I => charx_if_generate_plus_mult1_un47_sum_i
        );

    \I__5023\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22456\
        );

    \I__5022\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22453\
        );

    \I__5021\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22450\
        );

    \I__5020\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22446\
        );

    \I__5019\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22443\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22440\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__22453\,
            I => \N__22437\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__22450\,
            I => \N__22434\
        );

    \I__5015\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22431\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__22446\,
            I => \N__22428\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__22443\,
            I => \N__22425\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__22440\,
            I => \N__22422\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__22437\,
            I => \N__22413\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__22434\,
            I => \N__22413\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22413\
        );

    \I__5008\ : Span4Mux_s3_h
    port map (
            O => \N__22428\,
            I => \N__22413\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__22425\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__22422\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__22413\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__5004\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__22400\,
            I => charx_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__5000\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__22391\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\
        );

    \I__4998\ : InMux
    port map (
            O => \N__22388\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__4997\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__4995\ : Odrv12
    port map (
            O => \N__22379\,
            I => column_1_if_generate_plus_mult1_un47_sum1_2
        );

    \I__4994\ : InMux
    port map (
            O => \N__22376\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_1
        );

    \I__4993\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__22364\,
            I => column_1_if_generate_plus_mult1_un47_sum1_3
        );

    \I__4989\ : InMux
    port map (
            O => \N__22361\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_2
        );

    \I__4988\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__22352\,
            I => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__4984\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__22337\,
            I => column_1_if_generate_plus_mult1_un47_sum1_4
        );

    \I__4980\ : InMux
    port map (
            O => \N__22334\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_3
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22327\
        );

    \I__4978\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22324\
        );

    \I__4977\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22321\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22314\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22314\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22311\
        );

    \I__4973\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22306\
        );

    \I__4972\ : Span4Mux_s3_v
    port map (
            O => \N__22314\,
            I => \N__22302\
        );

    \I__4971\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22299\
        );

    \I__4970\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22296\
        );

    \I__4969\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22293\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__22306\,
            I => \N__22290\
        );

    \I__4967\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22287\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__22302\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__22299\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__22296\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__22293\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__22290\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__22287\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__4960\ : InMux
    port map (
            O => \N__22274\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_4
        );

    \I__4959\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22265\
        );

    \I__4958\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22265\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__22262\,
            I => column_1_if_generate_plus_mult1_un47_sum1_5
        );

    \I__4955\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22246\
        );

    \I__4954\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22246\
        );

    \I__4953\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22243\
        );

    \I__4952\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22238\
        );

    \I__4951\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22238\
        );

    \I__4950\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22235\
        );

    \I__4949\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22232\
        );

    \I__4948\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22229\
        );

    \I__4947\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22226\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22223\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__22243\,
            I => \N__22220\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__22238\,
            I => \N__22217\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__22235\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__22232\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__22229\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__22226\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4939\ : Odrv12
    port map (
            O => \N__22223\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__22220\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4937\ : Odrv4
    port map (
            O => \N__22217\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__4936\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__22196\,
            I => un5_visiblex_i_0_25
        );

    \I__4933\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22189\
        );

    \I__4932\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22185\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22182\
        );

    \I__4930\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22179\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__22185\,
            I => \N__22176\
        );

    \I__4928\ : Span4Mux_s3_h
    port map (
            O => \N__22182\,
            I => \N__22171\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__22179\,
            I => \N__22171\
        );

    \I__4926\ : Span4Mux_s2_h
    port map (
            O => \N__22176\,
            I => \N__22168\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__22171\,
            I => \N_56\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__22168\,
            I => \N_56\
        );

    \I__4923\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22159\
        );

    \I__4922\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22154\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__22151\
        );

    \I__4920\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22148\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__22157\,
            I => \N__22144\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__22154\,
            I => \N__22137\
        );

    \I__4917\ : Span4Mux_s2_v
    port map (
            O => \N__22151\,
            I => \N__22132\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__22148\,
            I => \N__22132\
        );

    \I__4915\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22127\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22127\
        );

    \I__4913\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22120\
        );

    \I__4912\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22120\
        );

    \I__4911\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22120\
        );

    \I__4910\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22117\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__22137\,
            I => \N__22112\
        );

    \I__4908\ : Span4Mux_h
    port map (
            O => \N__22132\,
            I => \N__22112\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__22127\,
            I => \N__22107\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22107\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__22117\,
            I => \N_32_i\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__22112\,
            I => \N_32_i\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__22107\,
            I => \N_32_i\
        );

    \I__4902\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__22097\,
            I => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__22094\,
            I => \N__22089\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__22093\,
            I => \N__22081\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22078\
        );

    \I__4897\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22068\
        );

    \I__4896\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22060\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22060\
        );

    \I__4894\ : InMux
    port map (
            O => \N__22086\,
            I => \N__22060\
        );

    \I__4893\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22057\
        );

    \I__4892\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22048\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22048\
        );

    \I__4890\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22048\
        );

    \I__4889\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22048\
        );

    \I__4888\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22045\
        );

    \I__4887\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22036\
        );

    \I__4886\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22036\
        );

    \I__4885\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22036\
        );

    \I__4884\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22036\
        );

    \I__4883\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22033\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__22068\,
            I => \N__22029\
        );

    \I__4881\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22026\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__22060\,
            I => \N__22013\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22013\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__22048\,
            I => \N__22013\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__22045\,
            I => \N__22006\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22006\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__22033\,
            I => \N__22006\
        );

    \I__4874\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22000\
        );

    \I__4873\ : Span4Mux_s0_v
    port map (
            O => \N__22029\,
            I => \N__21995\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__21995\
        );

    \I__4871\ : InMux
    port map (
            O => \N__22025\,
            I => \N__21984\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22024\,
            I => \N__21984\
        );

    \I__4869\ : InMux
    port map (
            O => \N__22023\,
            I => \N__21984\
        );

    \I__4868\ : InMux
    port map (
            O => \N__22022\,
            I => \N__21984\
        );

    \I__4867\ : InMux
    port map (
            O => \N__22021\,
            I => \N__21984\
        );

    \I__4866\ : InMux
    port map (
            O => \N__22020\,
            I => \N__21981\
        );

    \I__4865\ : Span4Mux_s3_v
    port map (
            O => \N__22013\,
            I => \N__21978\
        );

    \I__4864\ : Span4Mux_h
    port map (
            O => \N__22006\,
            I => \N__21975\
        );

    \I__4863\ : InMux
    port map (
            O => \N__22005\,
            I => \N__21968\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22004\,
            I => \N__21968\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21968\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__22000\,
            I => \CO3_0\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__21995\,
            I => \CO3_0\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__21984\,
            I => \CO3_0\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__21981\,
            I => \CO3_0\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__21978\,
            I => \CO3_0\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__21975\,
            I => \CO3_0\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__21968\,
            I => \CO3_0\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__4852\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__21947\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3_i
        );

    \I__4850\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21940\
        );

    \I__4849\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21937\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__21940\,
            I => \un113_pixel_1_0_3__N_10_mux\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__21937\,
            I => \un113_pixel_1_0_3__N_10_mux\
        );

    \I__4846\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__21929\,
            I => \beamY_RNIMR86ES2Z0Z_0\
        );

    \I__4844\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__21920\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254\
        );

    \I__4841\ : InMux
    port map (
            O => \N__21917\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__21914\,
            I => \N__21909\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__21913\,
            I => \N__21905\
        );

    \I__4838\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21901\
        );

    \I__4837\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21893\
        );

    \I__4836\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21893\
        );

    \I__4835\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21893\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__21904\,
            I => \N__21889\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21884\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__21900\,
            I => \N__21881\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__21893\,
            I => \N__21878\
        );

    \I__4830\ : IoInMux
    port map (
            O => \N__21892\,
            I => \N__21875\
        );

    \I__4829\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21872\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__21888\,
            I => \N__21867\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__21887\,
            I => \N__21863\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__21884\,
            I => \N__21860\
        );

    \I__4825\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21857\
        );

    \I__4824\ : IoSpan4Mux
    port map (
            O => \N__21878\,
            I => \N__21852\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21852\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21848\
        );

    \I__4821\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21845\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__21870\,
            I => \N__21841\
        );

    \I__4819\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21838\
        );

    \I__4818\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21833\
        );

    \I__4817\ : InMux
    port map (
            O => \N__21863\,
            I => \N__21833\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__21860\,
            I => \N__21828\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21828\
        );

    \I__4814\ : IoSpan4Mux
    port map (
            O => \N__21852\,
            I => \N__21825\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__21851\,
            I => \N__21822\
        );

    \I__4812\ : Span4Mux_s2_v
    port map (
            O => \N__21848\,
            I => \N__21819\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21816\
        );

    \I__4810\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21811\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21811\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__21838\,
            I => \N__21808\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21805\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__21828\,
            I => \N__21802\
        );

    \I__4805\ : Span4Mux_s1_v
    port map (
            O => \N__21825\,
            I => \N__21799\
        );

    \I__4804\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21796\
        );

    \I__4803\ : Sp12to4
    port map (
            O => \N__21819\,
            I => \N__21789\
        );

    \I__4802\ : Span12Mux_v
    port map (
            O => \N__21816\,
            I => \N__21789\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21789\
        );

    \I__4800\ : Odrv12
    port map (
            O => \N__21808\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4799\ : Odrv12
    port map (
            O => \N__21805\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__21802\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__21799\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__21796\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4795\ : Odrv12
    port map (
            O => \N__21789\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__4793\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__21767\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464\
        );

    \I__4790\ : InMux
    port map (
            O => \N__21764\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__4789\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__21755\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21752\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__4785\ : InMux
    port map (
            O => \N__21749\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21737\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21737\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__21734\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__21728\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf
        );

    \I__4777\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__21722\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\
        );

    \I__4775\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__21716\,
            I => m17
        );

    \I__4773\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21710\,
            I => m12
        );

    \I__4771\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__21704\,
            I => un115_pixel_5_ns_x1_0
        );

    \I__4769\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__21698\,
            I => un115_pixel_5_ns_x0_0
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__21695\,
            I => \N_1325_cascade_\
        );

    \I__4766\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__21683\,
            I => un115_pixel_7_bm_0
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__21680\,
            I => \N_1315_cascade_\
        );

    \I__4761\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__21674\,
            I => \N_1322\
        );

    \I__4759\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N_1329\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__21665\,
            I => \N_1294_cascade_\
        );

    \I__4756\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__21659\,
            I => \beamY_RNICJUESD2_1Z0Z_0\
        );

    \I__4754\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N_1308\
        );

    \I__4752\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__21647\,
            I => un115_pixel_5_d_2
        );

    \I__4750\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N_1286_0_0_0\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21635\,
            I => \N_1289\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__21626\,
            I => \N__21620\
        );

    \I__4743\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21615\
        );

    \I__4742\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21615\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21612\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__21620\,
            I => font_un3_pixel_29
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__21615\,
            I => font_un3_pixel_29
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__21612\,
            I => font_un3_pixel_29
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__21605\,
            I => \N_4562_0_0_0_cascade_\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21596\
        );

    \I__4734\ : Odrv12
    port map (
            O => \N__21596\,
            I => \N_1340_0\
        );

    \I__4733\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__21590\,
            I => \beamY_RNICJUESD2_0Z0Z_0\
        );

    \I__4731\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__21578\,
            I => \beamY_RNI1H36941Z0Z_0\
        );

    \I__4727\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__21572\,
            I => font_un125_pixel_1_bm
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__21569\,
            I => \un113_pixel_6_1_5__N_11_cascade_\
        );

    \I__4724\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__21563\,
            I => \un113_pixel_2_0_3__N_8\
        );

    \I__4722\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__21557\,
            I => \beamY_RNICJUESD2_2Z0Z_0\
        );

    \I__4720\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21551\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__21551\,
            I => un115_pixel_5_s_7
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__21548\,
            I => \un115_pixel_5_am_7_cascade_\
        );

    \I__4717\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__21542\,
            I => un115_pixel_5_bm_7
        );

    \I__4715\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N_1288\
        );

    \I__4713\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__21530\,
            I => \N__21520\
        );

    \I__4711\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21517\
        );

    \I__4710\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21510\
        );

    \I__4709\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21510\
        );

    \I__4708\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21510\
        );

    \I__4707\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21503\
        );

    \I__4706\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21503\
        );

    \I__4705\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21503\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__21520\,
            I => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__21517\,
            I => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__21510\,
            I => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__21503\,
            I => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\
        );

    \I__4700\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4698\ : Span4Mux_s3_h
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__21485\,
            I => \un113_pixel_4_0_15__g1Z0Z_0\
        );

    \I__4696\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__4694\ : Span4Mux_s3_h
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__21473\,
            I => m9
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \m9_cascade_\
        );

    \I__4691\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__21464\,
            I => m6
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__21461\,
            I => \m6_cascade_\
        );

    \I__4688\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__4686\ : Odrv12
    port map (
            O => \N__21452\,
            I => \beamY_RNICJUESD2Z0Z_0\
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \un115_pixel_2_s_6_cascade_\
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__21446\,
            I => \un115_pixel_2_d_0_6_cascade_\
        );

    \I__4683\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__21440\,
            I => un115_pixel_3_bm_6
        );

    \I__4681\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21433\
        );

    \I__4680\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21430\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21425\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21425\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__21425\,
            I => \ScreenBuffer_1_2Z0Z_1\
        );

    \I__4676\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21418\
        );

    \I__4675\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21415\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__21418\,
            I => \ScreenBuffer_1_0Z0Z_1\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__21415\,
            I => \ScreenBuffer_1_0Z0Z_1\
        );

    \I__4672\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N_1_7_0\
        );

    \I__4670\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21400\
        );

    \I__4669\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21397\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21392\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21392\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__21389\,
            I => \ScreenBuffer_1_3Z0Z_1\
        );

    \I__4664\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21382\
        );

    \I__4663\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21379\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21374\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21374\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__21368\,
            I => \ScreenBuffer_1_1Z0Z_1\
        );

    \I__4657\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__21362\,
            I => m8
        );

    \I__4655\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21352\
        );

    \I__4653\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__21352\,
            I => \N__21346\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__21349\,
            I => \ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__21346\,
            I => \ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1\
        );

    \I__4649\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21337\
        );

    \I__4648\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21334\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21331\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__21334\,
            I => \ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__21331\,
            I => \ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1\
        );

    \I__4644\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21317\
        );

    \I__4643\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21317\
        );

    \I__4642\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21317\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__21317\,
            I => \N__21313\
        );

    \I__4640\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21310\
        );

    \I__4639\ : Odrv4
    port map (
            O => \N__21313\,
            I => \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__21310\,
            I => \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__21305\,
            I => \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_\
        );

    \I__4636\ : InMux
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__21299\,
            I => \un113_pixel_3_0_11__gZ0Z1\
        );

    \I__4634\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N__21290\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__21290\,
            I => \N__21286\
        );

    \I__4631\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__21286\,
            I => font_un3_pixel_28
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__21283\,
            I => font_un3_pixel_28
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__4627\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__21272\,
            I => \N_1342\
        );

    \I__4625\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__4623\ : Odrv12
    port map (
            O => \N__21263\,
            I => \un113_pixel_4_0_15__g0_5Z0Z_1\
        );

    \I__4622\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21255\
        );

    \I__4621\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21250\
        );

    \I__4620\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21250\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__21255\,
            I => font_un71_pixellt7_0_1
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__21250\,
            I => font_un71_pixellt7_0_1
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__4616\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__21239\,
            I => font_un64_pixel_ac0_5_0
        );

    \I__4614\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21232\
        );

    \I__4613\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21229\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__21229\,
            I => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__21226\,
            I => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3\
        );

    \I__4609\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__21212\,
            I => font_un3_pixel_0_29
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \un113_pixel_4_0_15__g0_5Z0Z_4_cascade_\
        );

    \I__4604\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N_9\
        );

    \I__4602\ : CascadeMux
    port map (
            O => \N__21200\,
            I => \un113_pixel_4_0_15__g2Z0Z_0_cascade_\
        );

    \I__4601\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__21188\,
            I => \N_4566_0\
        );

    \I__4597\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__21182\,
            I => un115_pixel_4
        );

    \I__4595\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__21176\,
            I => \N_4564_0\
        );

    \I__4593\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N_5_0\
        );

    \I__4591\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21160\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__21163\,
            I => \N__21154\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__21160\,
            I => \N__21151\
        );

    \I__4587\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21148\
        );

    \I__4586\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21141\
        );

    \I__4585\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21141\
        );

    \I__4584\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21141\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__21151\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__21148\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__21141\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1\
        );

    \I__4580\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__4578\ : Span4Mux_s3_h
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__21125\,
            I => \N_4561_0\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__4575\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__4572\ : Span4Mux_s3_h
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__21107\,
            I => g1_0
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__4569\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__21098\,
            I => \N_2075\
        );

    \I__4567\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__21086\,
            I => \N_11\
        );

    \I__4563\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__21080\,
            I => \un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0\
        );

    \I__4561\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__21074\,
            I => \un113_pixel_4_0_15__g0_i_a3_2\
        );

    \I__4559\ : IoInMux
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__4557\ : Odrv12
    port map (
            O => \N__21065\,
            I => \Pixel_c\
        );

    \I__4556\ : ClkMux
    port map (
            O => \N__21062\,
            I => \N__21029\
        );

    \I__4555\ : ClkMux
    port map (
            O => \N__21061\,
            I => \N__21029\
        );

    \I__4554\ : ClkMux
    port map (
            O => \N__21060\,
            I => \N__21029\
        );

    \I__4553\ : ClkMux
    port map (
            O => \N__21059\,
            I => \N__21029\
        );

    \I__4552\ : ClkMux
    port map (
            O => \N__21058\,
            I => \N__21029\
        );

    \I__4551\ : ClkMux
    port map (
            O => \N__21057\,
            I => \N__21029\
        );

    \I__4550\ : ClkMux
    port map (
            O => \N__21056\,
            I => \N__21029\
        );

    \I__4549\ : ClkMux
    port map (
            O => \N__21055\,
            I => \N__21029\
        );

    \I__4548\ : ClkMux
    port map (
            O => \N__21054\,
            I => \N__21029\
        );

    \I__4547\ : ClkMux
    port map (
            O => \N__21053\,
            I => \N__21029\
        );

    \I__4546\ : ClkMux
    port map (
            O => \N__21052\,
            I => \N__21029\
        );

    \I__4545\ : GlobalMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__4544\ : gio2CtrlBuf
    port map (
            O => \N__21026\,
            I => \PixelClock_g\
        );

    \I__4543\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__21017\,
            I => \un113_pixel_7_1_7__g0_6Z0Z_0\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__4539\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__4537\ : Sp12to4
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__4536\ : Odrv12
    port map (
            O => \N__21002\,
            I => \N_3078_0\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__20999\,
            I => \N_1297_0_cascade_\
        );

    \I__4534\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__20987\,
            I => font_un67_pixel_ac0_5_0
        );

    \I__4530\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20978\
        );

    \I__4529\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20975\
        );

    \I__4528\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20970\
        );

    \I__4527\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20970\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20967\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20963\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__20970\,
            I => \N__20960\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__20967\,
            I => \N__20957\
        );

    \I__4522\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20954\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__20963\,
            I => \N__20951\
        );

    \I__4520\ : Span4Mux_h
    port map (
            O => \N__20960\,
            I => \N__20948\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__20957\,
            I => chary_if_generate_plus_mult1_un68_sum_c5
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20954\,
            I => chary_if_generate_plus_mult1_un68_sum_c5
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__20951\,
            I => chary_if_generate_plus_mult1_un68_sum_c5
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__20948\,
            I => chary_if_generate_plus_mult1_un68_sum_c5
        );

    \I__4515\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20930\
        );

    \I__4513\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20925\
        );

    \I__4512\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20925\
        );

    \I__4511\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20921\
        );

    \I__4510\ : Span4Mux_s3_h
    port map (
            O => \N__20930\,
            I => \N__20916\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20916\
        );

    \I__4508\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20913\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__20921\,
            I => \N__20910\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__20916\,
            I => \N__20907\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__20913\,
            I => chary_if_generate_plus_mult1_un1_sum_axbxc3_2
        );

    \I__4504\ : Odrv12
    port map (
            O => \N__20910\,
            I => chary_if_generate_plus_mult1_un1_sum_axbxc3_2
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__20907\,
            I => chary_if_generate_plus_mult1_un1_sum_axbxc3_2
        );

    \I__4502\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__20897\,
            I => \un113_pixel_4_0_15__g0_4_0Z0Z_0\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__20894\,
            I => \N__20889\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__20893\,
            I => \N__20879\
        );

    \I__4498\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20876\
        );

    \I__4497\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20873\
        );

    \I__4496\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20866\
        );

    \I__4495\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20866\
        );

    \I__4494\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20866\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__20885\,
            I => \N__20862\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__20884\,
            I => \N__20859\
        );

    \I__4491\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20855\
        );

    \I__4490\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20850\
        );

    \I__4489\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20850\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20847\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20842\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20842\
        );

    \I__4485\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20833\
        );

    \I__4484\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20833\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20833\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__20858\,
            I => \N__20828\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__20855\,
            I => \N__20822\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20819\
        );

    \I__4479\ : Span4Mux_v
    port map (
            O => \N__20847\,
            I => \N__20816\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__20842\,
            I => \N__20813\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20810\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20807\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20804\
        );

    \I__4474\ : InMux
    port map (
            O => \N__20832\,
            I => \N__20801\
        );

    \I__4473\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20798\
        );

    \I__4472\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20791\
        );

    \I__4471\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20791\
        );

    \I__4470\ : InMux
    port map (
            O => \N__20826\,
            I => \N__20791\
        );

    \I__4469\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20786\
        );

    \I__4468\ : Span4Mux_v
    port map (
            O => \N__20822\,
            I => \N__20783\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__20819\,
            I => \N__20780\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__20816\,
            I => \N__20773\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__20813\,
            I => \N__20773\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__20810\,
            I => \N__20773\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20770\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__20804\,
            I => \N__20767\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__20801\,
            I => \N__20764\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__20798\,
            I => \N__20759\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__20791\,
            I => \N__20759\
        );

    \I__4458\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20756\
        );

    \I__4457\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20748\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20745\
        );

    \I__4455\ : Span4Mux_h
    port map (
            O => \N__20783\,
            I => \N__20742\
        );

    \I__4454\ : Span4Mux_h
    port map (
            O => \N__20780\,
            I => \N__20739\
        );

    \I__4453\ : Span4Mux_h
    port map (
            O => \N__20773\,
            I => \N__20736\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__20770\,
            I => \N__20725\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__20767\,
            I => \N__20725\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__20764\,
            I => \N__20725\
        );

    \I__4449\ : Span4Mux_v
    port map (
            O => \N__20759\,
            I => \N__20725\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20725\
        );

    \I__4447\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20720\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20720\
        );

    \I__4445\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20717\
        );

    \I__4444\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20712\
        );

    \I__4443\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20712\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__20748\,
            I => \beamYZ0Z_2\
        );

    \I__4441\ : Odrv4
    port map (
            O => \N__20745\,
            I => \beamYZ0Z_2\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__20742\,
            I => \beamYZ0Z_2\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__20739\,
            I => \beamYZ0Z_2\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__20736\,
            I => \beamYZ0Z_2\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__20725\,
            I => \beamYZ0Z_2\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20720\,
            I => \beamYZ0Z_2\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__20717\,
            I => \beamYZ0Z_2\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__20712\,
            I => \beamYZ0Z_2\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20682\
        );

    \I__4432\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20682\
        );

    \I__4431\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20682\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__20690\,
            I => \N__20679\
        );

    \I__4429\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20673\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20669\
        );

    \I__4427\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20664\
        );

    \I__4426\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20664\
        );

    \I__4425\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20659\
        );

    \I__4424\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20659\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20656\
        );

    \I__4422\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20653\
        );

    \I__4421\ : Span4Mux_s3_h
    port map (
            O => \N__20669\,
            I => \N__20648\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20648\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20641\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__20656\,
            I => \N__20641\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20641\
        );

    \I__4416\ : Span4Mux_h
    port map (
            O => \N__20648\,
            I => \N__20638\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__20641\,
            I => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__20638\,
            I => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__20633\,
            I => \un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__4411\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__20624\,
            I => charx_if_generate_plus_mult1_un61_sum_i
        );

    \I__4409\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20616\
        );

    \I__4408\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20613\
        );

    \I__4407\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20610\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20616\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__20613\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__20610\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0\
        );

    \I__4403\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20597\
        );

    \I__4402\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20597\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__20597\,
            I => charx_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__4400\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__20591\,
            I => \N_2096_i\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__4397\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__20582\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__4395\ : InMux
    port map (
            O => \N__20579\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__4394\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20569\
        );

    \I__4392\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20566\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__20569\,
            I => \N__20562\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20559\
        );

    \I__4389\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20556\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__20562\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__20559\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__20556\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__4385\ : CascadeMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__4384\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__20543\,
            I => \N__20540\
        );

    \I__4382\ : Odrv12
    port map (
            O => \N__20540\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__4380\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__20531\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__4378\ : InMux
    port map (
            O => \N__20528\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__20525\,
            I => \N__20521\
        );

    \I__4376\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__4375\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20515\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__20518\,
            I => \N__20510\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20510\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__20510\,
            I => column_1_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__4370\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__20501\,
            I => \N__20498\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__20498\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__4367\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__20492\,
            I => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__4365\ : InMux
    port map (
            O => \N__20489\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__4364\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__20480\,
            I => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__4361\ : InMux
    port map (
            O => \N__20477\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__4360\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__4359\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20468\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__20468\,
            I => column_1_i_i_3
        );

    \I__4357\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20459\
        );

    \I__4356\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20459\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__20459\,
            I => charx_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__4354\ : InMux
    port map (
            O => \N__20456\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__4353\ : InMux
    port map (
            O => \N__20453\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__4351\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__20444\,
            I => charx_if_generate_plus_mult1_un54_sum_i
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__4348\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__20435\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0\
        );

    \I__4346\ : InMux
    port map (
            O => \N__20432\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__4344\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__20423\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__4341\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__20414\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0\
        );

    \I__4339\ : InMux
    port map (
            O => \N__20411\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__4337\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__20402\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0\
        );

    \I__4335\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__20396\,
            I => charx_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__4333\ : InMux
    port map (
            O => \N__20393\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__4332\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__20387\,
            I => charx_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__4330\ : InMux
    port map (
            O => \N__20384\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__4329\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20376\
        );

    \I__4328\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20373\
        );

    \I__4327\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20370\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__20376\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__20373\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__20370\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0\
        );

    \I__4323\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__20357\,
            I => if_generate_plus_mult1_un54_sum_axb_2_l_fx
        );

    \I__4320\ : InMux
    port map (
            O => \N__20354\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__4319\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20345\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__20350\,
            I => \N__20341\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__20349\,
            I => \N__20338\
        );

    \I__4316\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20334\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20331\
        );

    \I__4314\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20328\
        );

    \I__4313\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20321\
        );

    \I__4312\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20321\
        );

    \I__4311\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20321\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__20334\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__20331\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__20328\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__20321\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__4305\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__20303\,
            I => if_generate_plus_mult1_un54_sum_axb_3_l_fx
        );

    \I__4302\ : InMux
    port map (
            O => \N__20300\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__4301\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20294\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__20294\,
            I => if_generate_plus_mult1_un54_sum_axb_4_l_fx
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__20291\,
            I => \N__20287\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__20290\,
            I => \N__20284\
        );

    \I__4297\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20279\
        );

    \I__4296\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20279\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20275\
        );

    \I__4294\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20272\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__20275\,
            I => \N_2110_i\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__20272\,
            I => \N_2110_i\
        );

    \I__4291\ : InMux
    port map (
            O => \N__20267\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__4290\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__20261\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__4288\ : InMux
    port map (
            O => \N__20258\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__20255\,
            I => \if_generate_plus_mult1_un54_sum_s_5_cascade_\
        );

    \I__4286\ : InMux
    port map (
            O => \N__20252\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__4285\ : InMux
    port map (
            O => \N__20249\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__4284\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__20243\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2\
        );

    \I__4282\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__20237\,
            I => column_1_if_generate_plus_mult1_un47_sum0_3
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__4279\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__20228\,
            I => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx
        );

    \I__4277\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__20222\,
            I => column_1_if_generate_plus_mult1_un47_sum0_2
        );

    \I__4275\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20211\
        );

    \I__4274\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20211\
        );

    \I__4273\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20200\
        );

    \I__4272\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20196\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20190\
        );

    \I__4270\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20187\
        );

    \I__4269\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20178\
        );

    \I__4268\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20178\
        );

    \I__4267\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20178\
        );

    \I__4266\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20178\
        );

    \I__4265\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20175\
        );

    \I__4264\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20170\
        );

    \I__4263\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20170\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20167\
        );

    \I__4261\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20164\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20158\
        );

    \I__4259\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20155\
        );

    \I__4258\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20150\
        );

    \I__4257\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20150\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__20190\,
            I => \N__20145\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__20187\,
            I => \N__20145\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20142\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__20175\,
            I => \N__20137\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__20170\,
            I => \N__20137\
        );

    \I__4251\ : Span4Mux_s1_h
    port map (
            O => \N__20167\,
            I => \N__20132\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20132\
        );

    \I__4249\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20125\
        );

    \I__4248\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20125\
        );

    \I__4247\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20125\
        );

    \I__4246\ : Sp12to4
    port map (
            O => \N__20158\,
            I => \N__20122\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__20155\,
            I => \N__20117\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20117\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__20145\,
            I => \N__20114\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__20142\,
            I => \N__20111\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__20137\,
            I => \N__20104\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__20132\,
            I => \N__20104\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20104\
        );

    \I__4238\ : Span12Mux_v
    port map (
            O => \N__20122\,
            I => \N__20099\
        );

    \I__4237\ : Span12Mux_s9_h
    port map (
            O => \N__20117\,
            I => \N__20099\
        );

    \I__4236\ : IoSpan4Mux
    port map (
            O => \N__20114\,
            I => \N__20096\
        );

    \I__4235\ : Span4Mux_h
    port map (
            O => \N__20111\,
            I => \N__20091\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__20104\,
            I => \N__20091\
        );

    \I__4233\ : Odrv12
    port map (
            O => \N__20099\,
            I => \SDATA1_c\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__20096\,
            I => \SDATA1_c\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__20091\,
            I => \SDATA1_c\
        );

    \I__4230\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__4228\ : Span4Mux_v
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__20075\,
            I => \N__20071\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20068\
        );

    \I__4225\ : Span4Mux_v
    port map (
            O => \N__20071\,
            I => \N__20063\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__20068\,
            I => \N__20063\
        );

    \I__4223\ : Span4Mux_h
    port map (
            O => \N__20063\,
            I => \N__20058\
        );

    \I__4222\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20052\
        );

    \I__4221\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20052\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__20058\,
            I => \N__20049\
        );

    \I__4219\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20046\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__20052\,
            I => un1_sclk17_9_0_3
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__20049\,
            I => un1_sclk17_9_0_3
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__20046\,
            I => un1_sclk17_9_0_3
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__4214\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__20021\,
            I => un1_sclk17_5_1_0
        );

    \I__4208\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__4206\ : Span4Mux_h
    port map (
            O => \N__20012\,
            I => \N__20008\
        );

    \I__4205\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20005\,
            I => \ScreenBuffer_0_9Z0Z_0\
        );

    \I__4202\ : Odrv4
    port map (
            O => \N__20002\,
            I => \ScreenBuffer_0_9Z0Z_0\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19990\
        );

    \I__4199\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19987\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__19987\,
            I => \N__19957\
        );

    \I__4196\ : Glb2LocalMux
    port map (
            O => \N__19984\,
            I => \N__19892\
        );

    \I__4195\ : ClkMux
    port map (
            O => \N__19983\,
            I => \N__19892\
        );

    \I__4194\ : ClkMux
    port map (
            O => \N__19982\,
            I => \N__19892\
        );

    \I__4193\ : ClkMux
    port map (
            O => \N__19981\,
            I => \N__19892\
        );

    \I__4192\ : ClkMux
    port map (
            O => \N__19980\,
            I => \N__19892\
        );

    \I__4191\ : ClkMux
    port map (
            O => \N__19979\,
            I => \N__19892\
        );

    \I__4190\ : ClkMux
    port map (
            O => \N__19978\,
            I => \N__19892\
        );

    \I__4189\ : ClkMux
    port map (
            O => \N__19977\,
            I => \N__19892\
        );

    \I__4188\ : ClkMux
    port map (
            O => \N__19976\,
            I => \N__19892\
        );

    \I__4187\ : ClkMux
    port map (
            O => \N__19975\,
            I => \N__19892\
        );

    \I__4186\ : ClkMux
    port map (
            O => \N__19974\,
            I => \N__19892\
        );

    \I__4185\ : ClkMux
    port map (
            O => \N__19973\,
            I => \N__19892\
        );

    \I__4184\ : ClkMux
    port map (
            O => \N__19972\,
            I => \N__19892\
        );

    \I__4183\ : ClkMux
    port map (
            O => \N__19971\,
            I => \N__19892\
        );

    \I__4182\ : ClkMux
    port map (
            O => \N__19970\,
            I => \N__19892\
        );

    \I__4181\ : ClkMux
    port map (
            O => \N__19969\,
            I => \N__19892\
        );

    \I__4180\ : ClkMux
    port map (
            O => \N__19968\,
            I => \N__19892\
        );

    \I__4179\ : ClkMux
    port map (
            O => \N__19967\,
            I => \N__19892\
        );

    \I__4178\ : ClkMux
    port map (
            O => \N__19966\,
            I => \N__19892\
        );

    \I__4177\ : ClkMux
    port map (
            O => \N__19965\,
            I => \N__19892\
        );

    \I__4176\ : ClkMux
    port map (
            O => \N__19964\,
            I => \N__19892\
        );

    \I__4175\ : ClkMux
    port map (
            O => \N__19963\,
            I => \N__19892\
        );

    \I__4174\ : ClkMux
    port map (
            O => \N__19962\,
            I => \N__19892\
        );

    \I__4173\ : ClkMux
    port map (
            O => \N__19961\,
            I => \N__19892\
        );

    \I__4172\ : ClkMux
    port map (
            O => \N__19960\,
            I => \N__19892\
        );

    \I__4171\ : Glb2LocalMux
    port map (
            O => \N__19957\,
            I => \N__19892\
        );

    \I__4170\ : ClkMux
    port map (
            O => \N__19956\,
            I => \N__19892\
        );

    \I__4169\ : ClkMux
    port map (
            O => \N__19955\,
            I => \N__19892\
        );

    \I__4168\ : ClkMux
    port map (
            O => \N__19954\,
            I => \N__19892\
        );

    \I__4167\ : ClkMux
    port map (
            O => \N__19953\,
            I => \N__19892\
        );

    \I__4166\ : GlobalMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4165\ : gio2CtrlBuf
    port map (
            O => \N__19889\,
            I => \Clock12MHz_c_g\
        );

    \I__4164\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__19883\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4\
        );

    \I__4162\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__19874\,
            I => column_1_if_generate_plus_mult1_un47_sum0_4
        );

    \I__4159\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__19868\,
            I => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx
        );

    \I__4157\ : InMux
    port map (
            O => \N__19865\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_1
        );

    \I__4156\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__19859\,
            I => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__4153\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__19850\,
            I => if_generate_plus_mult1_un47_sum_0_cry_3_ma
        );

    \I__4151\ : InMux
    port map (
            O => \N__19847\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_2
        );

    \I__4150\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N_1184_0_i\
        );

    \I__4148\ : InMux
    port map (
            O => \N__19838\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_3
        );

    \I__4147\ : InMux
    port map (
            O => \N__19835\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_4
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__4145\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__19826\,
            I => un5_visiblex_i_25
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \N_2110_i_cascade_\
        );

    \I__4142\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19814\
        );

    \I__4141\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19814\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__19814\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__19811\,
            I => \un115_pixel_6_bm_2_cascade_\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4136\ : Odrv12
    port map (
            O => \N__19802\,
            I => \N_1330\
        );

    \I__4135\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__19796\,
            I => un115_pixel_6_am_2
        );

    \I__4133\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19789\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__19792\,
            I => \N__19786\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__19789\,
            I => \N__19783\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19786\,
            I => \N__19780\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__19783\,
            I => un5_visiblex_i_24
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__19780\,
            I => un5_visiblex_i_24
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4126\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4124\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__19763\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0\
        );

    \I__4122\ : InMux
    port map (
            O => \N__19760\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \N__19753\
        );

    \I__4120\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19748\
        );

    \I__4119\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19748\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__19742\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0\
        );

    \I__4115\ : InMux
    port map (
            O => \N__19739\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__4114\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4112\ : Span4Mux_h
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__19727\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__4110\ : InMux
    port map (
            O => \N__19724\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__4109\ : InMux
    port map (
            O => \N__19721\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__4108\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19712\
        );

    \I__4107\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19709\
        );

    \I__4106\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19706\
        );

    \I__4105\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19703\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19698\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19698\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19691\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19691\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__19698\,
            I => \N__19691\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__19691\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0\
        );

    \I__4098\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__19685\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \N__19678\
        );

    \I__4095\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19670\
        );

    \I__4094\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19670\
        );

    \I__4093\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19670\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__19670\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__19667\,
            I => \m14_cascade_\
        );

    \I__4090\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__19661\,
            I => \beamY_RNI7RM4IFZ0Z_0\
        );

    \I__4088\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__19655\,
            I => \un113_pixel_3_0_11__g1_1_0\
        );

    \I__4086\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__19649\,
            I => \beamY_RNIPQEDM42Z0Z_0\
        );

    \I__4084\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N_1293\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__19640\,
            I => \N_1306_cascade_\
        );

    \I__4081\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N_1327_0\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__19631\,
            I => \m11_cascade_\
        );

    \I__4078\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__19625\,
            I => \un113_pixel_4_0_15__N_17\
        );

    \I__4076\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__19619\,
            I => un115_pixel_4_am_7
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__19616\,
            I => \N_1287_cascade_\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__19613\,
            I => \currentchar_1_0_cascade_\
        );

    \I__4072\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__19607\,
            I => un115_pixel_4_bm_7
        );

    \I__4070\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19595\
        );

    \I__4068\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19590\
        );

    \I__4067\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19590\
        );

    \I__4066\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19587\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__19595\,
            I => \ScreenBuffer_0_7_RNII0GVLQZ0Z_0\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__19590\,
            I => \ScreenBuffer_0_7_RNII0GVLQZ0Z_0\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__19587\,
            I => \ScreenBuffer_0_7_RNII0GVLQZ0Z_0\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__19580\,
            I => \un113_pixel_1_0_3__N_10_mux_cascade_\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__19577\,
            I => \N_1285_0_0_0_cascade_\
        );

    \I__4060\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__19562\,
            I => \un113_pixel_3_0_11__g1_0_0_0\
        );

    \I__4055\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__19556\,
            I => m14
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__19550\,
            I => \currentchar_m7_0_cascade_\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__19547\,
            I => \N__19543\
        );

    \I__4050\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19540\
        );

    \I__4049\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19537\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19529\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__19534\,
            I => \N__19529\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__19529\,
            I => \ScreenBuffer_0_7Z0Z_0\
        );

    \I__4044\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19522\
        );

    \I__4043\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__19519\,
            I => \ScreenBuffer_0_5Z0Z_0\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__19516\,
            I => \ScreenBuffer_0_5Z0Z_0\
        );

    \I__4039\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19507\
        );

    \I__4038\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__19507\,
            I => \N__19500\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__19504\,
            I => \N__19497\
        );

    \I__4035\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19494\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__19500\,
            I => \un113_pixel_3_0_11__currentchar_N_13\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__19497\,
            I => \un113_pixel_3_0_11__currentchar_N_13\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__19494\,
            I => \un113_pixel_3_0_11__currentchar_N_13\
        );

    \I__4031\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__19484\,
            I => un112_pixel_1_2_x1
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \un112_pixel_2_8_cascade_\
        );

    \I__4028\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__19472\,
            I => \ScreenBuffer_1_2Z0Z_3\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__19469\,
            I => \un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__19466\,
            I => \un113_pixel_3_0_11__currentchar_N_13_cascade_\
        );

    \I__4023\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19459\
        );

    \I__4022\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19451\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__19456\,
            I => \N__19451\
        );

    \I__4019\ : Span12Mux_s11_v
    port map (
            O => \N__19451\,
            I => \N__19446\
        );

    \I__4018\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19443\
        );

    \I__4017\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19440\
        );

    \I__4016\ : Odrv12
    port map (
            O => \N__19446\,
            I => \voltage_3Z0Z_3\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__19443\,
            I => \voltage_3Z0Z_3\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__19440\,
            I => \voltage_3Z0Z_3\
        );

    \I__4013\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19429\
        );

    \I__4012\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__4009\ : Span4Mux_v
    port map (
            O => \N__19423\,
            I => \N__19413\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__19420\,
            I => \N__19413\
        );

    \I__4007\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19407\
        );

    \I__4006\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19407\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__19413\,
            I => \N__19404\
        );

    \I__4004\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19401\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19398\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__19404\,
            I => \voltage_0Z0Z_3\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__19401\,
            I => \voltage_0Z0Z_3\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__19398\,
            I => \voltage_0Z0Z_3\
        );

    \I__3999\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__19388\,
            I => \ScreenBuffer_1_0Z0Z_3\
        );

    \I__3997\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__19382\,
            I => \un113_pixel_4_0_15__g0_1Z0Z_0\
        );

    \I__3995\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__19376\,
            I => \un113_pixel_4_0_15__g0_3_0\
        );

    \I__3993\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19365\
        );

    \I__3991\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19362\
        );

    \I__3990\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19359\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__19365\,
            I => \N__19356\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__19362\,
            I => \N__19353\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19349\
        );

    \I__3986\ : Span4Mux_h
    port map (
            O => \N__19356\,
            I => \N__19344\
        );

    \I__3985\ : Span4Mux_s3_h
    port map (
            O => \N__19353\,
            I => \N__19344\
        );

    \I__3984\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19341\
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__19349\,
            I => \voltage_3Z0Z_1\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__19344\,
            I => \voltage_3Z0Z_1\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__19341\,
            I => \voltage_3Z0Z_1\
        );

    \I__3980\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19323\
        );

    \I__3979\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19315\
        );

    \I__3978\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19310\
        );

    \I__3977\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19310\
        );

    \I__3976\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19296\
        );

    \I__3975\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19293\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__19328\,
            I => \N__19285\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__19327\,
            I => \N__19281\
        );

    \I__3972\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19277\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__19323\,
            I => \N__19274\
        );

    \I__3970\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19265\
        );

    \I__3969\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19265\
        );

    \I__3968\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19265\
        );

    \I__3967\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19265\
        );

    \I__3966\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19262\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__19315\,
            I => \N__19257\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__19310\,
            I => \N__19257\
        );

    \I__3963\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19252\
        );

    \I__3962\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19252\
        );

    \I__3961\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19243\
        );

    \I__3960\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19243\
        );

    \I__3959\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19234\
        );

    \I__3958\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19234\
        );

    \I__3957\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19234\
        );

    \I__3956\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19234\
        );

    \I__3955\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19229\
        );

    \I__3954\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19229\
        );

    \I__3953\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19226\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19221\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__19293\,
            I => \N__19221\
        );

    \I__3950\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19218\
        );

    \I__3949\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19213\
        );

    \I__3948\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19213\
        );

    \I__3947\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19210\
        );

    \I__3946\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19203\
        );

    \I__3945\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19203\
        );

    \I__3944\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19203\
        );

    \I__3943\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19198\
        );

    \I__3942\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19198\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__19277\,
            I => \N__19187\
        );

    \I__3940\ : Span4Mux_h
    port map (
            O => \N__19274\,
            I => \N__19187\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19187\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__19262\,
            I => \N__19187\
        );

    \I__3937\ : Span4Mux_s3_v
    port map (
            O => \N__19257\,
            I => \N__19187\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__19252\,
            I => \N__19184\
        );

    \I__3935\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19167\
        );

    \I__3934\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19167\
        );

    \I__3933\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19167\
        );

    \I__3932\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19167\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__19243\,
            I => \N__19146\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__19234\,
            I => \N__19146\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__19229\,
            I => \N__19146\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19146\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__19221\,
            I => \N__19146\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19146\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__19213\,
            I => \N__19146\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19146\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__19203\,
            I => \N__19146\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__19198\,
            I => \N__19146\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__19187\,
            I => \N__19143\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__19184\,
            I => \N__19140\
        );

    \I__3919\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19135\
        );

    \I__3918\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19135\
        );

    \I__3917\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19132\
        );

    \I__3916\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19127\
        );

    \I__3915\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19127\
        );

    \I__3914\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19124\
        );

    \I__3913\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19121\
        );

    \I__3912\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19118\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__19167\,
            I => \N__19115\
        );

    \I__3910\ : Span4Mux_v
    port map (
            O => \N__19146\,
            I => \N__19107\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__19143\,
            I => \N__19102\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__19140\,
            I => \N__19102\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__19135\,
            I => \N__19093\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19093\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19093\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19093\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19086\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19086\
        );

    \I__3901\ : Span4Mux_h
    port map (
            O => \N__19115\,
            I => \N__19086\
        );

    \I__3900\ : InMux
    port map (
            O => \N__19114\,
            I => \N__19081\
        );

    \I__3899\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19081\
        );

    \I__3898\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19074\
        );

    \I__3897\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19074\
        );

    \I__3896\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19074\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__19107\,
            I => \N__19071\
        );

    \I__3894\ : Sp12to4
    port map (
            O => \N__19102\,
            I => \N__19066\
        );

    \I__3893\ : Span12Mux_s11_v
    port map (
            O => \N__19093\,
            I => \N__19066\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__19086\,
            I => \N__19063\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__19081\,
            I => \slaveselectZ0\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__19074\,
            I => \slaveselectZ0\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__19071\,
            I => \slaveselectZ0\
        );

    \I__3888\ : Odrv12
    port map (
            O => \N__19066\,
            I => \slaveselectZ0\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__19063\,
            I => \slaveselectZ0\
        );

    \I__3886\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19048\
        );

    \I__3885\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19043\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19040\
        );

    \I__3883\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19037\
        );

    \I__3882\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19034\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__19031\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__19040\,
            I => \N__19027\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19024\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__19034\,
            I => \N__19021\
        );

    \I__3877\ : Span4Mux_v
    port map (
            O => \N__19031\,
            I => \N__19018\
        );

    \I__3876\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19015\
        );

    \I__3875\ : Span4Mux_h
    port map (
            O => \N__19027\,
            I => \N__19010\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__19024\,
            I => \N__19010\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__19021\,
            I => \N__19005\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__19018\,
            I => \N__19005\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__19015\,
            I => \voltage_0Z0Z_1\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__19010\,
            I => \voltage_0Z0Z_1\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__19005\,
            I => \voltage_0Z0Z_1\
        );

    \I__3868\ : CEMux
    port map (
            O => \N__18998\,
            I => \N__18994\
        );

    \I__3867\ : CEMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__18985\,
            I => \N__18979\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__18982\,
            I => \un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__18979\,
            I => \un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0\
        );

    \I__3860\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18970\
        );

    \I__3859\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18967\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__18967\,
            I => \ScreenBuffer_0_12Z0Z_0\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__18964\,
            I => \ScreenBuffer_0_12Z0Z_0\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18955\
        );

    \I__3854\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__18952\,
            I => \ScreenBuffer_0_4Z0Z_0\
        );

    \I__3851\ : Odrv12
    port map (
            O => \N__18949\,
            I => \ScreenBuffer_0_4Z0Z_0\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__18944\,
            I => \ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18937\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__3846\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18928\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__18928\,
            I => \ScreenBuffer_0_6Z0Z_0\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__18925\,
            I => \ScreenBuffer_0_6Z0Z_0\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \beamY_RNIOEPPEK1Z0Z_0_cascade_\
        );

    \I__3841\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__18914\,
            I => un112_pixel_1_2
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__18911\,
            I => \N_3461_0_cascade_\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__18908\,
            I => \N_4568_0_cascade_\
        );

    \I__3837\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N_1305_0\
        );

    \I__3835\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__18896\,
            I => \un113_pixel_4_0_15__g0_0Z0Z_2\
        );

    \I__3833\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__3831\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__18884\,
            I => \Pixel_3_sqmuxa_0\
        );

    \I__3829\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__18878\,
            I => g0_1_1
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__18875\,
            I => \N_1_0_cascade_\
        );

    \I__3826\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__3824\ : Odrv12
    port map (
            O => \N__18866\,
            I => \ScreenBuffer_1_3Z0Z_3\
        );

    \I__3823\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__18854\,
            I => \ScreenBuffer_1_1Z0Z_3\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__3818\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__18845\,
            I => \column_1_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__3815\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18835\
        );

    \I__3814\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18832\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__18835\,
            I => chary_24
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__18832\,
            I => chary_24
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__3810\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__18818\,
            I => \un113_pixel_4_0_15__gZ0Z2\
        );

    \I__3807\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18811\
        );

    \I__3806\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__18811\,
            I => font_un3_pixel_30
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__18808\,
            I => font_un3_pixel_30
        );

    \I__3803\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__18800\,
            I => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__18797\,
            I => \font_un57_pixel_cascade_\
        );

    \I__3800\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__18791\,
            I => currentchar_1_5
        );

    \I__3798\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__18782\,
            I => font_un67_pixel_ac0_5
        );

    \I__3795\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__18776\,
            I => font_un64_pixel_ac0_5
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__18773\,
            I => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_\
        );

    \I__3792\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__18761\,
            I => \N_12\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__18749\,
            I => \un113_pixel_4_0_15__g0_iZ0Z_2\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__18746\,
            I => \un113_pixel_4_0_15__g0_iZ0Z_5_cascade_\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__18743\,
            I => \N__18737\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__18742\,
            I => \N__18733\
        );

    \I__3781\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18726\
        );

    \I__3780\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18726\
        );

    \I__3779\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18726\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__18736\,
            I => \N__18721\
        );

    \I__3777\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18717\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18714\
        );

    \I__3775\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18711\
        );

    \I__3774\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18708\
        );

    \I__3773\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18705\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \N__18701\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__18717\,
            I => \N__18695\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__18714\,
            I => \N__18692\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18687\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18687\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__18705\,
            I => \N__18684\
        );

    \I__3766\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18679\
        );

    \I__3765\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18679\
        );

    \I__3764\ : InMux
    port map (
            O => \N__18700\,
            I => \N__18676\
        );

    \I__3763\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18673\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18670\
        );

    \I__3761\ : Span4Mux_s2_v
    port map (
            O => \N__18695\,
            I => \N__18667\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__18692\,
            I => \N__18664\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__18687\,
            I => \N__18661\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__18684\,
            I => \N__18656\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__18679\,
            I => \N__18656\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__18676\,
            I => \N__18653\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__18673\,
            I => \beamXZ0Z_0\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__18670\,
            I => \beamXZ0Z_0\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__18667\,
            I => \beamXZ0Z_0\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__18664\,
            I => \beamXZ0Z_0\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__18661\,
            I => \beamXZ0Z_0\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__18656\,
            I => \beamXZ0Z_0\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__18653\,
            I => \beamXZ0Z_0\
        );

    \I__3748\ : InMux
    port map (
            O => \N__18638\,
            I => \N__18632\
        );

    \I__3747\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18632\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__18632\,
            I => \un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6\
        );

    \I__3745\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18623\
        );

    \I__3744\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18623\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__18623\,
            I => charx_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__3742\ : InMux
    port map (
            O => \N__18620\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__3741\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18602\
        );

    \I__3740\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18602\
        );

    \I__3739\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18602\
        );

    \I__3738\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18602\
        );

    \I__3737\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18602\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__18602\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__3734\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__18593\,
            I => charx_if_generate_plus_mult1_un68_sum_i
        );

    \I__3732\ : InMux
    port map (
            O => \N__18590\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__3731\ : InMux
    port map (
            O => \N__18587\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__3730\ : InMux
    port map (
            O => \N__18584\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__3729\ : InMux
    port map (
            O => \N__18581\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__3728\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18572\
        );

    \I__3727\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18572\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__18569\,
            I => \N__18565\
        );

    \I__3724\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18562\
        );

    \I__3723\ : Span4Mux_h
    port map (
            O => \N__18565\,
            I => \N__18559\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__18562\,
            I => \N__18556\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__18559\,
            I => \N__18551\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__18556\,
            I => \N__18551\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__18551\,
            I => un1_counter_1_0
        );

    \I__3718\ : SRMux
    port map (
            O => \N__18548\,
            I => \N__18524\
        );

    \I__3717\ : SRMux
    port map (
            O => \N__18547\,
            I => \N__18524\
        );

    \I__3716\ : SRMux
    port map (
            O => \N__18546\,
            I => \N__18524\
        );

    \I__3715\ : SRMux
    port map (
            O => \N__18545\,
            I => \N__18524\
        );

    \I__3714\ : SRMux
    port map (
            O => \N__18544\,
            I => \N__18524\
        );

    \I__3713\ : SRMux
    port map (
            O => \N__18543\,
            I => \N__18524\
        );

    \I__3712\ : SRMux
    port map (
            O => \N__18542\,
            I => \N__18524\
        );

    \I__3711\ : SRMux
    port map (
            O => \N__18541\,
            I => \N__18524\
        );

    \I__3710\ : GlobalMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__3709\ : gio2CtrlBuf
    port map (
            O => \N__18521\,
            I => voltage_0_0_sqmuxa_1_g
        );

    \I__3708\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__3705\ : Span4Mux_h
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__3704\ : Span4Mux_h
    port map (
            O => \N__18506\,
            I => \N__18500\
        );

    \I__3703\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18497\
        );

    \I__3702\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18494\
        );

    \I__3701\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18491\
        );

    \I__3700\ : Odrv4
    port map (
            O => \N__18500\,
            I => \voltage_3Z0Z_0\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__18497\,
            I => \voltage_3Z0Z_0\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__18494\,
            I => \voltage_3Z0Z_0\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__18491\,
            I => \voltage_3Z0Z_0\
        );

    \I__3696\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18469\
        );

    \I__3695\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18469\
        );

    \I__3694\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18469\
        );

    \I__3693\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18469\
        );

    \I__3692\ : InMux
    port map (
            O => \N__18478\,
            I => \N__18466\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18460\
        );

    \I__3689\ : Span4Mux_s3_h
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__18460\,
            I => \N__18453\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__18457\,
            I => \N__18450\
        );

    \I__3686\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18447\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__18453\,
            I => \N__18444\
        );

    \I__3684\ : Span4Mux_v
    port map (
            O => \N__18450\,
            I => \N__18441\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__18447\,
            I => \voltage_0Z0Z_0\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__18444\,
            I => \voltage_0Z0Z_0\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__18441\,
            I => \voltage_0Z0Z_0\
        );

    \I__3680\ : CEMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18427\
        );

    \I__3678\ : CEMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__3677\ : Span4Mux_h
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__18421\,
            I => \N__18415\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__18415\,
            I => \un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__18412\,
            I => \un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18403\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__18406\,
            I => \N__18399\
        );

    \I__3669\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18389\
        );

    \I__3668\ : InMux
    port map (
            O => \N__18402\,
            I => \N__18389\
        );

    \I__3667\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18389\
        );

    \I__3666\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18389\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__18389\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__3664\ : InMux
    port map (
            O => \N__18386\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__3663\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18374\
        );

    \I__3662\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18374\
        );

    \I__3661\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18374\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__18374\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1\
        );

    \I__3659\ : InMux
    port map (
            O => \N__18371\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__3658\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18364\
        );

    \I__3657\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18361\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__18364\,
            I => \N__18354\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18354\
        );

    \I__3654\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18351\
        );

    \I__3653\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18348\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__18354\,
            I => \N__18343\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__18351\,
            I => \N__18343\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__18348\,
            I => \beamXZ0Z_8\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__18343\,
            I => \beamXZ0Z_8\
        );

    \I__3648\ : InMux
    port map (
            O => \N__18338\,
            I => \bfn_8_4_0_\
        );

    \I__3647\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18331\
        );

    \I__3646\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18328\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18321\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18321\
        );

    \I__3643\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__3642\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18315\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__18321\,
            I => \N__18310\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18310\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__18315\,
            I => \beamXZ0Z_9\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__18310\,
            I => \beamXZ0Z_9\
        );

    \I__3637\ : InMux
    port map (
            O => \N__18305\,
            I => un5_visiblex_cry_8
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \CO3_0_cascade_\
        );

    \I__3635\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__18296\,
            I => charx_if_generate_plus_mult1_un26_sum_s_2_sf
        );

    \I__3633\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18288\
        );

    \I__3632\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18280\
        );

    \I__3631\ : InMux
    port map (
            O => \N__18291\,
            I => \N__18277\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18274\
        );

    \I__3629\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18271\
        );

    \I__3628\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18266\
        );

    \I__3627\ : InMux
    port map (
            O => \N__18285\,
            I => \N__18266\
        );

    \I__3626\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18263\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__18283\,
            I => \N__18257\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18250\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__18277\,
            I => \N__18247\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__18274\,
            I => \N__18242\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18242\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__18266\,
            I => \N__18237\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__18263\,
            I => \N__18237\
        );

    \I__3618\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18230\
        );

    \I__3617\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18230\
        );

    \I__3616\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18230\
        );

    \I__3615\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18227\
        );

    \I__3614\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18213\
        );

    \I__3613\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18213\
        );

    \I__3612\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18213\
        );

    \I__3611\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18213\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__18250\,
            I => \N__18202\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__18247\,
            I => \N__18202\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__18242\,
            I => \N__18202\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__18237\,
            I => \N__18202\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__18230\,
            I => \N__18202\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18199\
        );

    \I__3604\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18196\
        );

    \I__3603\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18193\
        );

    \I__3602\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18186\
        );

    \I__3601\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18186\
        );

    \I__3600\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18186\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18183\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__18202\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__18199\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__18196\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__18193\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__18186\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__18183\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3592\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18165\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__18169\,
            I => \N__18159\
        );

    \I__3590\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18154\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__18165\,
            I => \N__18151\
        );

    \I__3588\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18146\
        );

    \I__3587\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18146\
        );

    \I__3586\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18143\
        );

    \I__3585\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18132\
        );

    \I__3584\ : InMux
    port map (
            O => \N__18158\,
            I => \N__18129\
        );

    \I__3583\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18126\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__18154\,
            I => \N__18121\
        );

    \I__3581\ : Span4Mux_v
    port map (
            O => \N__18151\,
            I => \N__18121\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18116\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__18143\,
            I => \N__18116\
        );

    \I__3578\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18109\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18109\
        );

    \I__3576\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18109\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__18139\,
            I => \N__18103\
        );

    \I__3574\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18093\
        );

    \I__3573\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18093\
        );

    \I__3572\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18093\
        );

    \I__3571\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18093\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__18132\,
            I => \N__18088\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__18129\,
            I => \N__18088\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__18126\,
            I => \N__18085\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__18121\,
            I => \N__18078\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__18116\,
            I => \N__18078\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__18109\,
            I => \N__18078\
        );

    \I__3564\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18073\
        );

    \I__3563\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18073\
        );

    \I__3562\ : InMux
    port map (
            O => \N__18106\,
            I => \N__18066\
        );

    \I__3561\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18066\
        );

    \I__3560\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18066\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__18093\,
            I => \N__18063\
        );

    \I__3558\ : Odrv12
    port map (
            O => \N__18088\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__18085\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__18078\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__18073\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__18066\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__18063\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__3551\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N_13\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__3548\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__18032\,
            I => \N__18029\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__18029\,
            I => \un113_pixel_4_0_15__un4_rowZ0Z_1\
        );

    \I__3544\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18023\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__18011\,
            I => un1_voltage_0_axb_0
        );

    \I__3538\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__17993\,
            I => voltage_0_10_iv_0_0
        );

    \I__3532\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17984\
        );

    \I__3531\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17984\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__17984\,
            I => \N__17980\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__17983\,
            I => \N__17977\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__17980\,
            I => \N__17973\
        );

    \I__3527\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17970\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17967\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__17973\,
            I => \N__17964\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__17970\,
            I => un1_voltage_012_2_0
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__17967\,
            I => un1_voltage_012_2_0
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__17964\,
            I => un1_voltage_012_2_0
        );

    \I__3521\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__3519\ : Span12Mux_s10_h
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__3518\ : Odrv12
    port map (
            O => \N__17948\,
            I => voltage_0_10_iv_0_1
        );

    \I__3517\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__3515\ : Span12Mux_s8_v
    port map (
            O => \N__17939\,
            I => \N__17936\
        );

    \I__3514\ : Odrv12
    port map (
            O => \N__17936\,
            I => \voltage_0_RNO_0Z0Z_1\
        );

    \I__3513\ : IoInMux
    port map (
            O => \N__17933\,
            I => \N__17929\
        );

    \I__3512\ : IoInMux
    port map (
            O => \N__17932\,
            I => \N__17926\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__17929\,
            I => \N__17921\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17921\
        );

    \I__3509\ : Span4Mux_s3_v
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__3507\ : Span4Mux_v
    port map (
            O => \N__17915\,
            I => \N__17911\
        );

    \I__3506\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17908\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__17911\,
            I => \nCS1_c\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__17908\,
            I => \nCS1_c\
        );

    \I__3503\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17897\
        );

    \I__3502\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17892\
        );

    \I__3501\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17892\
        );

    \I__3500\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17888\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17885\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__17892\,
            I => \N__17882\
        );

    \I__3497\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17879\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__17888\,
            I => \beamXZ0Z_1\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__17885\,
            I => \beamXZ0Z_1\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__17882\,
            I => \beamXZ0Z_1\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__17879\,
            I => \beamXZ0Z_1\
        );

    \I__3492\ : InMux
    port map (
            O => \N__17870\,
            I => un5_visiblex_cry_0
        );

    \I__3491\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17861\
        );

    \I__3490\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17861\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17856\
        );

    \I__3488\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17853\
        );

    \I__3487\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17850\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__17856\,
            I => \N__17847\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__17853\,
            I => \N__17844\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__17850\,
            I => \beamXZ0Z_2\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__17847\,
            I => \beamXZ0Z_2\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__17844\,
            I => \beamXZ0Z_2\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17837\,
            I => un5_visiblex_cry_1
        );

    \I__3480\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17825\
        );

    \I__3478\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17820\
        );

    \I__3477\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17820\
        );

    \I__3476\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17816\
        );

    \I__3475\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17811\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__17820\,
            I => \N__17811\
        );

    \I__3473\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17808\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17803\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__17811\,
            I => \N__17803\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17800\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__17803\,
            I => \beamXZ0Z_3\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__17800\,
            I => \beamXZ0Z_3\
        );

    \I__3467\ : InMux
    port map (
            O => \N__17795\,
            I => un5_visiblex_cry_2
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__17792\,
            I => \N__17787\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \N__17784\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__17790\,
            I => \N__17780\
        );

    \I__3463\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17777\
        );

    \I__3462\ : InMux
    port map (
            O => \N__17784\,
            I => \N__17772\
        );

    \I__3461\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17772\
        );

    \I__3460\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17769\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__17777\,
            I => \N__17764\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__17772\,
            I => \N__17764\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__17769\,
            I => \N__17759\
        );

    \I__3456\ : Span4Mux_h
    port map (
            O => \N__17764\,
            I => \N__17756\
        );

    \I__3455\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17753\
        );

    \I__3454\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17750\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17747\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__17756\,
            I => \N__17744\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17741\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__17750\,
            I => \beamXZ0Z_4\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__17747\,
            I => \beamXZ0Z_4\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__17744\,
            I => \beamXZ0Z_4\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__17741\,
            I => \beamXZ0Z_4\
        );

    \I__3446\ : InMux
    port map (
            O => \N__17732\,
            I => un5_visiblex_cry_3
        );

    \I__3445\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17717\
        );

    \I__3444\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17717\
        );

    \I__3443\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17717\
        );

    \I__3442\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17717\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__17714\,
            I => \N__17709\
        );

    \I__3439\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17706\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17703\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__17709\,
            I => \N__17700\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__17706\,
            I => \N__17697\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__17703\,
            I => \beamXZ0Z_5\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__17700\,
            I => \beamXZ0Z_5\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__17697\,
            I => \beamXZ0Z_5\
        );

    \I__3432\ : InMux
    port map (
            O => \N__17690\,
            I => un5_visiblex_cry_4
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \N__17681\
        );

    \I__3430\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17676\
        );

    \I__3429\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17673\
        );

    \I__3428\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17668\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17668\
        );

    \I__3426\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17665\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__17679\,
            I => \N__17662\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__17676\,
            I => \N__17658\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__17673\,
            I => \N__17653\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17653\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17650\
        );

    \I__3420\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17647\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17644\
        );

    \I__3418\ : Span4Mux_v
    port map (
            O => \N__17658\,
            I => \N__17641\
        );

    \I__3417\ : Span12Mux_s7_h
    port map (
            O => \N__17653\,
            I => \N__17638\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__17650\,
            I => \N__17633\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17633\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__17644\,
            I => \beamXZ0Z_6\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__17641\,
            I => \beamXZ0Z_6\
        );

    \I__3412\ : Odrv12
    port map (
            O => \N__17638\,
            I => \beamXZ0Z_6\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__17633\,
            I => \beamXZ0Z_6\
        );

    \I__3410\ : InMux
    port map (
            O => \N__17624\,
            I => un5_visiblex_cry_5
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__17621\,
            I => \N__17616\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__17620\,
            I => \N__17611\
        );

    \I__3407\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17608\
        );

    \I__3406\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17601\
        );

    \I__3405\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17601\
        );

    \I__3404\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17601\
        );

    \I__3403\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17598\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__17608\,
            I => \N__17591\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__17601\,
            I => \N__17591\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__17598\,
            I => \N__17588\
        );

    \I__3399\ : InMux
    port map (
            O => \N__17597\,
            I => \N__17585\
        );

    \I__3398\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17582\
        );

    \I__3397\ : Span12Mux_v
    port map (
            O => \N__17591\,
            I => \N__17579\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__17588\,
            I => \N__17576\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__17585\,
            I => \N__17573\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__17582\,
            I => \beamXZ0Z_7\
        );

    \I__3393\ : Odrv12
    port map (
            O => \N__17579\,
            I => \beamXZ0Z_7\
        );

    \I__3392\ : Odrv4
    port map (
            O => \N__17576\,
            I => \beamXZ0Z_7\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__17573\,
            I => \beamXZ0Z_7\
        );

    \I__3390\ : InMux
    port map (
            O => \N__17564\,
            I => un5_visiblex_cry_6
        );

    \I__3389\ : InMux
    port map (
            O => \N__17561\,
            I => un8_beamx_cry_4
        );

    \I__3388\ : InMux
    port map (
            O => \N__17558\,
            I => un8_beamx_cry_5
        );

    \I__3387\ : InMux
    port map (
            O => \N__17555\,
            I => un8_beamx_cry_6
        );

    \I__3386\ : InMux
    port map (
            O => \N__17552\,
            I => un8_beamx_cry_7
        );

    \I__3385\ : InMux
    port map (
            O => \N__17549\,
            I => \bfn_8_2_0_\
        );

    \I__3384\ : CEMux
    port map (
            O => \N__17546\,
            I => \N__17542\
        );

    \I__3383\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17537\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__17542\,
            I => \N__17534\
        );

    \I__3381\ : CEMux
    port map (
            O => \N__17541\,
            I => \N__17530\
        );

    \I__3380\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17526\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17523\
        );

    \I__3378\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17520\
        );

    \I__3377\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17516\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__17530\,
            I => \N__17513\
        );

    \I__3375\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17510\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__17526\,
            I => \N__17507\
        );

    \I__3373\ : Span4Mux_h
    port map (
            O => \N__17523\,
            I => \N__17504\
        );

    \I__3372\ : Span4Mux_s1_h
    port map (
            O => \N__17520\,
            I => \N__17501\
        );

    \I__3371\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17498\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__17516\,
            I => \N__17495\
        );

    \I__3369\ : Span4Mux_s2_h
    port map (
            O => \N__17513\,
            I => \N__17492\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17487\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__17507\,
            I => \N__17487\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__17504\,
            I => \N__17482\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__17501\,
            I => \N__17482\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__17498\,
            I => un3_beamx_0
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__17495\,
            I => un3_beamx_0
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__17492\,
            I => un3_beamx_0
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__17487\,
            I => un3_beamx_0
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__17482\,
            I => un3_beamx_0
        );

    \I__3359\ : InMux
    port map (
            O => \N__17471\,
            I => un8_beamx_cry_9
        );

    \I__3358\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17463\
        );

    \I__3357\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17459\
        );

    \I__3356\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17456\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__17463\,
            I => \N__17453\
        );

    \I__3354\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17450\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__17459\,
            I => \N__17445\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17445\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__17453\,
            I => \N__17442\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17437\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__17445\,
            I => \N__17437\
        );

    \I__3348\ : Span4Mux_v
    port map (
            O => \N__17442\,
            I => \N__17434\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__17437\,
            I => \beamXZ0Z_10\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__17434\,
            I => \beamXZ0Z_10\
        );

    \I__3345\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__17426\,
            I => \ScreenBuffer_0_7_RNIHMH43T2Z0Z_0\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__17423\,
            I => \beamY_RNIDQUNU91Z0Z_0_cascade_\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \un115_pixel_2_sn_5_cascade_\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \un112_pixel_7_cascade_\
        );

    \I__3340\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__17411\,
            I => \beamY_RNIINK7J73Z0Z_0\
        );

    \I__3338\ : InMux
    port map (
            O => \N__17408\,
            I => un8_beamx_cry_1
        );

    \I__3337\ : InMux
    port map (
            O => \N__17405\,
            I => un8_beamx_cry_2
        );

    \I__3336\ : InMux
    port map (
            O => \N__17402\,
            I => un8_beamx_cry_3
        );

    \I__3335\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__17393\,
            I => \slaveselect_RNILOQC2Z0Z_0\
        );

    \I__3332\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17386\
        );

    \I__3331\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__17383\,
            I => \ScreenBuffer_1_2Z0Z_4\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__17380\,
            I => \ScreenBuffer_1_2Z0Z_4\
        );

    \I__3327\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__17372\,
            I => \ScreenBuffer_1_3Z0Z_2\
        );

    \I__3325\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__3323\ : Span4Mux_v
    port map (
            O => \N__17363\,
            I => \N__17360\
        );

    \I__3322\ : Span4Mux_h
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__17357\,
            I => \ScreenBuffer_1_0Z0Z_2\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__17354\,
            I => \un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__17351\,
            I => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_\
        );

    \I__3318\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__17345\,
            I => m10_0_x1
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__17342\,
            I => \un112_pixel_2_2_cascade_\
        );

    \I__3315\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17336\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__17336\,
            I => \un113_pixel_3_0_11__g0_0Z0Z_0\
        );

    \I__3313\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17329\
        );

    \I__3312\ : InMux
    port map (
            O => \N__17332\,
            I => \N__17326\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__17329\,
            I => \N__17323\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__17326\,
            I => \N__17318\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__17323\,
            I => \N__17318\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__17318\,
            I => \ScreenBuffer_1_3Z0Z_4\
        );

    \I__3307\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__17312\,
            I => \ScreenBuffer_1_3_RNIVS9G2FZ0Z_4\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__17309\,
            I => \g1Z0Z_1_cascade_\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__17306\,
            I => \N_1428_0_cascade_\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__17303\,
            I => \un113_pixel_4_0_15__g1_1_cascade_\
        );

    \I__3302\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17297\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__17297\,
            I => \N_1300_0\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__17294\,
            I => \un112_pixel_0_2_cascade_\
        );

    \I__3299\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17288\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__17288\,
            I => \N_1293_0\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__17285\,
            I => \ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__17282\,
            I => \ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_\
        );

    \I__3295\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17273\
        );

    \I__3294\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17273\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17270\
        );

    \I__3292\ : Span12Mux_s7_h
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__3291\ : Odrv12
    port map (
            O => \N__17267\,
            I => row_1_if_generate_plus_mult1_un75_sum_c5
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__3289\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17255\
        );

    \I__3288\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17255\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17252\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__17252\,
            I => \N__17248\
        );

    \I__3285\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17245\
        );

    \I__3284\ : Sp12to4
    port map (
            O => \N__17248\,
            I => \N__17240\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17240\
        );

    \I__3282\ : Odrv12
    port map (
            O => \N__17240\,
            I => \row_1_if_generate_plus_mult1_un68_sum_cZ0Z4\
        );

    \I__3281\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17231\
        );

    \I__3280\ : InMux
    port map (
            O => \N__17236\,
            I => \N__17231\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__3277\ : Span4Mux_h
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__17222\,
            I => row_1_if_generate_plus_mult1_un75_sum_axbxc5_0
        );

    \I__3275\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__17216\,
            I => \ScreenBuffer_1_2Z0Z_0\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__17213\,
            I => \un3_rowlto1_cascade_\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3271\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17203\
        );

    \I__3270\ : InMux
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__17203\,
            I => \N__17197\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__17200\,
            I => \N__17194\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__17197\,
            I => \ScreenBuffer_0_2Z0Z_0\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__17194\,
            I => \ScreenBuffer_0_2Z0Z_0\
        );

    \I__3265\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17182\
        );

    \I__3263\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__17176\,
            I => \ScreenBuffer_1_1_1_sqmuxa\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__17173\,
            I => \ScreenBuffer_1_1_1_sqmuxa\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__3257\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17161\
        );

    \I__3256\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__17161\,
            I => \ScreenBuffer_0_0Z0Z_0\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__17158\,
            I => \ScreenBuffer_0_0Z0Z_0\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__17150\,
            I => \N__17146\
        );

    \I__3251\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__17143\,
            I => \ScreenBuffer_1_1Z0Z_4\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__17140\,
            I => \ScreenBuffer_1_1Z0Z_4\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__17135\,
            I => \ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_\
        );

    \I__3246\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__17129\,
            I => currentchar_1_11_ns_1_4
        );

    \I__3244\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__17123\,
            I => \ScreenBuffer_1_2_RNIUP6F2FZ0Z_4\
        );

    \I__3242\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17110\
        );

    \I__3241\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17107\
        );

    \I__3240\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17104\
        );

    \I__3239\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17101\
        );

    \I__3238\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17092\
        );

    \I__3237\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17092\
        );

    \I__3236\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17092\
        );

    \I__3235\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17092\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__17110\,
            I => \N__17087\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__17107\,
            I => \N__17087\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__17104\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__17101\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__17092\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__17087\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\
        );

    \I__3228\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17074\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__17077\,
            I => \N__17070\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__17074\,
            I => \N__17062\
        );

    \I__3225\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17057\
        );

    \I__3224\ : InMux
    port map (
            O => \N__17070\,
            I => \N__17057\
        );

    \I__3223\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17054\
        );

    \I__3222\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17045\
        );

    \I__3221\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17045\
        );

    \I__3220\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17045\
        );

    \I__3219\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17045\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__17062\,
            I => \N__17040\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__17057\,
            I => \N__17040\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__17054\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__17045\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__17040\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__17033\,
            I => \N_9_i_cascade_\
        );

    \I__3212\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__17027\,
            I => \N_13_0\
        );

    \I__3210\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__17017\
        );

    \I__3208\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17014\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__17017\,
            I => \N__17011\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__17014\,
            I => \ScreenBuffer_0_8Z0Z_0\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__17011\,
            I => \ScreenBuffer_0_8Z0Z_0\
        );

    \I__3204\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__3202\ : Odrv12
    port map (
            O => \N__17000\,
            I => \ScreenBuffer_1_0Z0Z_0\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \currentchar_1_9_ns_1_0_cascade_\
        );

    \I__3200\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3198\ : Span4Mux_h
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__16985\,
            I => \ScreenBuffer_1_1Z0Z_0\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__16982\,
            I => \currentchar_1_6_ns_1_0_cascade_\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__16979\,
            I => \N__16975\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16972\
        );

    \I__3193\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16969\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__16972\,
            I => \N__16966\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__16969\,
            I => \N__16961\
        );

    \I__3190\ : Span4Mux_v
    port map (
            O => \N__16966\,
            I => \N__16961\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__16961\,
            I => \ScreenBuffer_0_1Z0Z_0\
        );

    \I__3188\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__16955\,
            I => \N__16951\
        );

    \I__3186\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16948\
        );

    \I__3185\ : Span4Mux_v
    port map (
            O => \N__16951\,
            I => \N__16945\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__16948\,
            I => \ScreenBuffer_1_0Z0Z_4\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__16945\,
            I => \ScreenBuffer_1_0Z0Z_4\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \font_un3_pixel_28_cascade_\
        );

    \I__3181\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16933\
        );

    \I__3180\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16930\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__16933\,
            I => \un113_pixel_4_0_15__un15_beamyZ0Z_2\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__16930\,
            I => \un113_pixel_4_0_15__un15_beamyZ0Z_2\
        );

    \I__3177\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__3175\ : Span4Mux_h
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__16916\,
            I => un13_beamy
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \font_un61_pixel_cascade_\
        );

    \I__3172\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__16907\,
            I => un4_row
        );

    \I__3170\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__16901\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__16898\,
            I => \N__16895\
        );

    \I__3167\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__16892\,
            I => \N__16889\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__16889\,
            I => \N__16885\
        );

    \I__3164\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__16885\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__16882\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__3161\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16871\
        );

    \I__3160\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16871\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__16871\,
            I => charx_23
        );

    \I__3158\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__16865\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__3155\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__16856\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\
        );

    \I__3153\ : InMux
    port map (
            O => \N__16853\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__3152\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__16847\,
            I => charx_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__3150\ : InMux
    port map (
            O => \N__16844\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__3149\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__16838\,
            I => \un113_pixel_4_0_15__un18_beamylto9Z0Z_2\
        );

    \I__3147\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16830\
        );

    \I__3146\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16827\
        );

    \I__3145\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16824\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__16830\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__16827\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__16824\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__3141\ : InMux
    port map (
            O => \N__16817\,
            I => \N__16811\
        );

    \I__3140\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16811\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__16811\,
            I => charx_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__3138\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16796\
        );

    \I__3137\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16796\
        );

    \I__3136\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16796\
        );

    \I__3135\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16796\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__16796\,
            I => un1_beamx_2
        );

    \I__3133\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__16790\,
            I => charx_i_24
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__16787\,
            I => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3129\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__16778\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\
        );

    \I__3127\ : InMux
    port map (
            O => \N__16775\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3125\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__16766\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\
        );

    \I__3123\ : InMux
    port map (
            O => \N__16763\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3121\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__16754\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\
        );

    \I__3119\ : InMux
    port map (
            O => \N__16751\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__3118\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16742\
        );

    \I__3117\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16742\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__16742\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__3115\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16735\
        );

    \I__3114\ : InMux
    port map (
            O => \N__16738\,
            I => \N__16732\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__16735\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__16732\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_\
        );

    \I__3110\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16721\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__16721\,
            I => charx_if_generate_plus_mult1_un26_sum_i_5
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__3107\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__16712\,
            I => charx_if_generate_plus_mult1_un33_sum_i
        );

    \I__3105\ : InMux
    port map (
            O => \N__16709\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__3103\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16700\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__16700\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\
        );

    \I__3101\ : InMux
    port map (
            O => \N__16697\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__3100\ : InMux
    port map (
            O => \N__16694\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__3099\ : InMux
    port map (
            O => \N__16691\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__3098\ : InMux
    port map (
            O => \N__16688\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__3097\ : InMux
    port map (
            O => \N__16685\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__3096\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__16679\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\
        );

    \I__3094\ : InMux
    port map (
            O => \N__16676\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__3093\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__16670\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3090\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__16661\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0\
        );

    \I__3088\ : InMux
    port map (
            O => \N__16658\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3086\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__16649\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91\
        );

    \I__3084\ : InMux
    port map (
            O => \N__16646\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__3083\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__16640\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__3081\ : InMux
    port map (
            O => \N__16637\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__3080\ : InMux
    port map (
            O => \N__16634\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__3079\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16626\
        );

    \I__3078\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16621\
        );

    \I__3077\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16621\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__16626\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__16621\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1\
        );

    \I__3074\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__16613\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__3071\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__16604\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3068\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__16595\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__3066\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__16586\,
            I => \N__16581\
        );

    \I__3063\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16578\
        );

    \I__3062\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16574\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__16581\,
            I => \N__16569\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16569\
        );

    \I__3059\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16566\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__16574\,
            I => \voltage_3Z0Z_2\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__16569\,
            I => \voltage_3Z0Z_2\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__16566\,
            I => \voltage_3Z0Z_2\
        );

    \I__3055\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__16556\,
            I => \N__16551\
        );

    \I__3053\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16548\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__16554\,
            I => \N__16545\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__16551\,
            I => \N__16538\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16538\
        );

    \I__3049\ : InMux
    port map (
            O => \N__16545\,
            I => \N__16535\
        );

    \I__3048\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16530\
        );

    \I__3047\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16530\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__16538\,
            I => \N__16527\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__16535\,
            I => \voltage_0Z0Z_2\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__16530\,
            I => \voltage_0Z0Z_2\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__16527\,
            I => \voltage_0Z0Z_2\
        );

    \I__3042\ : InMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__16517\,
            I => un1_sclk17_7_1
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__16514\,
            I => \N__16508\
        );

    \I__3039\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16500\
        );

    \I__3038\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16500\
        );

    \I__3037\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16500\
        );

    \I__3036\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16495\
        );

    \I__3035\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16492\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__16500\,
            I => \N__16489\
        );

    \I__3033\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16486\
        );

    \I__3032\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16483\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__16495\,
            I => \N__16473\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__16492\,
            I => \N__16473\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__16489\,
            I => \N__16473\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16473\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16470\
        );

    \I__3026\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16467\
        );

    \I__3025\ : Span4Mux_h
    port map (
            O => \N__16473\,
            I => \N__16463\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__16470\,
            I => \N__16458\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__16467\,
            I => \N__16458\
        );

    \I__3022\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16455\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__16463\,
            I => un5_slaveselect
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__16458\,
            I => un5_slaveselect
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__16455\,
            I => un5_slaveselect
        );

    \I__3018\ : IoInMux
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__3016\ : Span4Mux_s2_v
    port map (
            O => \N__16442\,
            I => \N__16438\
        );

    \I__3015\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16435\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__16438\,
            I => \SDATA2_c\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__16435\,
            I => \SDATA2_c\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__16430\,
            I => \un1_sclk17_9_1_cascade_\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__16427\,
            I => \N__16420\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__16425\,
            I => \N__16414\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__16424\,
            I => \N__16411\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__16423\,
            I => \N__16403\
        );

    \I__3006\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16394\
        );

    \I__3005\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16394\
        );

    \I__3004\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16388\
        );

    \I__3003\ : InMux
    port map (
            O => \N__16411\,
            I => \N__16388\
        );

    \I__3002\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16381\
        );

    \I__3001\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16381\
        );

    \I__3000\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16381\
        );

    \I__2999\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16378\
        );

    \I__2998\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16375\
        );

    \I__2997\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16366\
        );

    \I__2996\ : InMux
    port map (
            O => \N__16402\,
            I => \N__16366\
        );

    \I__2995\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16366\
        );

    \I__2994\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16366\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__16399\,
            I => \N__16363\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__16394\,
            I => \N__16357\
        );

    \I__2991\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16354\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16351\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__16381\,
            I => \N__16348\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__16378\,
            I => \N__16341\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16336\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__16366\,
            I => \N__16336\
        );

    \I__2985\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16333\
        );

    \I__2984\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16328\
        );

    \I__2983\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16328\
        );

    \I__2982\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16325\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__16357\,
            I => \N__16316\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__16354\,
            I => \N__16316\
        );

    \I__2979\ : Span4Mux_s3_v
    port map (
            O => \N__16351\,
            I => \N__16316\
        );

    \I__2978\ : Span4Mux_s3_v
    port map (
            O => \N__16348\,
            I => \N__16316\
        );

    \I__2977\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16311\
        );

    \I__2976\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16311\
        );

    \I__2975\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16306\
        );

    \I__2974\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16306\
        );

    \I__2973\ : Span4Mux_v
    port map (
            O => \N__16341\,
            I => \N__16297\
        );

    \I__2972\ : Span4Mux_s3_v
    port map (
            O => \N__16336\,
            I => \N__16297\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__16333\,
            I => \N__16297\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__16328\,
            I => \N__16297\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__16325\,
            I => \counterZ0Z_3\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__16316\,
            I => \counterZ0Z_3\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__16311\,
            I => \counterZ0Z_3\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__16306\,
            I => \counterZ0Z_3\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__16297\,
            I => \counterZ0Z_3\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__16286\,
            I => \N__16279\
        );

    \I__2963\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16270\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__16284\,
            I => \N__16262\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__16283\,
            I => \N__16252\
        );

    \I__2960\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16234\
        );

    \I__2959\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16234\
        );

    \I__2958\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16234\
        );

    \I__2957\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16231\
        );

    \I__2956\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16224\
        );

    \I__2955\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16224\
        );

    \I__2954\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16224\
        );

    \I__2953\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16218\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16209\
        );

    \I__2951\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16204\
        );

    \I__2950\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16204\
        );

    \I__2949\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16201\
        );

    \I__2948\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16198\
        );

    \I__2947\ : InMux
    port map (
            O => \N__16265\,
            I => \N__16189\
        );

    \I__2946\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16189\
        );

    \I__2945\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16189\
        );

    \I__2944\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16189\
        );

    \I__2943\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16182\
        );

    \I__2942\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16182\
        );

    \I__2941\ : InMux
    port map (
            O => \N__16257\,
            I => \N__16182\
        );

    \I__2940\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16174\
        );

    \I__2939\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16174\
        );

    \I__2938\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16174\
        );

    \I__2937\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16167\
        );

    \I__2936\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16167\
        );

    \I__2935\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16167\
        );

    \I__2934\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16160\
        );

    \I__2933\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16160\
        );

    \I__2932\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16160\
        );

    \I__2931\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16157\
        );

    \I__2930\ : InMux
    port map (
            O => \N__16244\,
            I => \N__16154\
        );

    \I__2929\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16151\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__16242\,
            I => \N__16147\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__16241\,
            I => \N__16144\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__16234\,
            I => \N__16141\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__16231\,
            I => \N__16138\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__16224\,
            I => \N__16135\
        );

    \I__2923\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16128\
        );

    \I__2922\ : InMux
    port map (
            O => \N__16222\,
            I => \N__16128\
        );

    \I__2921\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16128\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16125\
        );

    \I__2919\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16118\
        );

    \I__2918\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16118\
        );

    \I__2917\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16118\
        );

    \I__2916\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16113\
        );

    \I__2915\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16113\
        );

    \I__2914\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16110\
        );

    \I__2913\ : Span4Mux_s3_h
    port map (
            O => \N__16209\,
            I => \N__16106\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__16204\,
            I => \N__16101\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__16201\,
            I => \N__16101\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__16198\,
            I => \N__16098\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__16189\,
            I => \N__16093\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16093\
        );

    \I__2907\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16090\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16085\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16085\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__16160\,
            I => \N__16080\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16080\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__16154\,
            I => \N__16075\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__16151\,
            I => \N__16075\
        );

    \I__2900\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16072\
        );

    \I__2899\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16069\
        );

    \I__2898\ : InMux
    port map (
            O => \N__16144\,
            I => \N__16066\
        );

    \I__2897\ : Span4Mux_s3_h
    port map (
            O => \N__16141\,
            I => \N__16061\
        );

    \I__2896\ : Span4Mux_s3_h
    port map (
            O => \N__16138\,
            I => \N__16061\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__16135\,
            I => \N__16054\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16054\
        );

    \I__2893\ : Span4Mux_s2_h
    port map (
            O => \N__16125\,
            I => \N__16054\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__16118\,
            I => \N__16051\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__16113\,
            I => \N__16048\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__16110\,
            I => \N__16045\
        );

    \I__2889\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16042\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__16106\,
            I => \N__16037\
        );

    \I__2887\ : Span4Mux_s3_h
    port map (
            O => \N__16101\,
            I => \N__16037\
        );

    \I__2886\ : Span4Mux_h
    port map (
            O => \N__16098\,
            I => \N__16026\
        );

    \I__2885\ : Span4Mux_s3_h
    port map (
            O => \N__16093\,
            I => \N__16026\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__16090\,
            I => \N__16026\
        );

    \I__2883\ : Span4Mux_s3_h
    port map (
            O => \N__16085\,
            I => \N__16026\
        );

    \I__2882\ : Span4Mux_h
    port map (
            O => \N__16080\,
            I => \N__16026\
        );

    \I__2881\ : Span12Mux_s3_h
    port map (
            O => \N__16075\,
            I => \N__16023\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__16072\,
            I => \counterZ0Z_0\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__16069\,
            I => \counterZ0Z_0\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__16066\,
            I => \counterZ0Z_0\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__16061\,
            I => \counterZ0Z_0\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__16054\,
            I => \counterZ0Z_0\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__16051\,
            I => \counterZ0Z_0\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__16048\,
            I => \counterZ0Z_0\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__16045\,
            I => \counterZ0Z_0\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__16042\,
            I => \counterZ0Z_0\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__16037\,
            I => \counterZ0Z_0\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__16026\,
            I => \counterZ0Z_0\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__16023\,
            I => \counterZ0Z_0\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__15998\,
            I => \N__15985\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__15997\,
            I => \N__15982\
        );

    \I__2866\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15971\
        );

    \I__2865\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15964\
        );

    \I__2864\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15964\
        );

    \I__2863\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15964\
        );

    \I__2862\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15959\
        );

    \I__2861\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15959\
        );

    \I__2860\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15952\
        );

    \I__2859\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15952\
        );

    \I__2858\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15952\
        );

    \I__2857\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15947\
        );

    \I__2856\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15947\
        );

    \I__2855\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15938\
        );

    \I__2854\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15938\
        );

    \I__2853\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15938\
        );

    \I__2852\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15938\
        );

    \I__2851\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15930\
        );

    \I__2850\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15930\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__15975\,
            I => \N__15927\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__15974\,
            I => \N__15924\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15918\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__15964\,
            I => \N__15918\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N__15913\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15913\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15910\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__15938\,
            I => \N__15907\
        );

    \I__2841\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15902\
        );

    \I__2840\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15902\
        );

    \I__2839\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15899\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15896\
        );

    \I__2837\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15893\
        );

    \I__2836\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15890\
        );

    \I__2835\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15887\
        );

    \I__2834\ : Span4Mux_s3_v
    port map (
            O => \N__15918\,
            I => \N__15876\
        );

    \I__2833\ : Span4Mux_s3_v
    port map (
            O => \N__15913\,
            I => \N__15876\
        );

    \I__2832\ : Span4Mux_s3_v
    port map (
            O => \N__15910\,
            I => \N__15876\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__15907\,
            I => \N__15876\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__15902\,
            I => \N__15876\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__15899\,
            I => \counterZ0Z_2\
        );

    \I__2828\ : Odrv12
    port map (
            O => \N__15896\,
            I => \counterZ0Z_2\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__15893\,
            I => \counterZ0Z_2\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__15890\,
            I => \counterZ0Z_2\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__15887\,
            I => \counterZ0Z_2\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__15876\,
            I => \counterZ0Z_2\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \N__15858\
        );

    \I__2822\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15851\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__15861\,
            I => \N__15848\
        );

    \I__2820\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15845\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__15857\,
            I => \N__15842\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15838\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15833\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__15854\,
            I => \N__15829\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__15851\,
            I => \N__15826\
        );

    \I__2814\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15823\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__15845\,
            I => \N__15807\
        );

    \I__2812\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15804\
        );

    \I__2811\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15797\
        );

    \I__2810\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15797\
        );

    \I__2809\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15797\
        );

    \I__2808\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15794\
        );

    \I__2807\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15787\
        );

    \I__2806\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15787\
        );

    \I__2805\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15787\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__15826\,
            I => \N__15782\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__15823\,
            I => \N__15782\
        );

    \I__2802\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15773\
        );

    \I__2801\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15773\
        );

    \I__2800\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15773\
        );

    \I__2799\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15773\
        );

    \I__2798\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15770\
        );

    \I__2797\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15767\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \N__15760\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15757\
        );

    \I__2794\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15751\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__15813\,
            I => \N__15746\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__15812\,
            I => \N__15743\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__15811\,
            I => \N__15736\
        );

    \I__2790\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15730\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__15807\,
            I => \N__15723\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__15804\,
            I => \N__15723\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__15797\,
            I => \N__15723\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__15794\,
            I => \N__15715\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15708\
        );

    \I__2784\ : Span4Mux_s3_v
    port map (
            O => \N__15782\,
            I => \N__15708\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15708\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15703\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__15767\,
            I => \N__15703\
        );

    \I__2780\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15694\
        );

    \I__2779\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15694\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15764\,
            I => \N__15694\
        );

    \I__2777\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15694\
        );

    \I__2776\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15689\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15689\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__15756\,
            I => \N__15685\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__15755\,
            I => \N__15681\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__15754\,
            I => \N__15678\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15675\
        );

    \I__2770\ : InMux
    port map (
            O => \N__15750\,
            I => \N__15672\
        );

    \I__2769\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15665\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15665\
        );

    \I__2767\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15665\
        );

    \I__2766\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15659\
        );

    \I__2765\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15659\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15650\
        );

    \I__2763\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15650\
        );

    \I__2762\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15650\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15650\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15647\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__15733\,
            I => \N__15644\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15636\
        );

    \I__2757\ : Span4Mux_s3_v
    port map (
            O => \N__15723\,
            I => \N__15636\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15631\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15631\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15624\
        );

    \I__2753\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15624\
        );

    \I__2752\ : InMux
    port map (
            O => \N__15718\,
            I => \N__15624\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__15715\,
            I => \N__15615\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__15708\,
            I => \N__15615\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__15703\,
            I => \N__15615\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__15694\,
            I => \N__15615\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15612\
        );

    \I__2746\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15607\
        );

    \I__2745\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15607\
        );

    \I__2744\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15604\
        );

    \I__2743\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15601\
        );

    \I__2742\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15598\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__15675\,
            I => \N__15591\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__15672\,
            I => \N__15591\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15591\
        );

    \I__2738\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15588\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__15659\,
            I => \N__15583\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__15650\,
            I => \N__15583\
        );

    \I__2735\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15572\
        );

    \I__2734\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15572\
        );

    \I__2733\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15572\
        );

    \I__2732\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15572\
        );

    \I__2731\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15572\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__15636\,
            I => \N__15567\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__15631\,
            I => \N__15567\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__15624\,
            I => \N__15562\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__15615\,
            I => \N__15562\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__15612\,
            I => \counterZ0Z_1\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__15607\,
            I => \counterZ0Z_1\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__15604\,
            I => \counterZ0Z_1\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__15601\,
            I => \counterZ0Z_1\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__15598\,
            I => \counterZ0Z_1\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__15591\,
            I => \counterZ0Z_1\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__15588\,
            I => \counterZ0Z_1\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__15583\,
            I => \counterZ0Z_1\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__15572\,
            I => \counterZ0Z_1\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__15567\,
            I => \counterZ0Z_1\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__15562\,
            I => \counterZ0Z_1\
        );

    \I__2715\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15536\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__15536\,
            I => un1_sclk17_4_1
        );

    \I__2713\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15529\
        );

    \I__2712\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15526\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__15529\,
            I => \N_1505\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__15526\,
            I => \N_1505\
        );

    \I__2709\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15516\
        );

    \I__2708\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15513\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__15519\,
            I => \N__15509\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__15516\,
            I => \N__15506\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__15513\,
            I => \N__15503\
        );

    \I__2704\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15498\
        );

    \I__2703\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15498\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__15506\,
            I => \N__15495\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__15503\,
            I => \N__15492\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__15498\,
            I => \N_1509\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__15495\,
            I => \N_1509\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__15492\,
            I => \N_1509\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__15485\,
            I => \N__15482\
        );

    \I__2696\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__15476\,
            I => \un42_cry_2_c_RNOZ0\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \un1_sclk17_6_1_cascade_\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__15470\,
            I => \un1_sclk17_3_1_cascade_\
        );

    \I__2691\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__2689\ : Odrv12
    port map (
            O => \N__15461\,
            I => \ScreenBuffer_0_0_1_sqmuxa_0\
        );

    \I__2688\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15454\
        );

    \I__2687\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__15454\,
            I => \slaveselect_RNILOQCZ0Z2\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__15451\,
            I => \slaveselect_RNILOQCZ0Z2\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__15446\,
            I => \un1_sclk17_8_0_0_cascade_\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__2682\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__15437\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3\
        );

    \I__2680\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__15431\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5
        );

    \I__2678\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__15425\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\
        );

    \I__2676\ : InMux
    port map (
            O => \N__15422\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4
        );

    \I__2675\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15413\
        );

    \I__2674\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15413\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__15413\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__15410\,
            I => \N__15406\
        );

    \I__2671\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15398\
        );

    \I__2670\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15398\
        );

    \I__2669\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15398\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__15398\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\
        );

    \I__2667\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__15392\,
            I => \N__15386\
        );

    \I__2665\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15381\
        );

    \I__2664\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15381\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__15389\,
            I => \N__15376\
        );

    \I__2662\ : Span4Mux_h
    port map (
            O => \N__15386\,
            I => \N__15372\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15369\
        );

    \I__2660\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15366\
        );

    \I__2659\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15363\
        );

    \I__2658\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15358\
        );

    \I__2657\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15358\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__15372\,
            I => \N__15353\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__15369\,
            I => \N__15353\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__15366\,
            I => \voltage_2Z0Z_0\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__15363\,
            I => \voltage_2Z0Z_0\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__15358\,
            I => \voltage_2Z0Z_0\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__15353\,
            I => \voltage_2Z0Z_0\
        );

    \I__2650\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15340\
        );

    \I__2649\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15336\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15333\
        );

    \I__2647\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15330\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__15336\,
            I => \N__15325\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__15333\,
            I => \N__15322\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__15330\,
            I => \N__15319\
        );

    \I__2643\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15314\
        );

    \I__2642\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15314\
        );

    \I__2641\ : Odrv12
    port map (
            O => \N__15325\,
            I => \voltage_1Z0Z_0\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__15322\,
            I => \voltage_1Z0Z_0\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__15319\,
            I => \voltage_1Z0Z_0\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__15314\,
            I => \voltage_1Z0Z_0\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__2636\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15298\
        );

    \I__2635\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15295\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__15298\,
            I => \N__15290\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__15295\,
            I => \N__15287\
        );

    \I__2632\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15283\
        );

    \I__2631\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15280\
        );

    \I__2630\ : Span4Mux_v
    port map (
            O => \N__15290\,
            I => \N__15275\
        );

    \I__2629\ : Span4Mux_s1_h
    port map (
            O => \N__15287\,
            I => \N__15275\
        );

    \I__2628\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15272\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__15283\,
            I => \voltage_2Z0Z_2\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__15280\,
            I => \voltage_2Z0Z_2\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__15275\,
            I => \voltage_2Z0Z_2\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__15272\,
            I => \voltage_2Z0Z_2\
        );

    \I__2623\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15258\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__15262\,
            I => \N__15255\
        );

    \I__2621\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15252\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__15258\,
            I => \N__15249\
        );

    \I__2619\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15246\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__15252\,
            I => \N__15242\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__15249\,
            I => \N__15239\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__15246\,
            I => \N__15236\
        );

    \I__2615\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15233\
        );

    \I__2614\ : Odrv12
    port map (
            O => \N__15242\,
            I => \voltage_1Z0Z_2\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__15239\,
            I => \voltage_1Z0Z_2\
        );

    \I__2612\ : Odrv12
    port map (
            O => \N__15236\,
            I => \voltage_1Z0Z_2\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__15233\,
            I => \voltage_1Z0Z_2\
        );

    \I__2610\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15220\
        );

    \I__2609\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15216\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__15220\,
            I => \N__15213\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15210\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__15216\,
            I => \N__15206\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__15213\,
            I => \N__15202\
        );

    \I__2604\ : InMux
    port map (
            O => \N__15210\,
            I => \N__15197\
        );

    \I__2603\ : InMux
    port map (
            O => \N__15209\,
            I => \N__15197\
        );

    \I__2602\ : Span4Mux_v
    port map (
            O => \N__15206\,
            I => \N__15194\
        );

    \I__2601\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15191\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__15202\,
            I => \N__15188\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__15197\,
            I => \N__15185\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__15194\,
            I => \voltage_2Z0Z_3\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__15191\,
            I => \voltage_2Z0Z_3\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__15188\,
            I => \voltage_2Z0Z_3\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__15185\,
            I => \voltage_2Z0Z_3\
        );

    \I__2594\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15172\
        );

    \I__2593\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15169\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__15172\,
            I => \N__15164\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__15169\,
            I => \N__15164\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__15164\,
            I => \N__15159\
        );

    \I__2589\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15156\
        );

    \I__2588\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15153\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__15159\,
            I => \voltage_1Z0Z_3\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__15156\,
            I => \voltage_1Z0Z_3\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__15153\,
            I => \voltage_1Z0Z_3\
        );

    \I__2584\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15143\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__15143\,
            I => \N__15139\
        );

    \I__2582\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15136\
        );

    \I__2581\ : Span4Mux_s2_h
    port map (
            O => \N__15139\,
            I => \N__15130\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__15136\,
            I => \N__15130\
        );

    \I__2579\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15124\
        );

    \I__2578\ : Span4Mux_v
    port map (
            O => \N__15130\,
            I => \N__15121\
        );

    \I__2577\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15116\
        );

    \I__2576\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15116\
        );

    \I__2575\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15113\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__15124\,
            I => \voltage_2Z0Z_1\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__15121\,
            I => \voltage_2Z0Z_1\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__15116\,
            I => \voltage_2Z0Z_1\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__15113\,
            I => \voltage_2Z0Z_1\
        );

    \I__2570\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N__15096\
        );

    \I__2568\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15093\
        );

    \I__2567\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15090\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__15096\,
            I => \N__15087\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__15093\,
            I => \N__15083\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__15090\,
            I => \N__15078\
        );

    \I__2563\ : Span4Mux_s2_h
    port map (
            O => \N__15087\,
            I => \N__15078\
        );

    \I__2562\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15075\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__15083\,
            I => \voltage_1Z0Z_1\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__15078\,
            I => \voltage_1Z0Z_1\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__15075\,
            I => \voltage_1Z0Z_1\
        );

    \I__2558\ : CEMux
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__15065\,
            I => \N__15062\
        );

    \I__2556\ : Span4Mux_h
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__2555\ : Odrv4
    port map (
            O => \N__15059\,
            I => \un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0\
        );

    \I__2554\ : InMux
    port map (
            O => \N__15056\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1
        );

    \I__2553\ : InMux
    port map (
            O => \N__15053\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2
        );

    \I__2552\ : InMux
    port map (
            O => \N__15050\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3
        );

    \I__2551\ : InMux
    port map (
            O => \N__15047\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__2549\ : InMux
    port map (
            O => \N__15041\,
            I => \N__15038\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__15038\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_i
        );

    \I__2547\ : InMux
    port map (
            O => \N__15035\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1
        );

    \I__2546\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__15029\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3\
        );

    \I__2544\ : InMux
    port map (
            O => \N__15026\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2
        );

    \I__2543\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__15017\,
            I => un13_beamy_0
        );

    \I__2540\ : InMux
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__15008\,
            I => chessboardpixel_un174_pixel
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__15005\,
            I => \un4_row_cascade_\
        );

    \I__2536\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__14999\,
            I => \N__14995\
        );

    \I__2534\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14992\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__14995\,
            I => \N__14984\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14984\
        );

    \I__2531\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14980\
        );

    \I__2530\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14977\
        );

    \I__2529\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14974\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__14984\,
            I => \N__14969\
        );

    \I__2527\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14966\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__14980\,
            I => \N__14963\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__14977\,
            I => \N__14958\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14958\
        );

    \I__2523\ : InMux
    port map (
            O => \N__14973\,
            I => \N__14955\
        );

    \I__2522\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14952\
        );

    \I__2521\ : Sp12to4
    port map (
            O => \N__14969\,
            I => \N__14947\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14947\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__14963\,
            I => \N__14942\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__14958\,
            I => \N__14942\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14939\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__14952\,
            I => \beamYZ0Z_9\
        );

    \I__2515\ : Odrv12
    port map (
            O => \N__14947\,
            I => \beamYZ0Z_9\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__14942\,
            I => \beamYZ0Z_9\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__14939\,
            I => \beamYZ0Z_9\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__14930\,
            I => \N__14926\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \N__14922\
        );

    \I__2510\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14917\
        );

    \I__2509\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14914\
        );

    \I__2508\ : InMux
    port map (
            O => \N__14922\,
            I => \N__14911\
        );

    \I__2507\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14908\
        );

    \I__2506\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14905\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__14917\,
            I => \N__14898\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__14914\,
            I => \N__14898\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__14911\,
            I => \N__14898\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__14908\,
            I => \N__14893\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__14905\,
            I => \N__14893\
        );

    \I__2500\ : Span4Mux_v
    port map (
            O => \N__14898\,
            I => \N__14884\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__14893\,
            I => \N__14884\
        );

    \I__2498\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14881\
        );

    \I__2497\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14878\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__14890\,
            I => \N__14874\
        );

    \I__2495\ : InMux
    port map (
            O => \N__14889\,
            I => \N__14871\
        );

    \I__2494\ : Sp12to4
    port map (
            O => \N__14884\,
            I => \N__14866\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__14881\,
            I => \N__14866\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14863\
        );

    \I__2491\ : InMux
    port map (
            O => \N__14877\,
            I => \N__14860\
        );

    \I__2490\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14857\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__14871\,
            I => \beamYZ0Z_8\
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__14866\,
            I => \beamYZ0Z_8\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__14863\,
            I => \beamYZ0Z_8\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__14860\,
            I => \beamYZ0Z_8\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__14857\,
            I => \beamYZ0Z_8\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__14846\,
            I => \N__14842\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__14845\,
            I => \N__14839\
        );

    \I__2482\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14834\
        );

    \I__2481\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14831\
        );

    \I__2480\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14828\
        );

    \I__2479\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14825\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__14834\,
            I => \N__14821\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14818\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14813\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14813\
        );

    \I__2474\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14806\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__14821\,
            I => \N__14803\
        );

    \I__2472\ : Span4Mux_h
    port map (
            O => \N__14818\,
            I => \N__14800\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__14813\,
            I => \N__14797\
        );

    \I__2470\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14794\
        );

    \I__2469\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14791\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14786\
        );

    \I__2467\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14777\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__14806\,
            I => \N__14774\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__14803\,
            I => \N__14771\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__14800\,
            I => \N__14768\
        );

    \I__2463\ : Sp12to4
    port map (
            O => \N__14797\,
            I => \N__14761\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14761\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__14791\,
            I => \N__14761\
        );

    \I__2460\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14756\
        );

    \I__2459\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14756\
        );

    \I__2458\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14751\
        );

    \I__2457\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14751\
        );

    \I__2456\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14746\
        );

    \I__2455\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14746\
        );

    \I__2454\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14739\
        );

    \I__2453\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14739\
        );

    \I__2452\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14739\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__14777\,
            I => \beamYZ0Z_7\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__14774\,
            I => \beamYZ0Z_7\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__14771\,
            I => \beamYZ0Z_7\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__14768\,
            I => \beamYZ0Z_7\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__14761\,
            I => \beamYZ0Z_7\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__14756\,
            I => \beamYZ0Z_7\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__14751\,
            I => \beamYZ0Z_7\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__14746\,
            I => \beamYZ0Z_7\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__14739\,
            I => \beamYZ0Z_7\
        );

    \I__2442\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__14717\,
            I => un4_beamylt8_0
        );

    \I__2440\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14711\,
            I => un4_beamy_0
        );

    \I__2438\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__14705\,
            I => \un113_pixel_4_0_15__un8_beamylto9Z0Z_1\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14697\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__14701\,
            I => \N__14691\
        );

    \I__2434\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14684\
        );

    \I__2433\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14681\
        );

    \I__2432\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14678\
        );

    \I__2431\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14675\
        );

    \I__2430\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14672\
        );

    \I__2429\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14669\
        );

    \I__2428\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14662\
        );

    \I__2427\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14662\
        );

    \I__2426\ : InMux
    port map (
            O => \N__14688\,
            I => \N__14662\
        );

    \I__2425\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14654\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14651\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14648\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__14678\,
            I => \N__14645\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__14675\,
            I => \N__14640\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__14672\,
            I => \N__14640\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__14669\,
            I => \N__14637\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14634\
        );

    \I__2417\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14631\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__14660\,
            I => \N__14627\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__14659\,
            I => \N__14624\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__14658\,
            I => \N__14618\
        );

    \I__2413\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14614\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__14654\,
            I => \N__14611\
        );

    \I__2411\ : Span12Mux_s5_v
    port map (
            O => \N__14651\,
            I => \N__14606\
        );

    \I__2410\ : Span12Mux_s10_v
    port map (
            O => \N__14648\,
            I => \N__14606\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__14645\,
            I => \N__14601\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__14640\,
            I => \N__14601\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__14637\,
            I => \N__14596\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__14634\,
            I => \N__14596\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__14631\,
            I => \N__14593\
        );

    \I__2404\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14588\
        );

    \I__2403\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14588\
        );

    \I__2402\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14585\
        );

    \I__2401\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14580\
        );

    \I__2400\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14580\
        );

    \I__2399\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14573\
        );

    \I__2398\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14573\
        );

    \I__2397\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14573\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__14614\,
            I => \beamYZ0Z_4\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__14611\,
            I => \beamYZ0Z_4\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__14606\,
            I => \beamYZ0Z_4\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__14601\,
            I => \beamYZ0Z_4\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__14596\,
            I => \beamYZ0Z_4\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__14593\,
            I => \beamYZ0Z_4\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__14588\,
            I => \beamYZ0Z_4\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__14585\,
            I => \beamYZ0Z_4\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__14580\,
            I => \beamYZ0Z_4\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__14573\,
            I => \beamYZ0Z_4\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__2385\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__14543\,
            I => un8_beamy
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__14540\,
            I => \N__14537\
        );

    \I__2381\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14534\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__14534\,
            I => \N_6_i\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__14531\,
            I => \N_6_i_cascade_\
        );

    \I__2378\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__14522\,
            I => \N__14514\
        );

    \I__2375\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14511\
        );

    \I__2374\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14502\
        );

    \I__2373\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14502\
        );

    \I__2372\ : InMux
    port map (
            O => \N__14518\,
            I => \N__14502\
        );

    \I__2371\ : InMux
    port map (
            O => \N__14517\,
            I => \N__14502\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__14514\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__14511\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__14502\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\
        );

    \I__2367\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14491\
        );

    \I__2366\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14488\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14482\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14482\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__14487\,
            I => \N__14473\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__14482\,
            I => \N__14466\
        );

    \I__2361\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14459\
        );

    \I__2360\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14459\
        );

    \I__2359\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14459\
        );

    \I__2358\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14454\
        );

    \I__2357\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14454\
        );

    \I__2356\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14451\
        );

    \I__2355\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14442\
        );

    \I__2354\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14442\
        );

    \I__2353\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14442\
        );

    \I__2352\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14442\
        );

    \I__2351\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14437\
        );

    \I__2350\ : Sp12to4
    port map (
            O => \N__14466\,
            I => \N__14430\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14430\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14430\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__14451\,
            I => \N__14425\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14425\
        );

    \I__2345\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14422\
        );

    \I__2344\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14414\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14411\
        );

    \I__2342\ : Span12Mux_s11_h
    port map (
            O => \N__14430\,
            I => \N__14408\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__14425\,
            I => \N__14403\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__14422\,
            I => \N__14403\
        );

    \I__2339\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14400\
        );

    \I__2338\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14395\
        );

    \I__2337\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14395\
        );

    \I__2336\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14392\
        );

    \I__2335\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14389\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__14414\,
            I => \beamYZ0Z_3\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__14411\,
            I => \beamYZ0Z_3\
        );

    \I__2332\ : Odrv12
    port map (
            O => \N__14408\,
            I => \beamYZ0Z_3\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__14403\,
            I => \beamYZ0Z_3\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__14400\,
            I => \beamYZ0Z_3\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__14395\,
            I => \beamYZ0Z_3\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__14392\,
            I => \beamYZ0Z_3\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__14389\,
            I => \beamYZ0Z_3\
        );

    \I__2326\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14367\
        );

    \I__2325\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14364\
        );

    \I__2324\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14361\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__14367\,
            I => un4_beamylt6
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__14364\,
            I => un4_beamylt6
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__14361\,
            I => un4_beamylt6
        );

    \I__2320\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14351\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__14351\,
            I => \N__14348\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__14348\,
            I => if_m1_ns
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \if_m2_2_cascade_\
        );

    \I__2316\ : InMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__14339\,
            I => row_1_if_generate_plus_mult1_un82_sum_axbxc5_0
        );

    \I__2314\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14330\
        );

    \I__2313\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14330\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__14330\,
            I => un18_beamylt4
        );

    \I__2311\ : InMux
    port map (
            O => \N__14327\,
            I => \N__14324\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__14324\,
            I => \un113_pixel_4_0_15__un4_rowZ0Z_2\
        );

    \I__2309\ : InMux
    port map (
            O => \N__14321\,
            I => \N__14318\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__14318\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__2306\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14307\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__14311\,
            I => \N__14304\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__14310\,
            I => \N__14300\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__14307\,
            I => \N__14294\
        );

    \I__2302\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14289\
        );

    \I__2301\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14289\
        );

    \I__2300\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14284\
        );

    \I__2299\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14284\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__14298\,
            I => \N__14281\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__14297\,
            I => \N__14278\
        );

    \I__2296\ : Span4Mux_h
    port map (
            O => \N__14294\,
            I => \N__14273\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__14289\,
            I => \N__14273\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14270\
        );

    \I__2293\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14265\
        );

    \I__2292\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14265\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__14273\,
            I => \N__14260\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__14270\,
            I => \N__14260\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__14265\,
            I => \N__14257\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__14260\,
            I => \N__14254\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__14257\,
            I => \r_N_6\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__14254\,
            I => \r_N_6\
        );

    \I__2285\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__14246\,
            I => \un113_pixel_4_0_15__un3_beamxZ0Z_7\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__14243\,
            I => \un1_beamxlt10_0_cascade_\
        );

    \I__2282\ : IoInMux
    port map (
            O => \N__14240\,
            I => \N__14237\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__2280\ : IoSpan4Mux
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2279\ : Span4Mux_s3_v
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__14228\,
            I => \HSync_c\
        );

    \I__2277\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__14222\,
            I => un18_beamylt10_0
        );

    \I__2275\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14216\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__14216\,
            I => if_generate_plus_mult1_un82_sum_axbxc5_0_x1
        );

    \I__2273\ : InMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__14210\,
            I => if_generate_plus_mult1_un82_sum_axbxc5_0_x0
        );

    \I__2271\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14199\
        );

    \I__2269\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14196\
        );

    \I__2268\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14193\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__14199\,
            I => un1_beamy_4
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__14196\,
            I => un1_beamy_4
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__14193\,
            I => un1_beamy_4
        );

    \I__2264\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14181\
        );

    \I__2263\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14176\
        );

    \I__2262\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14176\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__14181\,
            I => \N__14171\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14171\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__14171\,
            I => \N__14168\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__14168\,
            I => row_1_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__14165\,
            I => \N__14162\
        );

    \I__2256\ : InMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__14159\,
            I => \un113_pixel_4_0_15__un4_rowZ0Z_5\
        );

    \I__2254\ : InMux
    port map (
            O => \N__14156\,
            I => \N__14153\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__14153\,
            I => \un113_pixel_4_0_15__un5_beamx_2Z0Z_0\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__14150\,
            I => \un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14147\,
            I => \N__14139\
        );

    \I__2250\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14139\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14136\
        );

    \I__2248\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14133\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__14139\,
            I => \N__14126\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__14136\,
            I => \N__14126\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__14133\,
            I => \N__14126\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__14126\,
            I => \N__14122\
        );

    \I__2243\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14119\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__14122\,
            I => \N__14116\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__14119\,
            I => un5_beamx_0
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__14116\,
            I => un5_beamx_0
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \un5_beamx_0_cascade_\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__14108\,
            I => \un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_\
        );

    \I__2237\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__14102\,
            I => un13_beamylt6_0
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__14099\,
            I => \un13_beamylt6_0_cascade_\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__14096\,
            I => \N__14093\
        );

    \I__2233\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__14090\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2\
        );

    \I__2231\ : InMux
    port map (
            O => \N__14087\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__2230\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14081\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__14081\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__2228\ : InMux
    port map (
            O => \N__14078\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__2227\ : InMux
    port map (
            O => \N__14075\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__2226\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14067\
        );

    \I__2225\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14062\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14062\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__14067\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__14062\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14051\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14051\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__14051\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__2217\ : InMux
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__14042\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__14039\,
            I => \N__14029\
        );

    \I__2214\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14025\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14037\,
            I => \N__14022\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__14036\,
            I => \N__14017\
        );

    \I__2211\ : InMux
    port map (
            O => \N__14035\,
            I => \N__14012\
        );

    \I__2210\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14012\
        );

    \I__2209\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14009\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14004\
        );

    \I__2207\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14004\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__14028\,
            I => \N__13998\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__14025\,
            I => \N__13993\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__14022\,
            I => \N__13990\
        );

    \I__2203\ : InMux
    port map (
            O => \N__14021\,
            I => \N__13983\
        );

    \I__2202\ : InMux
    port map (
            O => \N__14020\,
            I => \N__13983\
        );

    \I__2201\ : InMux
    port map (
            O => \N__14017\,
            I => \N__13983\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__14012\,
            I => \N__13976\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__13976\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__14004\,
            I => \N__13976\
        );

    \I__2197\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13971\
        );

    \I__2196\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13971\
        );

    \I__2195\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13966\
        );

    \I__2194\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13966\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__13997\,
            I => \N__13962\
        );

    \I__2192\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13959\
        );

    \I__2191\ : Span4Mux_h
    port map (
            O => \N__13993\,
            I => \N__13952\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__13990\,
            I => \N__13952\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13952\
        );

    \I__2188\ : Span12Mux_s11_h
    port map (
            O => \N__13976\,
            I => \N__13947\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__13971\,
            I => \N__13947\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13944\
        );

    \I__2185\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13939\
        );

    \I__2184\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13939\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__13959\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__13952\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2181\ : Odrv12
    port map (
            O => \N__13947\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__13944\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__13939\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__2177\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13918\
        );

    \I__2176\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13915\
        );

    \I__2175\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13912\
        );

    \I__2174\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13907\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13907\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__13918\,
            I => \counterZ0Z_9\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__13915\,
            I => \counterZ0Z_9\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__13912\,
            I => \counterZ0Z_9\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__13907\,
            I => \counterZ0Z_9\
        );

    \I__2168\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13892\
        );

    \I__2167\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13889\
        );

    \I__2166\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13884\
        );

    \I__2165\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13884\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__13892\,
            I => \counterZ0Z_7\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__13889\,
            I => \counterZ0Z_7\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__13884\,
            I => \counterZ0Z_7\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__13877\,
            I => \un1_counter_1lto9_2_cascade_\
        );

    \I__2160\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__13871\,
            I => un10_slaveselectlt4
        );

    \I__2158\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__13865\,
            I => \N__13856\
        );

    \I__2156\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13852\
        );

    \I__2155\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13849\
        );

    \I__2154\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13846\
        );

    \I__2153\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13843\
        );

    \I__2152\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13840\
        );

    \I__2151\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13837\
        );

    \I__2150\ : Span4Mux_s3_h
    port map (
            O => \N__13856\,
            I => \N__13834\
        );

    \I__2149\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13831\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__13852\,
            I => \N__13826\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__13849\,
            I => \N__13826\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__13846\,
            I => \counterZ0Z_4\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13843\,
            I => \counterZ0Z_4\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__13840\,
            I => \counterZ0Z_4\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__13837\,
            I => \counterZ0Z_4\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__13834\,
            I => \counterZ0Z_4\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__13831\,
            I => \counterZ0Z_4\
        );

    \I__2140\ : Odrv12
    port map (
            O => \N__13826\,
            I => \counterZ0Z_4\
        );

    \I__2139\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13807\
        );

    \I__2138\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__13807\,
            I => un1_counter_1lt9
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__13804\,
            I => un1_counter_1lt9
        );

    \I__2135\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13796\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__13796\,
            I => \N__13790\
        );

    \I__2133\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13787\
        );

    \I__2132\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13784\
        );

    \I__2131\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13781\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__13790\,
            I => \counterZ0Z_6\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__13787\,
            I => \counterZ0Z_6\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__13784\,
            I => \counterZ0Z_6\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__13781\,
            I => \counterZ0Z_6\
        );

    \I__2126\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13768\
        );

    \I__2125\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13760\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__13768\,
            I => \N__13757\
        );

    \I__2123\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13754\
        );

    \I__2122\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13751\
        );

    \I__2121\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13748\
        );

    \I__2120\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13745\
        );

    \I__2119\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13742\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__13760\,
            I => \N__13739\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__13757\,
            I => \counterZ0Z_5\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__13754\,
            I => \counterZ0Z_5\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__13751\,
            I => \counterZ0Z_5\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13748\,
            I => \counterZ0Z_5\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__13745\,
            I => \counterZ0Z_5\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__13742\,
            I => \counterZ0Z_5\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__13739\,
            I => \counterZ0Z_5\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__13721\,
            I => \N__13714\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13711\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13708\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13703\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13703\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__13714\,
            I => \counterZ0Z_8\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13711\,
            I => \counterZ0Z_8\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__13708\,
            I => \counterZ0Z_8\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__13703\,
            I => \counterZ0Z_8\
        );

    \I__2100\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__13688\,
            I => slaveselect_1lto9_4
        );

    \I__2097\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__13682\,
            I => slaveselect_1lto9_3
        );

    \I__2095\ : IoInMux
    port map (
            O => \N__13679\,
            I => \N__13675\
        );

    \I__2094\ : IoInMux
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__13675\,
            I => \N__13667\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__13672\,
            I => \N__13667\
        );

    \I__2091\ : IoSpan4Mux
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__2090\ : Span4Mux_s3_h
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__13661\,
            I => \SCLK1_0_i\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__2087\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__13652\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13649\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__13646\,
            I => \un1_sclk17_0_0_cascade_\
        );

    \I__2083\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13639\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13636\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__13639\,
            I => \N__13633\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__13636\,
            I => un39_0_3
        );

    \I__2079\ : Odrv12
    port map (
            O => \N__13633\,
            I => un39_0_3
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__13628\,
            I => \un39_0_3_cascade_\
        );

    \I__2077\ : InMux
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__13619\,
            I => un5_slaveselect_1
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__13616\,
            I => \un5_slaveselect_1_cascade_\
        );

    \I__2073\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13608\
        );

    \I__2072\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13603\
        );

    \I__2071\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13603\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__13608\,
            I => \ScreenBuffer_1_122_1\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__13603\,
            I => \ScreenBuffer_1_122_1\
        );

    \I__2068\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13591\
        );

    \I__2067\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13588\
        );

    \I__2066\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13581\
        );

    \I__2065\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13581\
        );

    \I__2064\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13581\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__13591\,
            I => \N__13578\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__13588\,
            I => un39_0_6
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__13581\,
            I => un39_0_6
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__13578\,
            I => un39_0_6
        );

    \I__2059\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__13568\,
            I => \ScreenBuffer_1_2_1_sqmuxa\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \ScreenBuffer_1_2_1_sqmuxa_cascade_\
        );

    \I__2056\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13558\
        );

    \I__2055\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13550\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13547\
        );

    \I__2053\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13540\
        );

    \I__2052\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13540\
        );

    \I__2051\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13540\
        );

    \I__2050\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13537\
        );

    \I__2049\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13534\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__13550\,
            I => \N__13527\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__13547\,
            I => \N__13527\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__13540\,
            I => \N__13527\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__13537\,
            I => un10_slaveselect
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__13534\,
            I => un10_slaveselect
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__13527\,
            I => un10_slaveselect
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__13520\,
            I => \slaveselect_RNILOQC2Z0Z_0_cascade_\
        );

    \I__2041\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13513\
        );

    \I__2040\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13510\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__13513\,
            I => \N__13507\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13503\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__13507\,
            I => \N__13500\
        );

    \I__2036\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13497\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__13503\,
            I => \Z_decfrac4_2\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__13500\,
            I => \Z_decfrac4_2\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__13497\,
            I => \Z_decfrac4_2\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \ScreenBuffer_1_122_1_cascade_\
        );

    \I__2031\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13481\
        );

    \I__2030\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13481\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__13481\,
            I => \ScreenBuffer_1_3_1_sqmuxa\
        );

    \I__2028\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__13472\,
            I => \ScreenBuffer_1_0_1_sqmuxa\
        );

    \I__2025\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13462\
        );

    \I__2024\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13462\
        );

    \I__2023\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13459\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__13462\,
            I => \N__13456\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__13459\,
            I => \Z_decfrac4\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__13456\,
            I => \Z_decfrac4\
        );

    \I__2019\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__13445\,
            I => voltage_2_9_iv_0_0
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__13442\,
            I => \un1_voltage_2_1_axb_0_cascade_\
        );

    \I__2015\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__13436\,
            I => voltage_2_9_iv_0_2
        );

    \I__2013\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__13424\,
            I => \voltage_2_RNO_0Z0Z_2\
        );

    \I__2009\ : InMux
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__13415\,
            I => \N__13409\
        );

    \I__2006\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13402\
        );

    \I__2005\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13402\
        );

    \I__2004\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13402\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__13409\,
            I => un1_voltage_012_3_0
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__13402\,
            I => un1_voltage_012_3_0
        );

    \I__2001\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__13394\,
            I => \N__13391\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__13391\,
            I => voltage_2_9_iv_0_1
        );

    \I__1998\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13385\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__13379\,
            I => \voltage_2_RNO_0Z0Z_1\
        );

    \I__1994\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__13373\,
            I => \un42_cry_1_c_RNOZ0\
        );

    \I__1992\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__13361\,
            I => \counter_RNIGLLH1Z0Z_0\
        );

    \I__1988\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__13355\,
            I => voltage_011_0
        );

    \I__1986\ : InMux
    port map (
            O => \N__13352\,
            I => un42_cry_3
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__13349\,
            I => \N__13344\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__13348\,
            I => \N__13340\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__13347\,
            I => \N__13337\
        );

    \I__1982\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13331\
        );

    \I__1981\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13331\
        );

    \I__1980\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13326\
        );

    \I__1979\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13326\
        );

    \I__1978\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13323\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N__13320\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13317\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__13323\,
            I => voltage_011
        );

    \I__1974\ : Odrv12
    port map (
            O => \N__13320\,
            I => voltage_011
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__13317\,
            I => voltage_011
        );

    \I__1972\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13302\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13309\,
            I => \N__13297\
        );

    \I__1970\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13297\
        );

    \I__1969\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13294\
        );

    \I__1968\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13289\
        );

    \I__1967\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13289\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__13302\,
            I => \N__13286\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__13297\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__13294\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__13289\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__13286\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__13277\,
            I => \N__13273\
        );

    \I__1960\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13259\
        );

    \I__1959\ : InMux
    port map (
            O => \N__13273\,
            I => \N__13256\
        );

    \I__1958\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13251\
        );

    \I__1957\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13251\
        );

    \I__1956\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13248\
        );

    \I__1955\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13239\
        );

    \I__1954\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13239\
        );

    \I__1953\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13239\
        );

    \I__1952\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13239\
        );

    \I__1951\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13232\
        );

    \I__1950\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13232\
        );

    \I__1949\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13232\
        );

    \I__1948\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13226\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__13259\,
            I => \N__13223\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13212\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__13251\,
            I => \N__13212\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__13248\,
            I => \N__13212\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__13239\,
            I => \N__13212\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__13232\,
            I => \N__13212\
        );

    \I__1941\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13208\
        );

    \I__1940\ : InMux
    port map (
            O => \N__13230\,
            I => \N__13203\
        );

    \I__1939\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13203\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13196\
        );

    \I__1937\ : Span4Mux_s3_v
    port map (
            O => \N__13223\,
            I => \N__13196\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__13212\,
            I => \N__13196\
        );

    \I__1935\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13193\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13190\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__13203\,
            I => \N__13187\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__13196\,
            I => \N__13182\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__13193\,
            I => \N__13182\
        );

    \I__1930\ : Odrv12
    port map (
            O => \N__13190\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__13187\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__13182\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1927\ : InMux
    port map (
            O => \N__13175\,
            I => \N__13171\
        );

    \I__1926\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13168\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__13171\,
            I => \beamY_RNIV42D31Z0Z_6\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__13168\,
            I => \beamY_RNIV42D31Z0Z_6\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__13163\,
            I => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13153\
        );

    \I__1921\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13150\
        );

    \I__1920\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13147\
        );

    \I__1919\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13142\
        );

    \I__1918\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13142\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__13153\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__13150\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__13147\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__13142\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__1913\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13130\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__13130\,
            I => \un113_pixel_3_0_11__g0_0_x2_0Z0Z_0\
        );

    \I__1911\ : CEMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__13121\,
            I => \un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0\
        );

    \I__1908\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13114\
        );

    \I__1907\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13111\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__13114\,
            I => \N__13108\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13103\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__13108\,
            I => \N__13103\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__13103\,
            I => \N_1520\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \N__13097\
        );

    \I__1901\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__1899\ : Span4Mux_s2_h
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__13088\,
            I => \N__13085\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__13085\,
            I => \un1_voltage_2_1_cry_0_c_RNOZ0\
        );

    \I__1896\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__13079\,
            I => \N__13076\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__13076\,
            I => if_generate_plus_mult1_un75_sum_c5_x0
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \if_generate_plus_mult1_un75_sum_c5_x1_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13065\
        );

    \I__1891\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13060\
        );

    \I__1890\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13060\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__13065\,
            I => \beamY_RNIPNEA3_0Z0Z_6\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__13060\,
            I => \beamY_RNIPNEA3_0Z0Z_6\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13049\
        );

    \I__1886\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13049\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__13049\,
            I => \beamY_RNI0K169Z0Z_6\
        );

    \I__1884\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13041\
        );

    \I__1883\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13036\
        );

    \I__1882\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13036\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__13041\,
            I => \N__13033\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__13036\,
            I => \N__13030\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__13033\,
            I => chary_if_generate_plus_mult1_un61_sum_c4
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__13030\,
            I => chary_if_generate_plus_mult1_un61_sum_c4
        );

    \I__1877\ : InMux
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__13022\,
            I => \N__13019\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__13019\,
            I => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__13016\,
            I => \chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\
        );

    \I__1873\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13008\
        );

    \I__1872\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13005\
        );

    \I__1871\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13002\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__12998\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__13005\,
            I => \N__12993\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13002\,
            I => \N__12993\
        );

    \I__1867\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12990\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__12998\,
            I => \N__12981\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__12993\,
            I => \N__12981\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__12990\,
            I => \N__12981\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__12989\,
            I => \N__12974\
        );

    \I__1862\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12967\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__12981\,
            I => \N__12964\
        );

    \I__1860\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12959\
        );

    \I__1859\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12959\
        );

    \I__1858\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12954\
        );

    \I__1857\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12954\
        );

    \I__1856\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12949\
        );

    \I__1855\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12949\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12942\
        );

    \I__1853\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12942\
        );

    \I__1852\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12942\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__12967\,
            I => \beamYZ0Z_6\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__12964\,
            I => \beamYZ0Z_6\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__12959\,
            I => \beamYZ0Z_6\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__12954\,
            I => \beamYZ0Z_6\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__12949\,
            I => \beamYZ0Z_6\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__12942\,
            I => \beamYZ0Z_6\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__12929\,
            I => \N__12925\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__12928\,
            I => \N__12922\
        );

    \I__1843\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12918\
        );

    \I__1842\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12915\
        );

    \I__1841\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12912\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__12918\,
            I => \N__12908\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__12915\,
            I => \N__12903\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__12912\,
            I => \N__12903\
        );

    \I__1837\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12900\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__12908\,
            I => \N__12891\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__12903\,
            I => \N__12891\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__12900\,
            I => \N__12891\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__12899\,
            I => \N__12887\
        );

    \I__1832\ : InMux
    port map (
            O => \N__12898\,
            I => \N__12876\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__12891\,
            I => \N__12873\
        );

    \I__1830\ : InMux
    port map (
            O => \N__12890\,
            I => \N__12866\
        );

    \I__1829\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12866\
        );

    \I__1828\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12866\
        );

    \I__1827\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12861\
        );

    \I__1826\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12861\
        );

    \I__1825\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12856\
        );

    \I__1824\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12856\
        );

    \I__1823\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12849\
        );

    \I__1822\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12849\
        );

    \I__1821\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12849\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__12876\,
            I => \beamYZ0Z_5\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__12873\,
            I => \beamYZ0Z_5\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__12866\,
            I => \beamYZ0Z_5\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__12861\,
            I => \beamYZ0Z_5\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__12856\,
            I => \beamYZ0Z_5\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__12849\,
            I => \beamYZ0Z_5\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__12833\,
            I => \chary_if_generate_plus_mult1_un75_sum_c5_N_9\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__12830\,
            I => \beamY_RNIPLAE31Z0Z_4_cascade_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__12824\,
            I => chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__12821\,
            I => \N__12814\
        );

    \I__1808\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12806\
        );

    \I__1807\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12806\
        );

    \I__1806\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12806\
        );

    \I__1805\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12803\
        );

    \I__1804\ : InMux
    port map (
            O => \N__12814\,
            I => \N__12798\
        );

    \I__1803\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12798\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__12806\,
            I => \beamY_RNIV42D31_0Z0Z_6\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__12803\,
            I => \beamY_RNIV42D31_0Z0Z_6\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__12798\,
            I => \beamY_RNIV42D31_0Z0Z_6\
        );

    \I__1799\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__12788\,
            I => \un113_pixel_3_0_11__N_4_i_0\
        );

    \I__1797\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__12782\,
            I => g1_0_0
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__12779\,
            I => \row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12772\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__12775\,
            I => \N__12769\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12765\
        );

    \I__1791\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12762\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__12768\,
            I => \N__12758\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__12765\,
            I => \N__12753\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__12762\,
            I => \N__12753\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12750\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12746\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__12753\,
            I => \N__12742\
        );

    \I__1784\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12737\
        );

    \I__1783\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12737\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__12746\,
            I => \N__12734\
        );

    \I__1781\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12731\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__12742\,
            I => un5_visibley_c5
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__12737\,
            I => un5_visibley_c5
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__12734\,
            I => un5_visibley_c5
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__12731\,
            I => un5_visibley_c5
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__12722\,
            I => \N__12716\
        );

    \I__1775\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12711\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12711\
        );

    \I__1773\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12708\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12705\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__12711\,
            I => \N__12702\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__12708\,
            I => \beamY_RNIJNLCZ0Z_9\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12705\,
            I => \beamY_RNIJNLCZ0Z_9\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__12702\,
            I => \beamY_RNIJNLCZ0Z_9\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__12695\,
            I => \beamY_RNIJNLCZ0Z_9_cascade_\
        );

    \I__1766\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12682\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12682\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12679\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12673\
        );

    \I__1762\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12670\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12665\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__12682\,
            I => \N__12660\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12657\
        );

    \I__1758\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12650\
        );

    \I__1757\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12650\
        );

    \I__1756\ : InMux
    port map (
            O => \N__12676\,
            I => \N__12650\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__12673\,
            I => \N__12645\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12645\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12640\
        );

    \I__1752\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12640\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__12665\,
            I => \N__12637\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__12664\,
            I => \N__12633\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__12663\,
            I => \N__12628\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__12660\,
            I => \N__12618\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__12657\,
            I => \N__12618\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__12650\,
            I => \N__12618\
        );

    \I__1745\ : Span4Mux_s1_v
    port map (
            O => \N__12645\,
            I => \N__12615\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__12640\,
            I => \N__12612\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__12637\,
            I => \N__12609\
        );

    \I__1742\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12606\
        );

    \I__1741\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12597\
        );

    \I__1740\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12597\
        );

    \I__1739\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12597\
        );

    \I__1738\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12597\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12590\
        );

    \I__1736\ : InMux
    port map (
            O => \N__12626\,
            I => \N__12590\
        );

    \I__1735\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12590\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__12618\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__12615\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1732\ : Odrv12
    port map (
            O => \N__12612\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__12609\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__12606\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__12597\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__12590\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \N__12571\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__1725\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12560\
        );

    \I__1724\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12560\
        );

    \I__1723\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12560\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__12560\,
            I => \beamY_RNIVGU01Z0Z_9\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__12557\,
            I => \N__12552\
        );

    \I__1720\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12549\
        );

    \I__1719\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12546\
        );

    \I__1718\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12541\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__12549\,
            I => \N__12536\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12536\
        );

    \I__1715\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12533\
        );

    \I__1714\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12530\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__12541\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__12536\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__12533\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__12530\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__12521\,
            I => \N__12517\
        );

    \I__1708\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12514\
        );

    \I__1707\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12511\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__12514\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__12511\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__12506\,
            I => \N__12502\
        );

    \I__1703\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12496\
        );

    \I__1702\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12496\
        );

    \I__1701\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12493\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12490\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__12493\,
            I => row_1_if_generate_plus_mult1_un75_sum_ac0_5
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__12490\,
            I => row_1_if_generate_plus_mult1_un75_sum_ac0_5
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__12485\,
            I => \N__12482\
        );

    \I__1696\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12474\
        );

    \I__1695\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12464\
        );

    \I__1694\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12459\
        );

    \I__1693\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12459\
        );

    \I__1692\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12450\
        );

    \I__1691\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12447\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12444\
        );

    \I__1689\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12439\
        );

    \I__1688\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12439\
        );

    \I__1687\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12432\
        );

    \I__1686\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12432\
        );

    \I__1685\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12432\
        );

    \I__1684\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12427\
        );

    \I__1683\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12427\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__12464\,
            I => \N__12422\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__12459\,
            I => \N__12422\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__12458\,
            I => \N__12419\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__12457\,
            I => \N__12416\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12412\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__12455\,
            I => \N__12409\
        );

    \I__1676\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12402\
        );

    \I__1675\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12402\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__12450\,
            I => \N__12397\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__12447\,
            I => \N__12397\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__12444\,
            I => \N__12394\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__12439\,
            I => \N__12391\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__12432\,
            I => \N__12386\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__12427\,
            I => \N__12386\
        );

    \I__1668\ : Span4Mux_h
    port map (
            O => \N__12422\,
            I => \N__12383\
        );

    \I__1667\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12374\
        );

    \I__1666\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12374\
        );

    \I__1665\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12374\
        );

    \I__1664\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12374\
        );

    \I__1663\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12367\
        );

    \I__1662\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12367\
        );

    \I__1661\ : InMux
    port map (
            O => \N__12407\,
            I => \N__12367\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12362\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__12397\,
            I => \N__12362\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__12394\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1657\ : Odrv12
    port map (
            O => \N__12391\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1656\ : Odrv12
    port map (
            O => \N__12386\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__12383\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__12374\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__12367\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__12362\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1651\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12344\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__1649\ : Odrv12
    port map (
            O => \N__12341\,
            I => \un113_pixel_4_0_15__un1_beamylto9_3\
        );

    \I__1648\ : IoInMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__12335\,
            I => \N__12332\
        );

    \I__1646\ : Span4Mux_s3_v
    port map (
            O => \N__12332\,
            I => \N__12329\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__12329\,
            I => \VSync_c\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__12326\,
            I => \un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_\
        );

    \I__1643\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12317\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__12317\,
            I => \beamY_RNII8O41Z0Z_9\
        );

    \I__1640\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12311\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__12311\,
            I => \un113_pixel_4_0_15__g0_i_a3_0Z0Z_4\
        );

    \I__1638\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__12305\,
            I => if_m1_5
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \if_generate_plus_mult1_un54_sum_axbxc5_cascade_\
        );

    \I__1635\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12294\
        );

    \I__1634\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12287\
        );

    \I__1633\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12287\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__12294\,
            I => \N__12283\
        );

    \I__1631\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12278\
        );

    \I__1630\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12278\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__12287\,
            I => \N__12275\
        );

    \I__1628\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12272\
        );

    \I__1627\ : Span4Mux_h
    port map (
            O => \N__12283\,
            I => \N__12269\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__12278\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\
        );

    \I__1625\ : Odrv12
    port map (
            O => \N__12275\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__12272\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__12269\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\
        );

    \I__1622\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__12257\,
            I => if_generate_plus_mult1_un75_sum_ac0_5_x1
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__12254\,
            I => \row_1_if_i2_mux_0_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__12248\,
            I => if_generate_plus_mult1_un75_sum_ac0_5_x0
        );

    \I__1617\ : InMux
    port map (
            O => \N__12245\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__1616\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12236\
        );

    \I__1615\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12236\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__12236\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579\
        );

    \I__1613\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__12230\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4\
        );

    \I__1611\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12221\
        );

    \I__1610\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12221\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__12221\,
            I => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36\
        );

    \I__1608\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__12215\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__12212\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_\
        );

    \I__1605\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__12206\,
            I => chessboardpixel_un173_pixellt10
        );

    \I__1603\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__12200\,
            I => chessboardpixel_un151_pixel_27
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__12197\,
            I => \chessboardpixel_un177_pixel_26_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12188\
        );

    \I__1599\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12188\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__12188\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0\
        );

    \I__1597\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12179\
        );

    \I__1596\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12179\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__12179\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0\
        );

    \I__1594\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12169\
        );

    \I__1593\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12162\
        );

    \I__1592\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12162\
        );

    \I__1591\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12162\
        );

    \I__1590\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12159\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__12169\,
            I => \beamY_i_2\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__12162\,
            I => \beamY_i_2\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__12159\,
            I => \beamY_i_2\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \N__12147\
        );

    \I__1585\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12144\
        );

    \I__1584\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12139\
        );

    \I__1583\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12139\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__12144\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__12139\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_\
        );

    \I__1579\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__12128\,
            I => chessboardpixel_un199_pixellt10
        );

    \I__1577\ : InMux
    port map (
            O => \N__12125\,
            I => counter_cry_4
        );

    \I__1576\ : InMux
    port map (
            O => \N__12122\,
            I => counter_cry_5
        );

    \I__1575\ : InMux
    port map (
            O => \N__12119\,
            I => counter_cry_6
        );

    \I__1574\ : InMux
    port map (
            O => \N__12116\,
            I => counter_cry_7
        );

    \I__1573\ : InMux
    port map (
            O => \N__12113\,
            I => \bfn_4_14_0_\
        );

    \I__1572\ : SRMux
    port map (
            O => \N__12110\,
            I => \N__12106\
        );

    \I__1571\ : SRMux
    port map (
            O => \N__12109\,
            I => \N__12103\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__12106\,
            I => \N__12099\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__12103\,
            I => \N__12096\
        );

    \I__1568\ : SRMux
    port map (
            O => \N__12102\,
            I => \N__12093\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__12099\,
            I => \N__12090\
        );

    \I__1566\ : Span4Mux_s3_v
    port map (
            O => \N__12096\,
            I => \N__12085\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__12093\,
            I => \N__12085\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__12090\,
            I => un1_counter_i_0
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__12085\,
            I => un1_counter_i_0
        );

    \I__1562\ : InMux
    port map (
            O => \N__12080\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1561\ : InMux
    port map (
            O => \N__12077\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__1560\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12068\
        );

    \I__1559\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12068\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__12068\,
            I => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__1557\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12059\
        );

    \I__1556\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12059\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__12059\,
            I => \slaveselect_RNILOQC2Z0Z_2\
        );

    \I__1554\ : InMux
    port map (
            O => \N__12056\,
            I => counter_cry_1
        );

    \I__1553\ : InMux
    port map (
            O => \N__12053\,
            I => counter_cry_2
        );

    \I__1552\ : InMux
    port map (
            O => \N__12050\,
            I => counter_cry_3
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__12047\,
            I => \un1_voltage_012_0_cascade_\
        );

    \I__1550\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12039\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__12043\,
            I => \N__12035\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__12042\,
            I => \N__12032\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12028\
        );

    \I__1546\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12025\
        );

    \I__1545\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12022\
        );

    \I__1544\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12017\
        );

    \I__1543\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12017\
        );

    \I__1542\ : Span4Mux_h
    port map (
            O => \N__12028\,
            I => \N__12014\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__12025\,
            I => un74_voltage_0
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__12022\,
            I => un74_voltage_0
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__12017\,
            I => un74_voltage_0
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__12014\,
            I => un74_voltage_0
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__12005\,
            I => \N__12000\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11997\
        );

    \I__1535\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11992\
        );

    \I__1534\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11992\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11987\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__11992\,
            I => \N__11987\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__11984\,
            I => \N_1153\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__11981\,
            I => \N__11977\
        );

    \I__1528\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11970\
        );

    \I__1527\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11970\
        );

    \I__1526\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11967\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__11975\,
            I => \N__11964\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__11970\,
            I => \N__11958\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__11967\,
            I => \N__11955\
        );

    \I__1522\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11952\
        );

    \I__1521\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11945\
        );

    \I__1520\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11945\
        );

    \I__1519\ : InMux
    port map (
            O => \N__11961\,
            I => \N__11945\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__11958\,
            I => voltage_0_1_sqmuxa_1
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__11955\,
            I => voltage_0_1_sqmuxa_1
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__11952\,
            I => voltage_0_1_sqmuxa_1
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__11945\,
            I => voltage_0_1_sqmuxa_1
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__11936\,
            I => \N_1153_cascade_\
        );

    \I__1513\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11928\
        );

    \I__1512\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11925\
        );

    \I__1511\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11922\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__11928\,
            I => \N__11916\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__11925\,
            I => \N__11916\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__11922\,
            I => \N__11909\
        );

    \I__1507\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11906\
        );

    \I__1506\ : Span4Mux_h
    port map (
            O => \N__11916\,
            I => \N__11903\
        );

    \I__1505\ : InMux
    port map (
            O => \N__11915\,
            I => \N__11898\
        );

    \I__1504\ : InMux
    port map (
            O => \N__11914\,
            I => \N__11898\
        );

    \I__1503\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11893\
        );

    \I__1502\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11893\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__11909\,
            I => voltage_3_1_sqmuxa
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__11906\,
            I => voltage_3_1_sqmuxa
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__11903\,
            I => voltage_3_1_sqmuxa
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__11898\,
            I => voltage_3_1_sqmuxa
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__11893\,
            I => voltage_3_1_sqmuxa
        );

    \I__1496\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11879\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__11876\,
            I => \N__11873\
        );

    \I__1493\ : Span4Mux_h
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__11870\,
            I => \voltage_3_RNO_0Z0Z_1\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__11867\,
            I => \voltage_3_9_iv_0_1_cascade_\
        );

    \I__1490\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11853\
        );

    \I__1489\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11853\
        );

    \I__1488\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11848\
        );

    \I__1487\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11848\
        );

    \I__1486\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11841\
        );

    \I__1485\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11841\
        );

    \I__1484\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11841\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11836\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__11848\,
            I => \N__11833\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__11841\,
            I => \N__11830\
        );

    \I__1480\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11825\
        );

    \I__1479\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11825\
        );

    \I__1478\ : Span4Mux_s3_h
    port map (
            O => \N__11836\,
            I => \N__11822\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__11833\,
            I => \N__11819\
        );

    \I__1476\ : Span4Mux_s3_h
    port map (
            O => \N__11830\,
            I => \N__11816\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__11825\,
            I => un1_voltage_012_0
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__11822\,
            I => un1_voltage_012_0
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__11819\,
            I => un1_voltage_012_0
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__11816\,
            I => un1_voltage_012_0
        );

    \I__1471\ : InMux
    port map (
            O => \N__11807\,
            I => \N__11804\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__11804\,
            I => \N__11801\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__11801\,
            I => voltage_1_9_iv_0_1
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__11798\,
            I => \N__11795\
        );

    \I__1467\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__11792\,
            I => \N__11789\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__11786\,
            I => \voltage_1_RNO_0Z0Z_1\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__11783\,
            I => \N_1504_cascade_\
        );

    \I__1462\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__11777\,
            I => \N_1504\
        );

    \I__1460\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11766\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11766\
        );

    \I__1458\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11762\
        );

    \I__1457\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11758\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11755\
        );

    \I__1455\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11752\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__11762\,
            I => \N__11749\
        );

    \I__1453\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11746\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__11758\,
            I => \N__11743\
        );

    \I__1451\ : Span4Mux_s3_h
    port map (
            O => \N__11755\,
            I => \N__11740\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__11752\,
            I => \N__11735\
        );

    \I__1449\ : Span4Mux_s3_h
    port map (
            O => \N__11749\,
            I => \N__11735\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__11746\,
            I => \counter_RNI8DLH1Z0Z_0\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__11743\,
            I => \counter_RNI8DLH1Z0Z_0\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__11740\,
            I => \counter_RNI8DLH1Z0Z_0\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__11735\,
            I => \counter_RNI8DLH1Z0Z_0\
        );

    \I__1444\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11721\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__11725\,
            I => \N__11718\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__11724\,
            I => \N__11715\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11711\
        );

    \I__1440\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11704\
        );

    \I__1439\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11704\
        );

    \I__1438\ : InMux
    port map (
            O => \N__11714\,
            I => \N__11704\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__11711\,
            I => \N_1508\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__11704\,
            I => \N_1508\
        );

    \I__1435\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11690\
        );

    \I__1434\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11690\
        );

    \I__1433\ : InMux
    port map (
            O => \N__11697\,
            I => \N__11690\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__11690\,
            I => \N__11687\
        );

    \I__1431\ : Odrv12
    port map (
            O => \N__11687\,
            I => \N_1159_i\
        );

    \I__1430\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__11681\,
            I => \N__11675\
        );

    \I__1428\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11668\
        );

    \I__1427\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11668\
        );

    \I__1426\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11668\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__11675\,
            I => \N__11665\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N_1154\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__11665\,
            I => \N_1154\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__11660\,
            I => \N_1159_i_cascade_\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__11657\,
            I => \N__11652\
        );

    \I__1420\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11649\
        );

    \I__1419\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11646\
        );

    \I__1418\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11639\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__11649\,
            I => \N__11634\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__11646\,
            I => \N__11634\
        );

    \I__1415\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11631\
        );

    \I__1414\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11624\
        );

    \I__1413\ : InMux
    port map (
            O => \N__11643\,
            I => \N__11624\
        );

    \I__1412\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11624\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__11639\,
            I => \N__11619\
        );

    \I__1410\ : Span4Mux_h
    port map (
            O => \N__11634\,
            I => \N__11619\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__11631\,
            I => voltage_2_1_sqmuxa
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__11624\,
            I => voltage_2_1_sqmuxa
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__11619\,
            I => voltage_2_1_sqmuxa
        );

    \I__1406\ : IoInMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1404\ : Span4Mux_s3_h
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__11603\,
            I => voltage_0_0_sqmuxa_1
        );

    \I__1402\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__11597\,
            I => \slaveselect_RNILOQC2Z0Z_1\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__11594\,
            I => \slaveselect_RNILOQC2Z0Z_1_cascade_\
        );

    \I__1399\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__11588\,
            I => \N__11584\
        );

    \I__1397\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__11584\,
            I => \N__11578\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__11581\,
            I => \counter_RNICHLH1Z0Z_0\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__11578\,
            I => \counter_RNICHLH1Z0Z_0\
        );

    \I__1393\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__11570\,
            I => un5_visibley_0_29
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__11567\,
            I => \chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__11564\,
            I => \if_m1_x1_cascade_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11557\
        );

    \I__1388\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11553\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__11557\,
            I => \N__11550\
        );

    \I__1386\ : InMux
    port map (
            O => \N__11556\,
            I => \N__11547\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__11553\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__11550\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__11547\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1382\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11534\
        );

    \I__1381\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11534\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__1379\ : Span4Mux_h
    port map (
            O => \N__11531\,
            I => \N__11523\
        );

    \I__1378\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11516\
        );

    \I__1377\ : InMux
    port map (
            O => \N__11529\,
            I => \N__11516\
        );

    \I__1376\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11516\
        );

    \I__1375\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11511\
        );

    \I__1374\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11511\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__11523\,
            I => row_1_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__11516\,
            I => row_1_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__11511\,
            I => row_1_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__1370\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__11501\,
            I => if_m1_x0
        );

    \I__1368\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__11495\,
            I => \un113_pixel_3_0_11__g1_0\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__11492\,
            I => \chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_\
        );

    \I__1365\ : IoInMux
    port map (
            O => \N__11489\,
            I => \N__11486\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__1363\ : Span4Mux_s3_h
    port map (
            O => \N__11483\,
            I => \N__11480\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__11477\,
            I => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__11474\,
            I => \beamY_RNIQTGS2Z0Z_8_cascade_\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__11471\,
            I => \chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__11468\,
            I => \chary_if_generate_plus_mult1_un61_sum_axb3_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11459\
        );

    \I__1356\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11459\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__11459\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__11456\,
            I => \N__11451\
        );

    \I__1353\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11438\
        );

    \I__1352\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11438\
        );

    \I__1351\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11438\
        );

    \I__1350\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11438\
        );

    \I__1349\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11438\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__11438\,
            I => \beamY_RNIQTGS2Z0Z_8\
        );

    \I__1347\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11429\
        );

    \I__1346\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11429\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__11429\,
            I => chary_if_generate_plus_mult1_un54_sum_c4
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__11426\,
            I => \beamY_RNI0K169Z0Z_6_cascade_\
        );

    \I__1343\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11420\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__11420\,
            I => chary_if_generate_plus_mult1_un61_sum_c4_3_1
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__11417\,
            I => \chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__11414\,
            I => \N__11410\
        );

    \I__1339\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11405\
        );

    \I__1338\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11405\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__11405\,
            I => \N__11401\
        );

    \I__1336\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11398\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__11401\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__11398\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0
        );

    \I__1333\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11390\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__11390\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_6_2
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__11387\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_\
        );

    \I__1330\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11378\
        );

    \I__1329\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11378\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__11378\,
            I => \N__11374\
        );

    \I__1327\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11371\
        );

    \I__1326\ : Span4Mux_h
    port map (
            O => \N__11374\,
            I => \N__11368\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__11371\,
            I => row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__11368\,
            I => row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__1322\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11353\
        );

    \I__1321\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11353\
        );

    \I__1320\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11350\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__11353\,
            I => \N__11347\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11344\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__11344\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__11341\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0\
        );

    \I__1314\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11331\
        );

    \I__1313\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11326\
        );

    \I__1312\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11326\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__11331\,
            I => \N__11323\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11320\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__11323\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__11320\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__1306\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__11309\,
            I => \beamY_RNIFS4TZ0Z_7\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__11306\,
            I => \beamY_RNIFS4TZ0Z_7_cascade_\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__11303\,
            I => \chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_\
        );

    \I__1302\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__11297\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__1300\ : InMux
    port map (
            O => \N__11294\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__1298\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__11285\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \N__11279\
        );

    \I__1295\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__11273\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__1292\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__11267\,
            I => \N__11264\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__11264\,
            I => \N__11260\
        );

    \I__1289\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11257\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__11260\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__11257\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0
        );

    \I__1286\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__11249\,
            I => \N__11242\
        );

    \I__1284\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11239\
        );

    \I__1283\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11236\
        );

    \I__1282\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11231\
        );

    \I__1281\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11231\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__11242\,
            I => un5_visibley_c2
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__11239\,
            I => un5_visibley_c2
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__11236\,
            I => un5_visibley_c2
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__11231\,
            I => un5_visibley_c2
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__11222\,
            I => \chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_\
        );

    \I__1275\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11216\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__11216\,
            I => \beamY_RNIEDF31Z0Z_6\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__11213\,
            I => \chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1271\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__11204\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246\
        );

    \I__1269\ : InMux
    port map (
            O => \N__11201\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__1268\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__11195\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__1266\ : InMux
    port map (
            O => \N__11192\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__11189\,
            I => \N__11184\
        );

    \I__1264\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11179\
        );

    \I__1263\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11170\
        );

    \I__1262\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11170\
        );

    \I__1261\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11170\
        );

    \I__1260\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11170\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__11179\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__11170\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8\
        );

    \I__1257\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__11162\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__1255\ : InMux
    port map (
            O => \N__11159\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1253\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__11150\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79\
        );

    \I__1251\ : InMux
    port map (
            O => \N__11147\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1249\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__11138\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0\
        );

    \I__1247\ : InMux
    port map (
            O => \N__11135\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__1245\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__11126\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0\
        );

    \I__1243\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11114\
        );

    \I__1242\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11114\
        );

    \I__1241\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11111\
        );

    \I__1240\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11106\
        );

    \I__1239\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11106\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__11114\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__11111\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__11106\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__11096\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1232\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1230\ : Odrv12
    port map (
            O => \N__11084\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1\
        );

    \I__1229\ : InMux
    port map (
            O => \N__11081\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1227\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__11069\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2\
        );

    \I__1224\ : InMux
    port map (
            O => \N__11066\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1222\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__11054\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513\
        );

    \I__1219\ : InMux
    port map (
            O => \N__11051\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__1218\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__11042\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__1215\ : InMux
    port map (
            O => \N__11039\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__1214\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11029\
        );

    \I__1213\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11022\
        );

    \I__1212\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11022\
        );

    \I__1211\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11022\
        );

    \I__1210\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11019\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__11029\,
            I => \N__11014\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__11022\,
            I => \N__11014\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__11019\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__11014\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73\
        );

    \I__1205\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__11006\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__1203\ : InMux
    port map (
            O => \N__11003\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__1202\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10997\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__10997\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404\
        );

    \I__1200\ : InMux
    port map (
            O => \N__10994\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__10991\,
            I => \N__10988\
        );

    \I__1198\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__10985\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45\
        );

    \I__1196\ : InMux
    port map (
            O => \N__10982\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1195\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__10976\,
            I => \counter_RNI2RBA2Z0Z_3\
        );

    \I__1193\ : InMux
    port map (
            O => \N__10973\,
            I => un1_voltage_2_1_cry_1
        );

    \I__1192\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__10967\,
            I => un1_voltage_2_1_axb_3
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1189\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__10955\,
            I => voltage_2_9_iv_0_3
        );

    \I__1186\ : InMux
    port map (
            O => \N__10952\,
            I => un1_voltage_2_1_cry_2
        );

    \I__1185\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10941\
        );

    \I__1184\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10941\
        );

    \I__1183\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10936\
        );

    \I__1182\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10936\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__10941\,
            I => \N__10933\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N_46_1\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__10933\,
            I => \N_46_1\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__10928\,
            I => \un1_sclk17_2_1_cascade_\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__10925\,
            I => \un1_sclk17_1_1_cascade_\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1175\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1173\ : Odrv12
    port map (
            O => \N__10913\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__1172\ : InMux
    port map (
            O => \N__10910\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__1170\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__10901\,
            I => \counter_RNILOUG2Z0Z_3\
        );

    \I__1168\ : InMux
    port map (
            O => \N__10898\,
            I => un1_voltage_1_1_cry_0
        );

    \I__1167\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__10892\,
            I => \counter_RNIT58K2Z0Z_2\
        );

    \I__1165\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1163\ : Odrv12
    port map (
            O => \N__10883\,
            I => \voltage_1_RNO_0Z0Z_2\
        );

    \I__1162\ : InMux
    port map (
            O => \N__10880\,
            I => un1_voltage_1_1_cry_1
        );

    \I__1161\ : InMux
    port map (
            O => \N__10877\,
            I => un1_voltage_1_1_cry_2
        );

    \I__1160\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__10871\,
            I => \voltage_1_RNO_0Z0Z_3\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__10868\,
            I => \un6_slaveselectlto9_1_cascade_\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__10865\,
            I => \un6_slaveselect_0_cascade_\
        );

    \I__1156\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__10859\,
            I => un3_slaveselectlt9
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1153\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__10847\,
            I => \voltage_2_RNIKG123Z0Z_1\
        );

    \I__1150\ : InMux
    port map (
            O => \N__10844\,
            I => un1_voltage_2_1_cry_0
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__10841\,
            I => \voltage_1_1_sqmuxa_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__10835\,
            I => voltage_1_9_iv_0_3
        );

    \I__1146\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__10829\,
            I => \voltage_3_RNO_0Z0Z_3\
        );

    \I__1144\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__10823\,
            I => voltage_3_9_iv_0_3
        );

    \I__1142\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10813\
        );

    \I__1140\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10810\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__10813\,
            I => \N_1510\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N_1510\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__10805\,
            I => \N_1506_cascade_\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__10802\,
            I => \counter_RNIGLLH1Z0Z_0_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__1133\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10783\
        );

    \I__1132\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10783\
        );

    \I__1131\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10783\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__10790\,
            I => \N_2063\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__10783\,
            I => \N_2063\
        );

    \I__1128\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__10772\,
            I => \N_1522\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__1124\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__10760\,
            I => \un1_voltage_1_1_cry_0_0_c_RNOZ0\
        );

    \I__1121\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10751\
        );

    \I__1120\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10751\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__10751\,
            I => \N_1521\
        );

    \I__1118\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10743\
        );

    \I__1117\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10738\
        );

    \I__1116\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10738\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__10743\,
            I => \counter_RNI49LH1_0Z0Z_0\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__10738\,
            I => \counter_RNI49LH1_0Z0Z_0\
        );

    \I__1113\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__10730\,
            I => voltage_1_9_iv_0_0
        );

    \I__1111\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10721\
        );

    \I__1110\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10721\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__10721\,
            I => \CO1_3\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10718\,
            I => \voltage_2_1_sqmuxa_cascade_\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10706\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10706\
        );

    \I__1105\ : InMux
    port map (
            O => \N__10713\,
            I => \N__10706\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N_1155\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__10703\,
            I => \N__10699\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__10702\,
            I => \N__10696\
        );

    \I__1101\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10689\
        );

    \I__1100\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10689\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__10695\,
            I => \N__10686\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__10694\,
            I => \N__10680\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__10689\,
            I => \N__10677\
        );

    \I__1096\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10674\
        );

    \I__1095\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10671\
        );

    \I__1094\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10666\
        );

    \I__1093\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10666\
        );

    \I__1092\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10663\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__10677\,
            I => voltage_1_1_sqmuxa
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__10674\,
            I => voltage_1_1_sqmuxa
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__10671\,
            I => voltage_1_1_sqmuxa
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__10666\,
            I => voltage_1_1_sqmuxa
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__10663\,
            I => voltage_1_1_sqmuxa
        );

    \I__1086\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__10646\,
            I => \voltage_3_RNO_0Z0Z_2\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__10643\,
            I => \voltage_3_9_iv_0_2_cascade_\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \CO2_3_cascade_\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__10637\,
            I => \N_1155_cascade_\
        );

    \I__1080\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__10631\,
            I => voltage_0_10_iv_0_3
        );

    \I__1078\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10624\
        );

    \I__1077\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__10624\,
            I => \N_1519\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__10621\,
            I => \N_1519\
        );

    \I__1074\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__10613\,
            I => if_generate_plus_mult1_un68_sum_axbxc5_x0
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__10610\,
            I => \if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10598\
        );

    \I__1070\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10598\
        );

    \I__1069\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10591\
        );

    \I__1068\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10591\
        );

    \I__1067\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10591\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__10598\,
            I => \N__10586\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10586\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__10586\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8\
        );

    \I__1063\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__10580\,
            I => if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__10577\,
            I => \if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10568\
        );

    \I__1059\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10565\
        );

    \I__1058\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10560\
        );

    \I__1057\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10560\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__10568\,
            I => \beamY_RNI75QM4Z0Z_5\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__10565\,
            I => \beamY_RNI75QM4Z0Z_5\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__10560\,
            I => \beamY_RNI75QM4Z0Z_5\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__10553\,
            I => \voltage_0_10_iv_0_2_cascade_\
        );

    \I__1052\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10547\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__10547\,
            I => \voltage_0_RNO_0Z0Z_2\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \voltage_1_9_iv_0_2_cascade_\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__10541\,
            I => \beamY_RNI9425Z0Z_6_cascade_\
        );

    \I__1048\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__10535\,
            I => if_generate_plus_mult1_un61_sum_ac0_x0
        );

    \I__1046\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__10529\,
            I => if_generate_plus_mult1_un61_sum_ac0_x1
        );

    \I__1044\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10523\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__10523\,
            I => row_1_if_generate_plus_mult1_un61_sum_ac0_6
        );

    \I__1042\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10517\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__10514\,
            I => row_1_if_generate_plus_mult1_un61_sum_c4_d
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__10511\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__10508\,
            I => \beamY_RNI75QM4Z0Z_5_cascade_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__10502\,
            I => row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__10499\,
            I => \chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__10496\,
            I => \beamY_RNI9425_0Z0Z_6_cascade_\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__10493\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__10490\,
            I => \chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_\
        );

    \I__1031\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__10484\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__1029\ : InMux
    port map (
            O => \N__10481\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1027\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__10472\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__10469\,
            I => \un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__10466\,
            I => \un5_visibley_axbxc7_1_cascade_\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__10463\,
            I => \chary_if_generate_plus_mult1_un33_sum_axb3_cascade_\
        );

    \I__1022\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__10454\,
            I => \N_41_i\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__10451\,
            I => \N_41_i_cascade_\
        );

    \I__1018\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10443\
        );

    \I__1017\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10438\
        );

    \I__1016\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10438\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10427\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__10438\,
            I => \N__10427\
        );

    \I__1013\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10422\
        );

    \I__1012\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10422\
        );

    \I__1011\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10415\
        );

    \I__1010\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10415\
        );

    \I__1009\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10415\
        );

    \I__1008\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10412\
        );

    \I__1007\ : Odrv12
    port map (
            O => \N__10427\,
            I => voltage_0_1_sqmuxa
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__10422\,
            I => voltage_0_1_sqmuxa
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__10415\,
            I => voltage_0_1_sqmuxa
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__10412\,
            I => voltage_0_1_sqmuxa
        );

    \I__1003\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__10400\,
            I => \ScreenBuffer_0_1_1_sqmuxa_2\
        );

    \I__1001\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__10388\,
            I => \un4_voltage_2_0__i2_mux\
        );

    \I__997\ : InMux
    port map (
            O => \N__10385\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__996\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__10379\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31\
        );

    \I__994\ : InMux
    port map (
            O => \N__10376\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10369\
        );

    \I__992\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10360\
        );

    \I__991\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10360\
        );

    \I__990\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10360\
        );

    \I__989\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10357\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__10360\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__10357\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__985\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__10346\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1\
        );

    \I__983\ : InMux
    port map (
            O => \N__10343\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__982\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__10337\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10330\
        );

    \I__979\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10327\
        );

    \I__978\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__10327\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__10324\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1\
        );

    \I__975\ : InMux
    port map (
            O => \N__10319\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__10316\,
            I => \un4_voltage_10_9__N_4_cascade_\
        );

    \I__973\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10306\
        );

    \I__971\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10303\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__10306\,
            I => \un4_voltage_2_0__N_5_iZ0\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__10303\,
            I => \un4_voltage_2_0__N_5_iZ0\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \voltage_0_1_sqmuxa_cascade_\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__966\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__964\ : Span4Mux_v
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__10283\,
            I => \un1_voltage_0_cry_0_0_c_RNOZ0\
        );

    \I__962\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N_34_0_i\
        );

    \I__960\ : InMux
    port map (
            O => \N__10274\,
            I => un1_voltage_3_1_cry_1
        );

    \I__959\ : InMux
    port map (
            O => \N__10271\,
            I => un1_voltage_3_1_cry_2
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__10268\,
            I => \N__10264\
        );

    \I__957\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__956\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__10261\,
            I => \ScreenBuffer_0_0_1_sqmuxa\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__10258\,
            I => \ScreenBuffer_0_0_1_sqmuxa\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__10253\,
            I => \un4_voltage_2_0__N_13_mux_iZ0_cascade_\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__951\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__10244\,
            I => \N__10241\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__10241\,
            I => \SDATA1_ibuf_RNI098KZ0Z2\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N_35_0_i_cascade_\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \un1_voltage_1_1_axb_0_cascade_\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__10232\,
            I => \voltage_0_1_sqmuxa_1_cascade_\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__10229\,
            I => \voltage_3_9_iv_0_0_cascade_\
        );

    \I__944\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10222\
        );

    \I__943\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10219\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N_1507\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__10219\,
            I => \N_1507\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__10214\,
            I => \N_1507_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__10208\,
            I => \voltage_3_RNO_0Z0Z_0\
        );

    \I__937\ : InMux
    port map (
            O => \N__10205\,
            I => un1_voltage_3_1_cry_0
        );

    \I__936\ : InMux
    port map (
            O => \N__10202\,
            I => un1_voltage_0_cry_2
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__10199\,
            I => \N_1503_cascade_\
        );

    \I__934\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__10193\,
            I => \SDATA1_ibuf_RNILOUGZ0Z2\
        );

    \I__932\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__10187\,
            I => if_generate_plus_mult1_un75_sum_axbxc5_0_x1
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__10184\,
            I => \if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__10181\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\
        );

    \I__928\ : InMux
    port map (
            O => \N__10178\,
            I => un1_voltage_0_cry_0
        );

    \I__927\ : InMux
    port map (
            O => \N__10175\,
            I => un1_voltage_0_cry_1
        );

    \I__926\ : InMux
    port map (
            O => \N__10172\,
            I => un20_beamy_cry_1
        );

    \I__925\ : InMux
    port map (
            O => \N__10169\,
            I => un20_beamy_cry_2
        );

    \I__924\ : InMux
    port map (
            O => \N__10166\,
            I => un20_beamy_cry_3
        );

    \I__923\ : InMux
    port map (
            O => \N__10163\,
            I => un20_beamy_cry_4
        );

    \I__922\ : InMux
    port map (
            O => \N__10160\,
            I => un20_beamy_cry_5
        );

    \I__921\ : InMux
    port map (
            O => \N__10157\,
            I => un20_beamy_cry_6
        );

    \I__920\ : InMux
    port map (
            O => \N__10154\,
            I => un20_beamy_cry_7
        );

    \I__919\ : InMux
    port map (
            O => \N__10151\,
            I => \bfn_1_7_0_\
        );

    \I__918\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__10145\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\
        );

    \I__916\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__10139\,
            I => \beamY_RNISI4A_0Z0Z_9\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__10136\,
            I => \beamY_RNIE925Z0Z_6_cascade_\
        );

    \I__913\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__10130\,
            I => \beamY_RNIKOP3_0Z0Z_6\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__10127\,
            I => \un5_visibley_c2_cascade_\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__10124\,
            I => \N__10120\
        );

    \I__909\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__908\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10114\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__10117\,
            I => un5_visibley_c6_0_0_0
        );

    \I__906\ : LocalMux
    port map (
            O => \N__10114\,
            I => un5_visibley_c6_0_0_0
        );

    \I__905\ : InMux
    port map (
            O => \N__10109\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__904\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10097\
        );

    \I__903\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10097\
        );

    \I__902\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10090\
        );

    \I__901\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10090\
        );

    \I__900\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10090\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__10097\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__10090\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__896\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__10079\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__894\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10071\
        );

    \I__893\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10066\
        );

    \I__892\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10066\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__10071\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__890\ : LocalMux
    port map (
            O => \N__10066\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__888\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__10055\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0\
        );

    \I__886\ : InMux
    port map (
            O => \N__10052\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__885\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__10046\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0\
        );

    \I__883\ : InMux
    port map (
            O => \N__10043\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__882\ : InMux
    port map (
            O => \N__10040\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__881\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10031\
        );

    \I__880\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10031\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__10031\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__878\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__10025\,
            I => \beamY_RNITSR8_0Z0Z_8\
        );

    \I__876\ : InMux
    port map (
            O => \N__10022\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__875\ : InMux
    port map (
            O => \N__10019\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__10016\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \N__10010\
        );

    \I__872\ : InMux
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__10007\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__869\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9998\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0\
        );

    \I__867\ : InMux
    port map (
            O => \N__9995\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__865\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__9986\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0\
        );

    \I__863\ : InMux
    port map (
            O => \N__9983\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__862\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__9977\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0\
        );

    \I__860\ : InMux
    port map (
            O => \N__9974\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__858\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__9965\,
            I => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__856\ : InMux
    port map (
            O => \N__9962\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__855\ : IoInMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__853\ : IoSpan4Mux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__852\ : IoSpan4Mux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__851\ : IoSpan4Mux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__9944\,
            I => \Clock50MHz.PixelClock\
        );

    \I__849\ : InMux
    port map (
            O => \N__9941\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__848\ : InMux
    port map (
            O => \N__9938\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__847\ : InMux
    port map (
            O => \N__9935\,
            I => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un20_beamy_cry_8,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => counter_cry_8,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_2_0_\
        );

    \IN_MUX_bfv_4_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_1_0_\
        );

    \IN_MUX_bfv_2_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_1_0_\
        );

    \IN_MUX_bfv_1_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_1_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \slaveselect_RNIO5RB1_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11612\,
            GLOBALBUFFEROUTPUT => voltage_0_0_sqmuxa_1_g
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9959\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12688\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_1_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01J31_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10103\,
            in2 => \N__10085\,
            in3 => \N__9941\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI01JZ0Z31\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQI1_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10105\,
            in2 => \N__10004\,
            in3 => \N__9938\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI9JQIZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9P1_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10104\,
            in2 => \N__9992\,
            in3 => \N__9935\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIJJ9PZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI8SH33_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10367\,
            in1 => \N__9980\,
            in2 => \N__10013\,
            in3 => \N__10022\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25A1_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10106\,
            in1 => \N__10076\,
            in2 => \N__9971\,
            in3 => \N__10019\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1\,
            ltout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNII25AZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5ME33_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__10333\,
            in1 => \_gnd_net_\,
            in2 => \N__10016\,
            in3 => \_gnd_net_\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI5MEZ0Z33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_0_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10102\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14002\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7K_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10028\,
            in2 => \N__21913\,
            in3 => \N__9995\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI4C7KZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQ_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21908\,
            in2 => \N__10061\,
            in3 => \N__9983\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDALQZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQ_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10049\,
            in2 => \N__21914\,
            in3 => \N__9974\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFENQZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10074\,
            in2 => \_gnd_net_\,
            in3 => \N__9962\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MG_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10037\,
            in2 => \_gnd_net_\,
            in3 => \N__10109\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIM1MGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14003\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__10075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10036\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10148\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8F_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10142\,
            in2 => \N__21887\,
            in3 => \N__10052\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI5P8FZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9F_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21866\,
            in2 => \N__18283\,
            in3 => \N__10043\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6R9FZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10040\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITSR8_0_8_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18157\,
            lcout => \beamY_RNITSR8_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100111000011"
        )
    port map (
            in0 => \N__14661\,
            in1 => \N__14891\,
            in2 => \N__10124\,
            in3 => \N__11247\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_0_9_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18225\,
            lcout => \beamY_RNISI4A_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIE925_6_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__14782\,
            in1 => \N__12972\,
            in2 => \N__14658\,
            in3 => \N__12881\,
            lcout => OPEN,
            ltout => \beamY_RNIE925Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0DB_6_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10133\,
            in2 => \N__10136\,
            in3 => \N__11248\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKOP3_0_6_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__14781\,
            in1 => \N__12971\,
            in2 => \_gnd_net_\,
            in3 => \N__12880\,
            lcout => \beamY_RNIKOP3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20751\,
            in2 => \_gnd_net_\,
            in3 => \N__14417\,
            lcout => un5_visibley_c2,
            ltout => \un5_visibley_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITSR8_8_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000010101"
        )
    port map (
            in0 => \N__10123\,
            in1 => \N__14617\,
            in2 => \N__10127\,
            in3 => \N__14877\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un40_sum_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKOP3_6_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__14780\,
            in1 => \N__12970\,
            in2 => \_gnd_net_\,
            in3 => \N__12879\,
            lcout => un5_visibley_c6_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_3_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__14621\,
            in2 => \_gnd_net_\,
            in3 => \N__14421\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un20_beamy_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23301\,
            in2 => \N__24859\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => un20_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20789\,
            in2 => \_gnd_net_\,
            in3 => \N__10172\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => un20_beamy_cry_1,
            carryout => un20_beamy_cry_2,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14146\,
            in1 => \N__14440\,
            in2 => \_gnd_net_\,
            in3 => \N__10169\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => un20_beamy_cry_2,
            carryout => un20_beamy_cry_3,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14145\,
            in1 => \N__14657\,
            in2 => \_gnd_net_\,
            in3 => \N__10166\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un20_beamy_cry_3,
            carryout => un20_beamy_cry_4,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12898\,
            in2 => \_gnd_net_\,
            in3 => \N__10163\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un20_beamy_cry_4,
            carryout => un20_beamy_cry_5,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12988\,
            in2 => \_gnd_net_\,
            in3 => \N__10160\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un20_beamy_cry_5,
            carryout => un20_beamy_cry_6,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14147\,
            in1 => \N__14809\,
            in2 => \_gnd_net_\,
            in3 => \N__10157\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => un20_beamy_cry_6,
            carryout => un20_beamy_cry_7,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14889\,
            in2 => \_gnd_net_\,
            in3 => \N__10154\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un20_beamy_cry_7,
            carryout => un20_beamy_cry_8,
            clk => \N__21053\,
            ce => \N__17541\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__14972\,
            in1 => \N__14144\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21052\,
            ce => \N__17546\,
            sr => \_gnd_net_\
        );

    \beamY_RNICE3U5_5_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10604\,
            in2 => \_gnd_net_\,
            in3 => \N__10573\,
            lcout => \r_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x1_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12292\,
            in1 => \N__14519\,
            in2 => \N__12457\,
            in3 => \N__11530\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc5_0_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_x0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12293\,
            in1 => \N__14520\,
            in2 => \N__12458\,
            in3 => \N__11529\,
            lcout => OPEN,
            ltout => \if_generate_plus_mult1_un75_sum_axbxc5_0_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_0_ns_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10190\,
            in2 => \N__10184\,
            in3 => \N__11560\,
            lcout => row_1_if_generate_plus_mult1_un75_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011101000"
        )
    port map (
            in0 => \N__10603\,
            in1 => \N__13211\,
            in2 => \N__12456\,
            in3 => \N__14517\,
            lcout => if_generate_plus_mult1_un68_sum_ac0_7_1_0_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_c4_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__14518\,
            in1 => \N__12415\,
            in2 => \_gnd_net_\,
            in3 => \N__10526\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4\,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_x0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__10605\,
            in1 => \N__10574\,
            in2 => \N__10181\,
            in3 => \N__11528\,
            lcout => if_generate_plus_mult1_un68_sum_axbxc5_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_0_cry_0_0_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18478\,
            in2 => \N__10295\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => un1_voltage_0_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_0_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19052\,
            in2 => \N__10250\,
            in3 => \N__10178\,
            lcout => \voltage_0_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => un1_voltage_0_cry_0,
            carryout => un1_voltage_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_0_2_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10196\,
            in2 => \N__16554\,
            in3 => \N__10175\,
            lcout => \voltage_0_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => un1_voltage_0_cry_1,
            carryout => un1_voltage_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_3_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011101011101"
        )
    port map (
            in0 => \N__10634\,
            in1 => \N__19412\,
            in2 => \N__17983\,
            in3 => \N__10202\,
            lcout => \voltage_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19953\,
            ce => 'H',
            sr => \N__18541\
        );

    \ScreenBuffer_1_0_e_0_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19182\,
            in1 => \N__18505\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => \ScreenBuffer_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19954\,
            ce => \N__18997\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_2_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16584\,
            in1 => \N__19183\,
            in2 => \_gnd_net_\,
            in3 => \N__16544\,
            lcout => \ScreenBuffer_1_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19954\,
            ce => \N__18997\,
            sr => \_gnd_net_\
        );

    \voltage_0_RNITQ2M_0_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15391\,
            in1 => \N__18480\,
            in2 => \_gnd_net_\,
            in3 => \N__15720\,
            lcout => OPEN,
            ltout => \N_1503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI49LH1_0_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16277\,
            in2 => \N__10199\,
            in3 => \N__10225\,
            lcout => \counter_RNI49LH1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNITQ2M_0_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15390\,
            in1 => \N__18479\,
            in2 => \_gnd_net_\,
            in3 => \N__15718\,
            lcout => \N_1519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNI1V2M_0_2_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15719\,
            in1 => \N__15301\,
            in2 => \_gnd_net_\,
            in3 => \N__16543\,
            lcout => \N_1521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_0_0_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10447\,
            in1 => \N__10313\,
            in2 => \_gnd_net_\,
            in3 => \N__18481\,
            lcout => un1_voltage_0_axb_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATA1_ibuf_RNILOUG2_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10397\,
            in2 => \_gnd_net_\,
            in3 => \N__10446\,
            lcout => \SDATA1_ibuf_RNILOUGZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI2ACM1_0_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19180\,
            in1 => \N__16251\,
            in2 => \N__13349\,
            in3 => \N__15739\,
            lcout => voltage_3_1_sqmuxa,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_0_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10460\,
            in1 => \N__15329\,
            in2 => \_gnd_net_\,
            in3 => \N__10448\,
            lcout => OPEN,
            ltout => \un1_voltage_1_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__10733\,
            in1 => \N__11862\,
            in2 => \N__10235\,
            in3 => \N__15740\,
            lcout => \voltage_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19956\,
            ce => 'H',
            sr => \N__18543\
        );

    \counter_RNI2ACM1_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16250\,
            in1 => \N__19179\,
            in2 => \N__15811\,
            in3 => \N__13343\,
            lcout => voltage_0_1_sqmuxa_1,
            ltout => \voltage_0_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_1_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__10226\,
            in1 => \N__11921\,
            in2 => \N__10232\,
            in3 => \N__12038\,
            lcout => OPEN,
            ltout => \voltage_3_9_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_0_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111111001111"
        )
    port map (
            in0 => \N__11861\,
            in1 => \N__10211\,
            in2 => \N__10229\,
            in3 => \N__15814\,
            lcout => \voltage_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19956\,
            ce => 'H',
            sr => \N__18543\
        );

    \voltage_1_RNIV09O_0_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15328\,
            in1 => \N__18503\,
            in2 => \_gnd_net_\,
            in3 => \N__15735\,
            lcout => \N_1507\,
            ltout => \N_1507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI49LH1_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16249\,
            in1 => \_gnd_net_\,
            in2 => \N__10214\,
            in3 => \N__10627\,
            lcout => un74_voltage_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_0_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18504\,
            in2 => \N__10268\,
            in3 => \N__10267\,
            lcout => \voltage_3_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => un1_voltage_3_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_0_1_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19369\,
            in2 => \_gnd_net_\,
            in3 => \N__10205\,
            lcout => \voltage_3_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => un1_voltage_3_1_cry_0,
            carryout => un1_voltage_3_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_0_2_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16585\,
            in2 => \_gnd_net_\,
            in3 => \N__10274\,
            lcout => \voltage_3_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => un1_voltage_3_1_cry_1,
            carryout => un1_voltage_3_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_0_3_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19450\,
            in2 => \_gnd_net_\,
            in3 => \N__10271\,
            lcout => \voltage_3_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI4CSO_3_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16244\,
            in1 => \N__16407\,
            in2 => \N__15755\,
            in3 => \N__15467\,
            lcout => \ScreenBuffer_0_0_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIAV5D_4_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__13864\,
            in1 => \N__16361\,
            in2 => \_gnd_net_\,
            in3 => \N__13506\,
            lcout => un3_slaveselectlt9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_voltage_2_0__N_13_mux_i_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011110000100"
        )
    port map (
            in0 => \N__15976\,
            in1 => \N__10948\,
            in2 => \N__15754\,
            in3 => \N__16362\,
            lcout => OPEN,
            ltout => \un4_voltage_2_0__N_13_mux_iZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATA1_ibuf_RNI098K2_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10253\,
            in3 => \N__10436\,
            lcout => \SDATA1_ibuf_RNI098KZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__16269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15688\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19960\,
            ce => 'H',
            sr => \N__12110\
        );

    \counter_RNIE8FG_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__10949\,
            in1 => \N__16268\,
            in2 => \N__15756\,
            in3 => \N__15977\,
            lcout => OPEN,
            ltout => \N_35_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIT58K2_2_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__10437\,
            in1 => \_gnd_net_\,
            in2 => \N__10238\,
            in3 => \_gnd_net_\,
            lcout => \counter_RNIT58K2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_voltage_2_0__N_5_i_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111110"
        )
    port map (
            in0 => \N__13868\,
            in1 => \N__16212\,
            in2 => \N__15997\,
            in3 => \N__15664\,
            lcout => \un4_voltage_2_0__N_5_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_0_3_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10403\,
            in1 => \N__15205\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => un1_voltage_2_1_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNILOUG2_3_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10280\,
            in2 => \_gnd_net_\,
            in3 => \N__10433\,
            lcout => \counter_RNILOUG2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI2RBA2_3_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10435\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10947\,
            lcout => \counter_RNI2RBA2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_voltage_10_9__m3_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__10946\,
            in1 => \N__16406\,
            in2 => \N__15998\,
            in3 => \N__16273\,
            lcout => OPEN,
            ltout => \un4_voltage_10_9__N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNIKG123_1_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__10434\,
            in1 => \N__15684\,
            in2 => \N__10316\,
            in3 => \N__15146\,
            lcout => \voltage_2_RNIKG123Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATA1_ibuf_RNIFTO32_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19178\,
            in1 => \N__20217\,
            in2 => \_gnd_net_\,
            in3 => \N__16466\,
            lcout => voltage_0_1_sqmuxa,
            ltout => \voltage_0_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_0_cry_0_0_c_RNO_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10309\,
            in2 => \N__10298\,
            in3 => \_gnd_net_\,
            lcout => \un1_voltage_0_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_1_3_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101000100"
        )
    port map (
            in0 => \N__16400\,
            in1 => \N__15989\,
            in2 => \N__15813\,
            in3 => \N__16261\,
            lcout => \N_34_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNICVT22_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19181\,
            in2 => \_gnd_net_\,
            in3 => \N__16482\,
            lcout => un1_sclk17_9_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_0_3_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__16401\,
            in1 => \N__15988\,
            in2 => \N__15812\,
            in3 => \N__16260\,
            lcout => \N_41_i\,
            ltout => \N_41_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_1_1_cry_0_0_c_RNO_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10451\,
            in3 => \N__10432\,
            lcout => \un1_voltage_1_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_2_3_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20195\,
            in1 => \N__16265\,
            in2 => \N__16423\,
            in3 => \N__15750\,
            lcout => \ScreenBuffer_0_1_1_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_voltage_2_0__m11_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000100011000"
        )
    port map (
            in0 => \N__15990\,
            in1 => \N__15749\,
            in2 => \N__16284\,
            in3 => \N__16402\,
            lcout => \un4_voltage_2_0__i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12472\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_1_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCI1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10368\,
            in2 => \N__10478\,
            in3 => \N__10385\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI1OCIZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSH2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10382\,
            in2 => \N__10373\,
            in3 => \N__10376\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIVHSHZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI96513_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10372\,
            in2 => \N__10352\,
            in3 => \N__10343\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIZ0Z96513\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIVCO88_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11032\,
            in1 => \N__10340\,
            in2 => \N__10334\,
            in3 => \N__10319\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10487\,
            in2 => \_gnd_net_\,
            in3 => \N__10481\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGPZ0Z73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12473\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12689\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un1_beamylto9_0_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14824\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__un1_beamylto9Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un1_beamylto9_3_0_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__23284\,
            in1 => \N__14687\,
            in2 => \N__10469\,
            in3 => \N__20825\,
            lcout => \un113_pixel_4_0_15__un1_beamylto9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIID25_8_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14783\,
            in1 => \N__12973\,
            in2 => \N__14890\,
            in3 => \N__12882\,
            lcout => OPEN,
            ltout => \un5_visibley_axbxc7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_9_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001011010"
        )
    port map (
            in0 => \N__14973\,
            in1 => \N__14622\,
            in2 => \N__10466\,
            in3 => \N__11245\,
            lcout => chary_if_generate_plus_mult1_un33_sum_axb3,
            ltout => \chary_if_generate_plus_mult1_un33_sum_axb3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_1_tz_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__12477\,
            in1 => \N__12636\,
            in2 => \N__10463\,
            in3 => \N__18107\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_tz,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_6_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010100000"
        )
    port map (
            in0 => \N__12883\,
            in1 => \N__14623\,
            in2 => \N__12989\,
            in3 => \N__11246\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFS4T_0_7_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000010"
        )
    port map (
            in0 => \N__18108\,
            in1 => \N__14784\,
            in2 => \N__12768\,
            in3 => \N__18226\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un40_sum_ac0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_sx_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__11404\,
            in1 => \N__10505\,
            in2 => \N__10499\,
            in3 => \N__13996\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_sxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9425_0_6_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100110011001"
        )
    port map (
            in0 => \N__12977\,
            in1 => \N__12884\,
            in2 => \N__14659\,
            in3 => \N__20753\,
            lcout => OPEN,
            ltout => \beamY_RNI9425_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPOR8_0_6_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011010001"
        )
    port map (
            in0 => \N__12885\,
            in1 => \N__14418\,
            in2 => \N__10496\,
            in3 => \N__12978\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum,
            ltout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un47_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIL62O_0_7_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000001"
        )
    port map (
            in0 => \N__12453\,
            in1 => \N__12749\,
            in2 => \N__10493\,
            in3 => \N__14789\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_6_a2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_c4_d_0_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001110110111"
        )
    port map (
            in0 => \N__18222\,
            in1 => \N__12626\,
            in2 => \N__18139\,
            in3 => \N__13965\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_c4_d,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_8_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001000"
        )
    port map (
            in0 => \N__12625\,
            in1 => \N__18102\,
            in2 => \N__13997\,
            in3 => \N__18223\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIL62O_7_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__14790\,
            in1 => \N__12454\,
            in2 => \N__12761\,
            in3 => \N__12627\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_ac0_6_a1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__11263\,
            in1 => \N__18106\,
            in2 => \N__10490\,
            in3 => \N__18224\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_ac0_7_c_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_x0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000111"
        )
    port map (
            in0 => \N__18135\,
            in1 => \N__14785\,
            in2 => \N__12663\,
            in3 => \N__18254\,
            lcout => if_generate_plus_mult1_un61_sum_ac0_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9425_6_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__12979\,
            in1 => \N__12886\,
            in2 => \N__14660\,
            in3 => \N__20755\,
            lcout => OPEN,
            ltout => \beamY_RNI9425Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPOR8_6_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__12890\,
            in1 => \N__14420\,
            in2 => \N__10541\,
            in3 => \N__12980\,
            lcout => un5_visibley_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_x1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011011"
        )
    port map (
            in0 => \N__18253\,
            in1 => \N__18136\,
            in2 => \N__14810\,
            in3 => \N__12631\,
            lcout => if_generate_plus_mult1_un61_sum_ac0_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__20754\,
            in1 => \N__14419\,
            in2 => \N__12899\,
            in3 => \N__14630\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011010000001"
        )
    port map (
            in0 => \N__18255\,
            in1 => \N__12632\,
            in2 => \N__14028\,
            in3 => \N__18138\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010010010"
        )
    port map (
            in0 => \N__18137\,
            in1 => \N__18256\,
            in2 => \N__12664\,
            in3 => \N__14001\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_ns_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12745\,
            in1 => \N__10538\,
            in2 => \_gnd_net_\,
            in3 => \N__10532\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_ac0_6,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_ac0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI75QM4_5_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__12407\,
            in1 => \N__10520\,
            in2 => \N__10511\,
            in3 => \N__11526\,
            lcout => \beamY_RNI75QM4Z0Z_5\,
            ltout => \beamY_RNI75QM4Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_x1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__11527\,
            in1 => \N__12286\,
            in2 => \N__10508\,
            in3 => \N__10606\,
            lcout => OPEN,
            ltout => \if_generate_plus_mult1_un68_sum_axbxc5_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_ns_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10616\,
            in2 => \N__10610\,
            in3 => \N__11556\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11358\,
            in1 => \N__11336\,
            in2 => \_gnd_net_\,
            in3 => \N__11377\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_c4_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001101"
        )
    port map (
            in0 => \N__10607\,
            in1 => \N__13230\,
            in2 => \N__12455\,
            in3 => \N__10572\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_cZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101110"
        )
    port map (
            in0 => \N__13229\,
            in1 => \N__12408\,
            in2 => \_gnd_net_\,
            in3 => \N__14521\,
            lcout => OPEN,
            ltout => \if_generate_plus_mult1_un68_sum_ac0_7_1_0_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0_ns_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10583\,
            in2 => \N__10577\,
            in3 => \N__10571\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_ac0_7_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_1_2_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__11697\,
            in1 => \N__11980\,
            in2 => \N__10702\,
            in3 => \N__11678\,
            lcout => OPEN,
            ltout => \voltage_0_10_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17976\,
            in2 => \N__10553\,
            in3 => \N__10550\,
            lcout => \voltage_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19955\,
            ce => 'H',
            sr => \N__18542\
        );

    \voltage_1_RNO_1_2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11698\,
            in1 => \N__11656\,
            in2 => \N__10703\,
            in3 => \N__11679\,
            lcout => OPEN,
            ltout => \voltage_1_9_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_2_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__11859\,
            in1 => \N__15766\,
            in2 => \N__10544\,
            in3 => \N__10889\,
            lcout => \voltage_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19955\,
            ce => 'H',
            sr => \N__18542\
        );

    \counter_RNIVSBN2_0_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__15764\,
            in1 => \N__16285\,
            in2 => \_gnd_net_\,
            in3 => \N__11858\,
            lcout => un1_voltage_012_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_1_2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__11680\,
            in1 => \N__11699\,
            in2 => \N__11981\,
            in3 => \N__11933\,
            lcout => OPEN,
            ltout => \voltage_3_9_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_2_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111101001111"
        )
    port map (
            in0 => \N__15765\,
            in1 => \N__10652\,
            in2 => \N__10643\,
            in3 => \N__11860\,
            lcout => \voltage_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19955\,
            ce => 'H',
            sr => \N__18542\
        );

    \voltage_1_RNI359O_2_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16577\,
            in1 => \N__15245\,
            in2 => \_gnd_net_\,
            in3 => \N__15763\,
            lcout => \N_1509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_1_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__11914\,
            in1 => \N__11645\,
            in2 => \N__12043\,
            in3 => \N__10746\,
            lcout => voltage_2_9_iv_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIO70L4_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__10756\,
            in1 => \N__15512\,
            in2 => \N__16286\,
            in3 => \N__10727\,
            lcout => OPEN,
            ltout => \CO2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI8TL66_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000111100"
        )
    port map (
            in0 => \N__10778\,
            in1 => \N__10820\,
            in2 => \N__10640\,
            in3 => \N__16282\,
            lcout => \N_1155\,
            ltout => \N_1155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_0_3_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10799\,
            in1 => \N__10684\,
            in2 => \N__10637\,
            in3 => \N__11963\,
            lcout => voltage_0_10_iv_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_1_1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__11915\,
            in1 => \N__11774\,
            in2 => \N__11657\,
            in3 => \N__12003\,
            lcout => voltage_2_9_iv_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_1_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__10747\,
            in1 => \N__11961\,
            in2 => \N__10694\,
            in3 => \N__10628\,
            lcout => voltage_0_10_iv_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIO70L4_0_0_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001011010"
        )
    port map (
            in0 => \N__10726\,
            in1 => \N__10757\,
            in2 => \N__15519\,
            in3 => \N__16278\,
            lcout => \N_1154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNO_1_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11773\,
            in1 => \N__10683\,
            in2 => \N__12005\,
            in3 => \N__11962\,
            lcout => voltage_0_10_iv_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_1_3_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__10714\,
            in1 => \N__11643\,
            in2 => \N__10695\,
            in3 => \N__10794\,
            lcout => voltage_1_9_iv_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_1_3_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__10795\,
            in1 => \N__11913\,
            in2 => \N__11975\,
            in3 => \N__10715\,
            lcout => voltage_3_9_iv_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_1_0_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__10748\,
            in1 => \N__10685\,
            in2 => \N__12042\,
            in3 => \N__11644\,
            lcout => voltage_1_9_iv_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNICMA33_0_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__13118\,
            in1 => \N__12031\,
            in2 => \N__16283\,
            in3 => \N__11726\,
            lcout => \CO1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI2ACM1_1_0_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19309\,
            in1 => \N__15742\,
            in2 => \N__13348\,
            in3 => \N__16256\,
            lcout => voltage_2_1_sqmuxa,
            ltout => \voltage_2_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_1_3_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10793\,
            in1 => \N__11912\,
            in2 => \N__10718\,
            in3 => \N__10713\,
            lcout => voltage_2_9_iv_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI2ACM1_2_0_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19308\,
            in1 => \N__15741\,
            in2 => \N__13347\,
            in3 => \N__16255\,
            lcout => voltage_1_1_sqmuxa,
            ltout => \voltage_1_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_1_1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__11642\,
            in1 => \N__12004\,
            in2 => \N__10841\,
            in3 => \N__11771\,
            lcout => voltage_1_9_iv_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_3_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101010101"
        )
    port map (
            in0 => \N__10838\,
            in1 => \N__11863\,
            in2 => \N__15733\,
            in3 => \N__10874\,
            lcout => \voltage_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19961\,
            ce => 'H',
            sr => \N__18544\
        );

    \voltage_1_RNI579O_3_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19449\,
            in1 => \N__15162\,
            in2 => \_gnd_net_\,
            in3 => \N__15641\,
            lcout => \N_1510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100111011"
        )
    port map (
            in0 => \N__10832\,
            in1 => \N__10826\,
            in2 => \N__15734\,
            in3 => \N__11864\,
            lcout => \voltage_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19961\,
            ce => 'H',
            sr => \N__18544\
        );

    \voltage_0_RNI313M_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15642\,
            in1 => \N__15209\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => OPEN,
            ltout => \N_1506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIGLLH1_0_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10816\,
            in2 => \N__10805\,
            in3 => \N__16243\,
            lcout => \counter_RNIGLLH1Z0Z_0\,
            ltout => \counter_RNIGLLH1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI4K0L4_0_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100101"
        )
    port map (
            in0 => \N__11591\,
            in1 => \_gnd_net_\,
            in2 => \N__10802\,
            in3 => \N__11772\,
            lcout => \N_2063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_RNI313M_0_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19419\,
            in1 => \_gnd_net_\,
            in2 => \N__15219\,
            in3 => \N__15643\,
            lcout => \N_1522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_1_1_cry_0_0_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15339\,
            in2 => \N__10769\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => un1_voltage_1_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_0_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15104\,
            in2 => \N__10907\,
            in3 => \N__10898\,
            lcout => \voltage_1_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => un1_voltage_1_1_cry_0,
            carryout => un1_voltage_1_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_0_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10895\,
            in2 => \N__15262\,
            in3 => \N__10880\,
            lcout => \voltage_1_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => un1_voltage_1_1_cry_1,
            carryout => un1_voltage_1_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNO_0_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10877\,
            lcout => \voltage_1_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIJTI6_2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__15936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15721\,
            lcout => \Z_decfrac4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI1SFG_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__13863\,
            in1 => \N__13771\,
            in2 => \N__16399\,
            in3 => \N__13643\,
            lcout => OPEN,
            ltout => \un6_slaveselectlto9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIS6CQ_2_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__15937\,
            in1 => \N__16267\,
            in2 => \N__10868\,
            in3 => \N__15722\,
            lcout => OPEN,
            ltout => \un6_slaveselect_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIHC2O1_2_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__13625\,
            in1 => \_gnd_net_\,
            in2 => \N__10865\,
            in3 => \N__10862\,
            lcout => un5_slaveselect,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_2_1_cry_0_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15395\,
            in2 => \N__13100\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => un1_voltage_2_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_0_1_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15142\,
            in2 => \N__10856\,
            in3 => \N__10844\,
            lcout => \voltage_2_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => un1_voltage_2_1_cry_0,
            carryout => un1_voltage_2_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_0_2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10979\,
            in2 => \N__15305\,
            in3 => \N__10973\,
            lcout => \voltage_2_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => un1_voltage_2_1_cry_1,
            carryout => un1_voltage_2_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100101111"
        )
    port map (
            in0 => \N__10970\,
            in1 => \N__13421\,
            in2 => \N__10964\,
            in3 => \N__10952\,
            lcout => \voltage_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19966\,
            ce => 'H',
            sr => \N__18547\
        );

    \counter_RNIJTI6_3_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__16257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16408\,
            lcout => \N_46_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_3_RNO_0_0_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__16410\,
            in1 => \N__15992\,
            in2 => \N__15816\,
            in3 => \N__16259\,
            lcout => OPEN,
            ltout => \un1_sclk17_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_3_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20194\,
            in1 => \N__20062\,
            in2 => \N__10928\,
            in3 => \N__23647\,
            lcout => \ScreenBuffer_0_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_10_RNO_0_0_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16409\,
            in1 => \N__15991\,
            in2 => \N__15815\,
            in3 => \N__16258\,
            lcout => OPEN,
            ltout => \un1_sclk17_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_10_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20193\,
            in1 => \N__20061\,
            in2 => \N__10925\,
            in3 => \N__23707\,
            lcout => \ScreenBuffer_0_10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13276\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_1_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3Q404_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11034\,
            in2 => \N__10922\,
            in3 => \N__10910\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI3QZ0Z404\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40I45_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11036\,
            in2 => \N__11093\,
            in3 => \N__11081\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI40IZ0Z45\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3S246_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11035\,
            in2 => \N__11078\,
            in3 => \N__11066\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3SZ0Z246\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIRSJ6F_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11188\,
            in1 => \N__11009\,
            in2 => \N__11063\,
            in3 => \N__11051\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11048\,
            in2 => \_gnd_net_\,
            in3 => \N__11039\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7JZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIOGP73_0_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11033\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12555\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_2_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIV79_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11183\,
            in2 => \N__11282\,
            in3 => \N__11003\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITIVZ0Z79\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80D_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11000\,
            in2 => \N__11189\,
            in3 => \N__10994\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI2G80DZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4E_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11187\,
            in2 => \N__10991\,
            in3 => \N__10982\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI4OM4EZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIK4SNU_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11121\,
            in1 => \N__11165\,
            in2 => \N__11210\,
            in3 => \N__11201\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJF_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11198\,
            in2 => \_gnd_net_\,
            in3 => \N__11192\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGEJJFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDA7J8_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11182\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12172\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11122\,
            in2 => \N__11291\,
            in3 => \N__11159\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTFZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUO_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11120\,
            in2 => \N__11156\,
            in3 => \N__11147\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNITLMUOZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NS_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11123\,
            in2 => \N__11144\,
            in3 => \N__11135\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3L0NSZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11099\,
            in2 => \N__11132\,
            in3 => \N__11119\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RU_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11300\,
            in2 => \_gnd_net_\,
            in3 => \N__11294\,
            lcout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI7V2RUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12556\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13262\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEDF31_6_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14037\,
            in1 => \N__12690\,
            in2 => \N__12485\,
            in3 => \N__18291\,
            lcout => \beamY_RNIEDF31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__12176\,
            in1 => \N__21871\,
            in2 => \_gnd_net_\,
            in3 => \N__20832\,
            lcout => \beamY_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6EUJ1_7_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__18261\,
            in1 => \N__11270\,
            in2 => \N__11414\,
            in3 => \N__14020\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c4_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m1_5_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100101"
        )
    port map (
            in0 => \N__12687\,
            in1 => \N__18140\,
            in2 => \N__14036\,
            in3 => \N__18260\,
            lcout => if_m1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_0_6_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__13001\,
            in1 => \N__12911\,
            in2 => \N__14701\,
            in3 => \N__11252\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_ac0_6_a6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4QBV1_6_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__14021\,
            in1 => \N__12323\,
            in2 => \N__11222\,
            in3 => \N__18141\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_c4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILILV4_8_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__18142\,
            in1 => \N__11219\,
            in2 => \N__11213\,
            in3 => \N__11423\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_c4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEG4HI_3_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__11393\,
            in1 => \N__13310\,
            in2 => \N__11417\,
            in3 => \N__13231\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIER061_6_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__12719\,
            in1 => \N__18262\,
            in2 => \N__18169\,
            in3 => \N__11413\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIED3U1_0_7_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__12677\,
            in1 => \N__12721\,
            in2 => \N__11315\,
            in3 => \N__14035\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14441\,
            in2 => \_gnd_net_\,
            in3 => \N__20790\,
            lcout => chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum,
            ltout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un68_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_ac0_5_x0_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11334\,
            in1 => \N__11359\,
            in2 => \N__11387\,
            in3 => \N__11383\,
            lcout => if_generate_plus_mult1_un75_sum_ac0_5_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_ac0_5_x1_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__11384\,
            in1 => \N__12544\,
            in2 => \N__11363\,
            in3 => \N__11335\,
            lcout => if_generate_plus_mult1_un75_sum_ac0_5_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFS4T_7_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__18163\,
            in1 => \N__14812\,
            in2 => \N__12776\,
            in3 => \N__18285\,
            lcout => \beamY_RNIFS4TZ0Z_7\,
            ltout => \beamY_RNIFS4TZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIED3U1_7_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101111011010"
        )
    port map (
            in0 => \N__12720\,
            in1 => \N__14033\,
            in2 => \N__11306\,
            in3 => \N__12676\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un47_sum_axbxc5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQTGS2_8_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101111000"
        )
    port map (
            in0 => \N__18164\,
            in1 => \N__14034\,
            in2 => \N__11303\,
            in3 => \N__18286\,
            lcout => \beamY_RNIQTGS2Z0Z_8\,
            ltout => \beamY_RNIQTGS2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPNEA3_6_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12481\,
            in2 => \N__11474\,
            in3 => \N__12678\,
            lcout => chary_if_generate_plus_mult1_un54_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIO8DB4_6_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__12471\,
            in1 => \N__11455\,
            in2 => \N__12575\,
            in3 => \N__12692\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc5_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIECMV4_5_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11449\,
            in1 => \N__11464\,
            in2 => \_gnd_net_\,
            in3 => \N__12469\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axb3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0JK7C_5_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__12567\,
            in1 => \N__11450\,
            in2 => \N__11471\,
            in3 => \N__11434\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb3,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axb3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIS0VDC_3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__13270\,
            in1 => \_gnd_net_\,
            in2 => \N__11468\,
            in3 => \N__12545\,
            lcout => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_1_0_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14476\,
            in2 => \_gnd_net_\,
            in3 => \N__20831\,
            lcout => un5_visibley_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPNEA3_0_6_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__12691\,
            in1 => \_gnd_net_\,
            in2 => \N__11456\,
            in3 => \N__12470\,
            lcout => \beamY_RNIPNEA3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0K169_6_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101001"
        )
    port map (
            in0 => \N__11465\,
            in1 => \N__11454\,
            in2 => \N__12574\,
            in3 => \N__11435\,
            lcout => \beamY_RNI0K169Z0Z_6\,
            ltout => \beamY_RNI0K169Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV42D31_0_6_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101001"
        )
    port map (
            in0 => \N__12520\,
            in1 => \N__13070\,
            in2 => \N__11426\,
            in3 => \N__13046\,
            lcout => \beamY_RNIV42D31_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g1_0_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20841\,
            in2 => \_gnd_net_\,
            in3 => \N__14479\,
            lcout => \un113_pixel_3_0_11__g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_5_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101100011010"
        )
    port map (
            in0 => \N__13309\,
            in1 => \N__12818\,
            in2 => \N__13277\,
            in3 => \N__11573\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un68_sum_c5_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_3_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12819\,
            in1 => \N__13159\,
            in2 => \N__11567\,
            in3 => \N__14481\,
            lcout => \un113_pixel_3_0_11__N_4_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m1_x1_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12298\,
            in1 => \N__11540\,
            in2 => \N__14298\,
            in3 => \N__14689\,
            lcout => OPEN,
            ltout => \if_m1_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m1_ns_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__11504\,
            in1 => \_gnd_net_\,
            in2 => \N__11564\,
            in3 => \N__11561\,
            lcout => if_m1_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m1_x0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12297\,
            in1 => \N__11539\,
            in2 => \N__14297\,
            in3 => \N__14688\,
            lcout => if_m1_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_7_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__13158\,
            in1 => \N__13308\,
            in2 => \_gnd_net_\,
            in3 => \N__14480\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un75_sum_c5_N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_2_0_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__11498\,
            in1 => \N__12820\,
            in2 => \N__11492\,
            in3 => \N__14690\,
            lcout => g1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19993\,
            lcout => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIKUA33_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11587\,
            in2 => \_gnd_net_\,
            in3 => \N__11765\,
            lcout => \N_1159_i\,
            ltout => \N_1159_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_1_2_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__11684\,
            in1 => \N__11932\,
            in2 => \N__11660\,
            in3 => \N__11655\,
            lcout => voltage_2_9_iv_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNIO5RB1_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19292\,
            in2 => \_gnd_net_\,
            in3 => \N__13562\,
            lcout => voltage_0_0_sqmuxa_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_4_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11600\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_ScreenBuffer_1_1_1_sqmuxa_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__13556\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__17185\,
            lcout => \slaveselect_RNILOQC2Z0Z_1\,
            ltout => \slaveselect_RNILOQC2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_4_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19288\,
            in2 => \N__11594\,
            in3 => \N__17149\,
            lcout => \ScreenBuffer_1_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNICHLH1_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16213\,
            in1 => \N__15521\,
            in2 => \_gnd_net_\,
            in3 => \N__15533\,
            lcout => \counter_RNICHLH1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNIQDU22_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001011100"
        )
    port map (
            in0 => \N__13557\,
            in1 => \N__18568\,
            in2 => \N__19328\,
            in3 => \_gnd_net_\,
            lcout => un1_counter_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNIE1PG2_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__13336\,
            in1 => \N__13555\,
            in2 => \_gnd_net_\,
            in3 => \N__19284\,
            lcout => un1_voltage_012_0,
            ltout => \un1_voltage_012_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIVSBN2_0_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__16214\,
            in1 => \_gnd_net_\,
            in2 => \N__12047\,
            in3 => \N__15862\,
            lcout => un1_voltage_012_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNICMA33_0_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011111011000"
        )
    port map (
            in0 => \N__16248\,
            in1 => \N__13117\,
            in2 => \N__11725\,
            in3 => \N__12044\,
            lcout => \N_1153\,
            ltout => \N_1153_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_RNO_1_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__11976\,
            in1 => \N__11761\,
            in2 => \N__11936\,
            in3 => \N__11931\,
            lcout => OPEN,
            ltout => \voltage_3_9_iv_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_3_1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111101001111"
        )
    port map (
            in0 => \N__15821\,
            in1 => \N__11882\,
            in2 => \N__11867\,
            in3 => \N__11840\,
            lcout => \voltage_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19964\,
            ce => 'H',
            sr => \N__18545\
        );

    \voltage_1_1_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__11839\,
            in1 => \N__11807\,
            in2 => \N__11798\,
            in3 => \N__15822\,
            lcout => \voltage_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19964\,
            ce => 'H',
            sr => \N__18545\
        );

    \voltage_0_RNIVS2M_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15820\,
            in1 => \N__15127\,
            in2 => \_gnd_net_\,
            in3 => \N__19051\,
            lcout => \N_1504\,
            ltout => \N_1504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_1_c_RNO_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16246\,
            in2 => \N__11783\,
            in3 => \N__11714\,
            lcout => \un42_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI8DLH1_0_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16247\,
            in1 => \_gnd_net_\,
            in2 => \N__11724\,
            in3 => \N__11780\,
            lcout => \counter_RNI8DLH1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_1_RNI139O_1_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19352\,
            in1 => \N__15086\,
            in2 => \_gnd_net_\,
            in3 => \N__15819\,
            lcout => \N_1508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_3_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12064\,
            lcout => \un1_ScreenBuffer_1_0_1_sqmuxa_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_4_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__19291\,
            in1 => \N__12065\,
            in2 => \_gnd_net_\,
            in3 => \N__16954\,
            lcout => \ScreenBuffer_1_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19967\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16181\,
            in1 => \N__16347\,
            in2 => \_gnd_net_\,
            in3 => \N__13517\,
            lcout => \Z_decfrac4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIE36D_0_5_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13855\,
            in1 => \N__16346\,
            in2 => \N__15974\,
            in3 => \N__13764\,
            lcout => voltage_011_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_2_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__13478\,
            in1 => \N__19290\,
            in2 => \_gnd_net_\,
            in3 => \N__13553\,
            lcout => \slaveselect_RNILOQC2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_cry_1_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15810\,
            in2 => \N__16242\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15935\,
            in2 => \_gnd_net_\,
            in3 => \N__12056\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => counter_cry_1,
            carryout => counter_cry_2,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16393\,
            in2 => \_gnd_net_\,
            in3 => \N__12053\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => counter_cry_2,
            carryout => counter_cry_3,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_4_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13862\,
            in2 => \_gnd_net_\,
            in3 => \N__12050\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => counter_cry_3,
            carryout => counter_cry_4,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_5_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13767\,
            in2 => \_gnd_net_\,
            in3 => \N__12125\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => counter_cry_4,
            carryout => counter_cry_5,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_6_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13795\,
            in2 => \_gnd_net_\,
            in3 => \N__12122\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => counter_cry_5,
            carryout => counter_cry_6,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_7_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13898\,
            in2 => \_gnd_net_\,
            in3 => \N__12119\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => counter_cry_6,
            carryout => counter_cry_7,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_8_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13720\,
            in2 => \_gnd_net_\,
            in3 => \N__12116\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => counter_cry_7,
            carryout => counter_cry_8,
            clk => \N__19970\,
            ce => 'H',
            sr => \N__12102\
        );

    \counter_9_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13924\,
            in2 => \_gnd_net_\,
            in3 => \N__12113\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19973\,
            ce => 'H',
            sr => \N__12109\
        );

    \counter_0_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16150\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19973\,
            ce => 'H',
            sr => \N__12109\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22611\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2579_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12073\,
            in2 => \N__14048\,
            in3 => \N__12080\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIZ0Z2579\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTAS4_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14071\,
            in2 => \N__13658\,
            in3 => \N__12077\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIVTASZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14070\,
            in1 => \N__12074\,
            in2 => \N__14096\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKP36_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14084\,
            in2 => \_gnd_net_\,
            in3 => \N__12245\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNISKPZ0Z36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un173_pixellto5_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010100001000"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__23088\,
            in2 => \N__22622\,
            in3 => \N__12242\,
            lcout => chessboardpixel_un173_pixellt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un151_pixel_if_generate_plus_mult1_remainder_0_6_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__12241\,
            in1 => \N__12233\,
            in2 => \N__22621\,
            in3 => \N__12226\,
            lcout => chessboardpixel_un151_pixel_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un177_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5DMTF_0_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12193\,
            lcout => OPEN,
            ltout => \chessboardpixel_un177_pixel_if_generate_plus_mult1_un1_rem_adjust_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un177_pixel_if_generate_plus_mult1_remainder_0_5_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100110101010"
        )
    port map (
            in0 => \N__12218\,
            in1 => \N__12185\,
            in2 => \N__12212\,
            in3 => \N__12151\,
            lcout => OPEN,
            ltout => \chessboardpixel_un177_pixel_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un174_pixel_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011110"
        )
    port map (
            in0 => \N__12209\,
            in1 => \N__12203\,
            in2 => \N__12197\,
            in3 => \N__12131\,
            lcout => chessboardpixel_un174_pixel,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_1_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101001000000"
        )
    port map (
            in0 => \N__12194\,
            in1 => \N__12173\,
            in2 => \N__12152\,
            in3 => \N__12184\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__chessboardpixel_un199_pixellto4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__chessboardpixel_un199_pixellto4_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__12174\,
            in1 => \N__12150\,
            in2 => \N__12134\,
            in3 => \N__23231\,
            lcout => chessboardpixel_un199_pixellt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSyncZ0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__14207\,
            in1 => \N__14991\,
            in2 => \N__14930\,
            in3 => \N__12347\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_a3_0_3_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__23264\,
            in1 => \N__14838\,
            in2 => \_gnd_net_\,
            in3 => \N__20840\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__g0_i_a3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_a3_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14495\,
            in1 => \N__12314\,
            in2 => \N__12326\,
            in3 => \N__13013\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII8O41_9_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__12478\,
            in1 => \N__18158\,
            in2 => \N__12722\,
            in3 => \N__18287\,
            lcout => \beamY_RNII8O41Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_a3_0_4_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14696\,
            in1 => \N__14925\,
            in2 => \N__12929\,
            in3 => \N__14990\,
            lcout => \un113_pixel_4_0_15__g0_i_a3_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001010101010"
        )
    port map (
            in0 => \N__23265\,
            in1 => \N__14125\,
            in2 => \N__24639\,
            in3 => \N__17519\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111010011"
        )
    port map (
            in0 => \N__12668\,
            in1 => \N__18162\,
            in2 => \N__14039\,
            in3 => \N__18284\,
            lcout => if_generate_plus_mult1_un54_sum_axbxc5,
            ltout => \if_generate_plus_mult1_un54_sum_axbxc5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m4_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010010101"
        )
    port map (
            in0 => \N__13263\,
            in1 => \N__12308\,
            in2 => \N__12302\,
            in3 => \N__12299\,
            lcout => OPEN,
            ltout => \row_1_if_i2_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_ac0_5_ns_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12260\,
            in2 => \N__12254\,
            in3 => \N__12251\,
            lcout => row_1_if_generate_plus_mult1_un75_sum_ac0_5,
            ltout => \row_1_if_generate_plus_mult1_un75_sum_ac0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_c5_x0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000101100100"
        )
    port map (
            in0 => \N__13264\,
            in1 => \N__14299\,
            in2 => \N__12779\,
            in3 => \N__12479\,
            lcout => if_generate_plus_mult1_un75_sum_c5_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x1_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12480\,
            in1 => \N__13265\,
            in2 => \N__14310\,
            in3 => \N__12501\,
            lcout => if_generate_plus_mult1_un82_sum_axbxc5_0_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un5_beamx_4_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13011\,
            in2 => \_gnd_net_\,
            in3 => \N__12921\,
            lcout => un1_beamy_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJNLC_9_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110111010101"
        )
    port map (
            in0 => \N__14989\,
            in1 => \N__14892\,
            in2 => \N__12775\,
            in3 => \N__14811\,
            lcout => \beamY_RNIJNLCZ0Z_9\,
            ltout => \beamY_RNIJNLCZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVGU01_9_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14032\,
            in2 => \N__12695\,
            in3 => \N__12669\,
            lcout => \beamY_RNIVGU01Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIR51RF1_3_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110111010"
        )
    port map (
            in0 => \N__13307\,
            in1 => \N__12817\,
            in2 => \N__12557\,
            in3 => \N__13269\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV42D31_6_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100011110"
        )
    port map (
            in0 => \N__13069\,
            in1 => \N__13055\,
            in2 => \N__12521\,
            in3 => \N__13045\,
            lcout => \beamY_RNIV42D31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_x0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110011001"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__14303\,
            in2 => \N__12506\,
            in3 => \N__13266\,
            lcout => if_generate_plus_mult1_un82_sum_axbxc5_0_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_c5_x1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__13267\,
            in1 => \N__12505\,
            in2 => \N__14311\,
            in3 => \N__12468\,
            lcout => OPEN,
            ltout => \if_generate_plus_mult1_un75_sum_c5_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_c5_ns_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__13082\,
            in1 => \N__14186\,
            in2 => \N__13073\,
            in3 => \_gnd_net_\,
            lcout => row_1_if_generate_plus_mult1_un75_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7SK1V_3_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__13054\,
            in2 => \_gnd_net_\,
            in3 => \N__13044\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axbxc5_0,
            ltout => \chary_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDHF0F2_3_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111010110100"
        )
    port map (
            in0 => \N__13025\,
            in1 => \N__13174\,
            in2 => \N__13016\,
            in3 => \N__13268\,
            lcout => chary_if_generate_plus_mult1_un75_sum_axbxc5_m6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_beamylto6_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14695\,
            in1 => \N__13012\,
            in2 => \N__12928\,
            in3 => \N__14371\,
            lcout => un4_beamylt8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0VHAB1_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__14471\,
            in1 => \N__13156\,
            in2 => \_gnd_net_\,
            in3 => \N__13305\,
            lcout => \chary_if_generate_plus_mult1_un75_sum_c5_N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPLAE31_4_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__12813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14694\,
            lcout => OPEN,
            ltout => \beamY_RNIPLAE31Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4TRT4_3_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001110101100"
        )
    port map (
            in0 => \N__14372\,
            in1 => \N__12836\,
            in2 => \N__12830\,
            in3 => \N__12827\,
            lcout => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVGVF22_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__13157\,
            in1 => \_gnd_net_\,
            in2 => \N__12821\,
            in3 => \N__14472\,
            lcout => chary_if_generate_plus_mult1_un1_sum_axbxc3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000011000"
        )
    port map (
            in0 => \N__13133\,
            in1 => \N__12791\,
            in2 => \N__20858\,
            in3 => \N__12785\,
            lcout => \un113_pixel_3_0_11__g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_1_3_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14470\,
            in2 => \_gnd_net_\,
            in3 => \N__20826\,
            lcout => un4_beamylt6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__20827\,
            in1 => \N__13271\,
            in2 => \N__14487\,
            in3 => \N__13306\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un75_sum_axbxc5_N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_0_x2_0_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001110101100"
        )
    port map (
            in0 => \N__13272\,
            in1 => \N__13175\,
            in2 => \N__13163\,
            in3 => \N__13160\,
            lcout => \un113_pixel_3_0_11__g0_0_x2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15344\,
            in1 => \N__15379\,
            in2 => \_gnd_net_\,
            in3 => \N__19305\,
            lcout => \ScreenBuffer_1_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19963\,
            ce => \N__13127\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_2_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19303\,
            in1 => \N__15261\,
            in2 => \_gnd_net_\,
            in3 => \N__15294\,
            lcout => \ScreenBuffer_1_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19963\,
            ce => \N__13127\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15224\,
            in1 => \N__19304\,
            in2 => \_gnd_net_\,
            in3 => \N__15176\,
            lcout => \ScreenBuffer_1_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19963\,
            ce => \N__13127\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_1_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19302\,
            in1 => \N__15129\,
            in2 => \_gnd_net_\,
            in3 => \N__15100\,
            lcout => \ScreenBuffer_1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19963\,
            ce => \N__13127\,
            sr => \_gnd_net_\
        );

    \voltage_0_RNIVS2M_0_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15128\,
            in1 => \N__19047\,
            in2 => \_gnd_net_\,
            in3 => \N__15836\,
            lcout => \N_1520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_voltage_2_1_cry_0_c_RNO_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20218\,
            in1 => \N__19280\,
            in2 => \N__15389\,
            in3 => \N__13468\,
            lcout => \un1_voltage_2_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_RNO_0_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13469\,
            in1 => \N__20219\,
            in2 => \N__19327\,
            in3 => \N__15375\,
            lcout => OPEN,
            ltout => \un1_voltage_2_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_2_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13451\,
            in2 => \N__13442\,
            in3 => \N__13412\,
            lcout => \voltage_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19965\,
            ce => 'H',
            sr => \N__18546\
        );

    \voltage_2_2_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__13414\,
            in1 => \N__13439\,
            in2 => \_gnd_net_\,
            in3 => \N__13433\,
            lcout => \voltage_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19965\,
            ce => 'H',
            sr => \N__18546\
        );

    \voltage_2_1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__13413\,
            in1 => \N__13397\,
            in2 => \_gnd_net_\,
            in3 => \N__13388\,
            lcout => \voltage_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19965\,
            ce => 'H',
            sr => \N__18546\
        );

    \voltage_0_RNI1V2M_2_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15286\,
            in1 => \N__16555\,
            in2 => \_gnd_net_\,
            in3 => \N__15817\,
            lcout => \N_1505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_1_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13376\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => un42_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_2_c_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21912\,
            in2 => \N__15485\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un42_cry_1,
            carryout => un42_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_3_c_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13370\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un42_cry_2,
            carryout => un42_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_3_c_RNIMRT41_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13358\,
            in1 => \N__13598\,
            in2 => \_gnd_net_\,
            in3 => \N__13352\,
            lcout => voltage_011,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__19306\,
            in1 => \N__15458\,
            in2 => \_gnd_net_\,
            in3 => \N__17332\,
            lcout => \ScreenBuffer_1_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_2_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__20205\,
            in1 => \N__13487\,
            in2 => \N__17210\,
            in3 => \N__19307\,
            lcout => \ScreenBuffer_0_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__19289\,
            in1 => \N__13486\,
            in2 => \_gnd_net_\,
            in3 => \N__13561\,
            lcout => \slaveselect_RNILOQCZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIE36D_5_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13859\,
            in1 => \N__16360\,
            in2 => \N__15975\,
            in3 => \N__13765\,
            lcout => \ScreenBuffer_1_122_1\,
            ltout => \ScreenBuffer_1_122_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNITIV01_0_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13594\,
            in1 => \N__16216\,
            in2 => \N__13490\,
            in3 => \N__15832\,
            lcout => \ScreenBuffer_1_3_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNITIV01_2_0_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16215\,
            in1 => \N__13612\,
            in2 => \N__15854\,
            in3 => \N__13596\,
            lcout => \ScreenBuffer_1_0_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_1_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__19301\,
            in1 => \N__13571\,
            in2 => \N__16979\,
            in3 => \N__20203\,
            lcout => \ScreenBuffer_0_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNITIV01_1_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__16217\,
            in1 => \N__13611\,
            in2 => \N__15855\,
            in3 => \N__13595\,
            lcout => \ScreenBuffer_1_1_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_4_RNO_0_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19300\,
            in2 => \_gnd_net_\,
            in3 => \N__13467\,
            lcout => OPEN,
            ltout => \un1_sclk17_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_4_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__18958\,
            in1 => \N__16498\,
            in2 => \N__13646\,
            in3 => \N__20204\,
            lcout => \ScreenBuffer_0_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIUJ6D_9_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13922\,
            in1 => \N__13718\,
            in2 => \_gnd_net_\,
            in3 => \N__13642\,
            lcout => un39_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIT7J6_6_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13895\,
            in2 => \_gnd_net_\,
            in3 => \N__13793\,
            lcout => un39_0_3,
            ltout => \un39_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIB6GG_9_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13921\,
            in1 => \N__13717\,
            in2 => \N__13628\,
            in3 => \N__13763\,
            lcout => un5_slaveselect_1,
            ltout => \un5_slaveselect_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNITIV01_4_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__13874\,
            in1 => \_gnd_net_\,
            in2 => \N__13616\,
            in3 => \N__13860\,
            lcout => un10_slaveselect,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNITIV01_0_0_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__13613\,
            in1 => \N__13597\,
            in2 => \N__16241\,
            in3 => \N__15818\,
            lcout => \ScreenBuffer_1_2_1_sqmuxa\,
            ltout => \ScreenBuffer_1_2_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_0_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19329\,
            in2 => \N__13565\,
            in3 => \N__13554\,
            lcout => \slaveselect_RNILOQC2Z0Z_0\,
            ltout => \slaveselect_RNILOQC2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_5_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13520\,
            in3 => \_gnd_net_\,
            lcout => \un1_ScreenBuffer_1_2_1_sqmuxa_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIAAPJ_7_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13516\,
            in1 => \N__13811\,
            in2 => \N__13928\,
            in3 => \N__13896\,
            lcout => slaveselect_1lto9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIEUS9_6_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13923\,
            in1 => \N__13897\,
            in2 => \_gnd_net_\,
            in3 => \N__13794\,
            lcout => OPEN,
            ltout => \un1_counter_1lto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI283N_8_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13810\,
            in1 => \N__13719\,
            in2 => \N__13877\,
            in3 => \N__13766\,
            lcout => un1_counter_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_6_0_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__16520\,
            in1 => \N__16507\,
            in2 => \N__18940\,
            in3 => \N__20199\,
            lcout => \ScreenBuffer_0_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19977\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_2_3_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16344\,
            in1 => \N__15923\,
            in2 => \N__15861\,
            in3 => \N__16109\,
            lcout => un10_slaveselectlt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIN1J6_4_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13861\,
            in2 => \_gnd_net_\,
            in3 => \N__16345\,
            lcout => un1_counter_1lt9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIBRS9_6_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13799\,
            in1 => \N__13772\,
            in2 => \_gnd_net_\,
            in3 => \N__13724\,
            lcout => slaveselect_1lto9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNIIRSC1_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__13694\,
            in1 => \N__13685\,
            in2 => \N__19997\,
            in3 => \N__19330\,
            lcout => \SCLK1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22462\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJE1_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14056\,
            in2 => \N__16610\,
            in3 => \N__13649\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9KJEZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LB2_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16630\,
            in2 => \N__16667\,
            in3 => \N__14087\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF6LBZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGAHS5_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14072\,
            in1 => \N__14057\,
            in2 => \N__16655\,
            in3 => \N__14078\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3H63_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16643\,
            in2 => \_gnd_net_\,
            in3 => \N__14075\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIC3HZ0Z63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_0_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16629\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22459\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17529\,
            in2 => \_gnd_net_\,
            in3 => \N__18698\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un5_beamx_2_0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23232\,
            in1 => \N__15002\,
            in2 => \_gnd_net_\,
            in3 => \N__14837\,
            lcout => \un113_pixel_4_0_15__un5_beamx_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_row_2_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001110000"
        )
    port map (
            in0 => \N__14038\,
            in1 => \N__18168\,
            in2 => \N__18041\,
            in3 => \N__18292\,
            lcout => \un113_pixel_4_0_15__un4_rowZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un5_beamx_4_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14700\,
            in1 => \N__14494\,
            in2 => \N__14929\,
            in3 => \N__20883\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__un5_beamxZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un5_beamx_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14156\,
            in1 => \N__24593\,
            in2 => \N__14150\,
            in3 => \N__14203\,
            lcout => un5_beamx_0,
            ltout => \un5_beamx_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010110101010"
        )
    port map (
            in0 => \N__24594\,
            in1 => \_gnd_net_\,
            in2 => \N__14111\,
            in3 => \N__17533\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un3_beamx_5_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17867\,
            in1 => \N__17902\,
            in2 => \N__17790\,
            in3 => \N__17466\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__un3_beamxZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un3_beamx_7_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__17830\,
            in1 => \N__18704\,
            in2 => \N__14108\,
            in3 => \N__17686\,
            lcout => \un113_pixel_4_0_15__un3_beamxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un13_beamylto3_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__17866\,
            in1 => \N__17901\,
            in2 => \N__18720\,
            in3 => \N__17829\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un13_beamylto10_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__14105\,
            in1 => \N__17614\,
            in2 => \N__17687\,
            in3 => \N__16805\,
            lcout => un13_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un13_beamylto5_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14335\,
            in1 => \N__17726\,
            in2 => \_gnd_net_\,
            in3 => \N__17783\,
            lcout => un13_beamylt6_0,
            ltout => \un13_beamylt6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_6_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__17684\,
            in1 => \N__17615\,
            in2 => \N__14099\,
            in3 => \N__16806\,
            lcout => un13_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un18_beamylto9_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__14336\,
            in1 => \N__17727\,
            in2 => \N__17792\,
            in3 => \N__16841\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_row_5_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14327\,
            in1 => \N__14321\,
            in2 => \N__14315\,
            in3 => \N__20576\,
            lcout => \un113_pixel_4_0_15__un4_rowZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un3_beamx_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16807\,
            in1 => \N__14249\,
            in2 => \N__17621\,
            in3 => \N__17728\,
            lcout => un3_beamx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un1_beamxlto6_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17729\,
            in1 => \N__17685\,
            in2 => \N__17791\,
            in3 => \N__17834\,
            lcout => OPEN,
            ltout => \un1_beamxlt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSyncZ0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__16808\,
            in1 => \N__17619\,
            in2 => \N__14243\,
            in3 => \N__17467\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un15_beamy_2_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14714\,
            in1 => \N__17468\,
            in2 => \N__14552\,
            in3 => \N__14225\,
            lcout => \un113_pixel_4_0_15__un15_beamyZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_0_ns_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14184\,
            in1 => \N__14219\,
            in2 => \_gnd_net_\,
            in3 => \N__14213\,
            lcout => row_1_if_generate_plus_mult1_un82_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un8_beamylto9_1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14983\,
            in1 => \N__14920\,
            in2 => \N__14845\,
            in3 => \N__14202\,
            lcout => \un113_pixel_4_0_15__un8_beamylto9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_row_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14185\,
            in1 => \N__23615\,
            in2 => \N__14165\,
            in3 => \N__23108\,
            lcout => un4_row,
            ltout => \un4_row_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_5_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15023\,
            in1 => \N__15014\,
            in2 => \N__15005\,
            in3 => \N__16937\,
            lcout => \Pixel_3_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_beamylto9_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__14998\,
            in1 => \N__14921\,
            in2 => \N__14846\,
            in3 => \N__14720\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un8_beamylto9_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__14708\,
            in1 => \N__20886\,
            in2 => \N__14702\,
            in3 => \N__14478\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_a9_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100100001"
        )
    port map (
            in0 => \N__20888\,
            in1 => \N__23244\,
            in2 => \N__14540\,
            in3 => \N__20677\,
            lcout => \N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_x4_0_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20966\,
            lcout => \N_6_i\,
            ltout => \N_6_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_a9_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__20887\,
            in1 => \N__23243\,
            in2 => \N__14531\,
            in3 => \N__20676\,
            lcout => \N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m2_2_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__17251\,
            in1 => \N__14528\,
            in2 => \_gnd_net_\,
            in3 => \N__14477\,
            lcout => OPEN,
            ltout => \if_m2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010001011"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__14354\,
            in2 => \N__14345\,
            in3 => \N__14342\,
            lcout => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16876\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PA3_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16793\,
            in2 => \_gnd_net_\,
            in3 => \N__15056\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI707PAZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PA3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16904\,
            in2 => \N__21888\,
            in3 => \N__15053\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI828PAZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16888\,
            in2 => \_gnd_net_\,
            in3 => \N__15050\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15047\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_0_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17077\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBS1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15419\,
            in2 => \N__15044\,
            in3 => \N__15035\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNINNKBSZ0Z1\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5B3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15032\,
            in2 => \N__15410\,
            in3 => \N__15026\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIHMC5BZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15434\,
            in2 => \N__15443\,
            in3 => \N__15405\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5B3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15409\,
            in1 => \N__15428\,
            in2 => \N__16898\,
            in3 => \N__15422\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNILUG5BZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15418\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_5_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111101"
        )
    port map (
            in0 => \N__17073\,
            in1 => \N__20996\,
            in2 => \N__18736\,
            in3 => \N__17117\,
            lcout => \un113_pixel_4_0_15__g0_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_e_0_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19319\,
            in1 => \N__15380\,
            in2 => \_gnd_net_\,
            in3 => \N__15343\,
            lcout => \ScreenBuffer_1_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19972\,
            ce => \N__15068\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_e_0_2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15293\,
            in1 => \N__19322\,
            in2 => \_gnd_net_\,
            in3 => \N__15263\,
            lcout => \ScreenBuffer_1_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19972\,
            ce => \N__15068\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_e_0_3_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19320\,
            in1 => \N__15223\,
            in2 => \_gnd_net_\,
            in3 => \N__15175\,
            lcout => \ScreenBuffer_1_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19972\,
            ce => \N__15068\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_e_0_1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__19321\,
            in2 => \_gnd_net_\,
            in3 => \N__15099\,
            lcout => \ScreenBuffer_1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19972\,
            ce => \N__15068\,
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_15_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__17078\,
            in1 => \N__21159\,
            in2 => \_gnd_net_\,
            in3 => \N__17118\,
            lcout => font_un3_pixel_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un42_cry_2_c_RNO_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15532\,
            in1 => \N__16245\,
            in2 => \_gnd_net_\,
            in3 => \N__15520\,
            lcout => \un42_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_11_RNO_0_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__16274\,
            in1 => \N__15980\,
            in2 => \N__16426\,
            in3 => \N__19249\,
            lcout => OPEN,
            ltout => \un1_sclk17_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_11_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16511\,
            in1 => \N__20207\,
            in2 => \N__15473\,
            in3 => \N__23686\,
            lcout => \ScreenBuffer_0_11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_12_RNO_0_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16275\,
            in1 => \N__15981\,
            in2 => \N__16427\,
            in3 => \N__19250\,
            lcout => OPEN,
            ltout => \un1_sclk17_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_12_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16512\,
            in1 => \N__20208\,
            in2 => \N__15470\,
            in3 => \N__18973\,
            lcout => \ScreenBuffer_0_12Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATA1_ibuf_RNI800F_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20206\,
            in1 => \N__19248\,
            in2 => \_gnd_net_\,
            in3 => \N__15978\,
            lcout => \ScreenBuffer_0_0_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNILOQC2_6_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15457\,
            lcout => \un1_ScreenBuffer_1_3_1_sqmuxa_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_5_RNO_0_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16276\,
            in1 => \N__15979\,
            in2 => \N__15863\,
            in3 => \N__19251\,
            lcout => OPEN,
            ltout => \un1_sclk17_8_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_5_0_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16513\,
            in1 => \N__20209\,
            in2 => \N__15446\,
            in3 => \N__19525\,
            lcout => \ScreenBuffer_0_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_e_0_2_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19334\,
            in1 => \N__16592\,
            in2 => \_gnd_net_\,
            in3 => \N__16559\,
            lcout => \ScreenBuffer_1_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19978\,
            ce => \N__18430\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_6_RNO_0_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16222\,
            in1 => \N__15994\,
            in2 => \N__15856\,
            in3 => \N__19331\,
            lcout => un1_sclk17_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_0_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__16499\,
            in1 => \N__15539\,
            in2 => \N__19547\,
            in3 => \N__20162\,
            lcout => \ScreenBuffer_0_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATAZ0Z2_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__20161\,
            in1 => \N__16441\,
            in2 => \N__16514\,
            in3 => \N__19332\,
            lcout => \SDATA2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_8_RNO_0_0_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15995\,
            in1 => \N__15841\,
            in2 => \N__16425\,
            in3 => \N__16223\,
            lcout => OPEN,
            ltout => \un1_sclk17_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_8_0_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20163\,
            in1 => \N__20074\,
            in2 => \N__16430\,
            in3 => \N__17020\,
            lcout => \ScreenBuffer_0_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_9_RNO_0_0_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15993\,
            in1 => \N__15837\,
            in2 => \N__16424\,
            in3 => \N__16221\,
            lcout => un1_sclk17_5_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNO_0_0_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16266\,
            in1 => \N__15996\,
            in2 => \N__15857\,
            in3 => \N__19333\,
            lcout => un1_sclk17_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_0_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19715\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22731\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3V_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16673\,
            in2 => \N__16601\,
            in3 => \N__16658\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0K3VZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKID91_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19718\,
            in2 => \N__19775\,
            in3 => \N__16646\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKIDZ0Z91\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIU1G53_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16631\,
            in1 => \N__16616\,
            in2 => \N__19757\,
            in3 => \N__16637\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIB1_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19736\,
            in2 => \_gnd_net_\,
            in3 => \N__16634\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI3LIBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30T_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19717\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ30TZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22732\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22253\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17900\,
            in2 => \_gnd_net_\,
            in3 => \N__18699\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22305\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18299\,
            in2 => \_gnd_net_\,
            in3 => \N__16694\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16682\,
            in2 => \N__21851\,
            in3 => \N__16691\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22004\,
            in2 => \_gnd_net_\,
            in3 => \N__16688\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16685\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22003\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__ANC4_0_i_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__22005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22140\,
            lcout => \N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__N_32_i_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22255\,
            in2 => \_gnd_net_\,
            in3 => \N__22309\,
            lcout => \N_32_i\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16748\,
            in2 => \N__19792\,
            in3 => \N__16676\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16738\,
            in2 => \N__16784\,
            in3 => \N__16775\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16834\,
            in1 => \N__16724\,
            in2 => \N__16772\,
            in3 => \N__16763\,
            lcout => charx_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16739\,
            in1 => \N__22020\,
            in2 => \N__16760\,
            in3 => \N__16751\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16747\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\,
            ltout => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16727\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un26_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22256\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22743\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16816\,
            in2 => \N__16718\,
            in3 => \N__16709\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16835\,
            in2 => \N__16706\,
            in3 => \N__16697\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__16817\,
            in2 => \N__16862\,
            in3 => \N__16853\,
            lcout => charx_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16850\,
            in2 => \_gnd_net_\,
            in3 => \N__16844\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un18_beamylto9_2_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18367\,
            in1 => \N__17680\,
            in2 => \N__17620\,
            in3 => \N__18334\,
            lcout => \un113_pixel_4_0_15__un18_beamylto9Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16833\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17069\,
            in2 => \_gnd_net_\,
            in3 => \N__17120\,
            lcout => g1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un3_beamx_2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18335\,
            in2 => \_gnd_net_\,
            in3 => \N__18368\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101001110101"
        )
    port map (
            in0 => \N__18614\,
            in1 => \N__24349\,
            in2 => \N__18406\,
            in3 => \N__18381\,
            lcout => charx_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI80GJR1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__24354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18617\,
            lcout => charx_if_generate_plus_mult1_un1_sum_axb1,
            ltout => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNITU0P65_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16787\,
            in3 => \N__17119\,
            lcout => font_un3_pixel_28,
            ltout => \font_un3_pixel_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un61_pixel_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18814\,
            in1 => \N__21623\,
            in2 => \N__16940\,
            in3 => \N__18724\,
            lcout => OPEN,
            ltout => \font_un61_pixel_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un125_pixel_m_6_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16936\,
            in1 => \N__16925\,
            in2 => \N__16913\,
            in3 => \N__16910\,
            lcout => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011001010101"
        )
    port map (
            in0 => \N__18382\,
            in1 => \N__18402\,
            in2 => \N__24358\,
            in3 => \N__18615\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIJT9MA3_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010110001010"
        )
    port map (
            in0 => \N__18616\,
            in1 => \N__24353\,
            in2 => \N__18407\,
            in3 => \N__18383\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIE3GVR1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__24348\,
            in1 => \N__18398\,
            in2 => \_gnd_net_\,
            in3 => \N__18613\,
            lcout => charx_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIKML437_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__17065\,
            in1 => \N__21157\,
            in2 => \_gnd_net_\,
            in3 => \N__17113\,
            lcout => font_un3_pixel_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNI5D2AEA_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011000110"
        )
    port map (
            in0 => \N__17114\,
            in1 => \N__16868\,
            in2 => \N__21163\,
            in3 => \N__17066\,
            lcout => font_un3_pixel_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9A68G8_0_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000011000"
        )
    port map (
            in0 => \N__20934\,
            in1 => \N__20678\,
            in2 => \N__20893\,
            in3 => \N__20981\,
            lcout => font_un28_pixel_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFBK6ED_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__23285\,
            in1 => \N__18838\,
            in2 => \N__20690\,
            in3 => \N__20882\,
            lcout => font_un67_pixel_ac0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__17068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17116\,
            lcout => \un113_pixel_4_0_15__gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_x2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__17115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17067\,
            lcout => OPEN,
            ltout => \N_9_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__18725\,
            in1 => \N__21158\,
            in2 => \N__17033\,
            in3 => \N__17030\,
            lcout => \un113_pixel_4_0_15__g0_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_6_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20935\,
            lcout => \un113_pixel_7_1_7__g0_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_8_RNIV2FB2F_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001111011"
        )
    port map (
            in0 => \N__23510\,
            in1 => \N__25958\,
            in2 => \N__23603\,
            in3 => \N__17024\,
            lcout => OPEN,
            ltout => \currentchar_1_9_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_RNIBIJQMK_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__25960\,
            in1 => \N__17006\,
            in2 => \N__16997\,
            in3 => \N__17164\,
            lcout => \ScreenBuffer_1_0_e_0_RNIBIJQMKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_9_RNI06IC2F_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001111011"
        )
    port map (
            in0 => \N__23511\,
            in1 => \N__25959\,
            in2 => \N__23604\,
            in3 => \N__20018\,
            lcout => OPEN,
            ltout => \currentchar_1_6_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_RNIEVE0NK_0_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__25961\,
            in1 => \N__16994\,
            in2 => \N__16982\,
            in3 => \N__16978\,
            lcout => \ScreenBuffer_1_1_e_0_RNIEVE0NKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_RNISJ0D2F_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110100101"
        )
    port map (
            in0 => \N__23512\,
            in1 => \N__25962\,
            in2 => \N__23605\,
            in3 => \N__16958\,
            lcout => OPEN,
            ltout => \ScreenBuffer_1_0_RNISJ0D2FZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_RNIQ3KT7J1_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100101010001"
        )
    port map (
            in0 => \N__17132\,
            in1 => \N__25539\,
            in2 => \N__17285\,
            in3 => \N__17126\,
            lcout => OPEN,
            ltout => \ScreenBuffer_1_0_RNIQ3KT7J1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_RNIVUON9Q2_4_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22984\,
            in2 => \N__17282\,
            in3 => \N__25396\,
            lcout => currentchar_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17237\,
            in1 => \N__17279\,
            in2 => \N__17264\,
            in3 => \N__23513\,
            lcout => un3_rowlto0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17278\,
            in1 => \N__17260\,
            in2 => \_gnd_net_\,
            in3 => \N__17236\,
            lcout => un3_rowlto1,
            ltout => \un3_rowlto1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_e_0_RNINV7VE9_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__17219\,
            in2 => \N__17213\,
            in3 => \N__17206\,
            lcout => \ScreenBuffer_1_2_e_0_RNINV7VE9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_0_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__19326\,
            in1 => \N__17189\,
            in2 => \N__17168\,
            in3 => \N__20210\,
            lcout => \ScreenBuffer_0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_RNITM3E2F_4_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110100101"
        )
    port map (
            in0 => \N__23503\,
            in1 => \N__25985\,
            in2 => \N__23607\,
            in3 => \N__17153\,
            lcout => OPEN,
            ltout => \ScreenBuffer_1_1_RNITM3E2FZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_RNI4PNO0E3_4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__25545\,
            in1 => \N__17315\,
            in2 => \N__17135\,
            in3 => \N__25740\,
            lcout => currentchar_1_11_ns_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_RNIUP6F2F_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110100101"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__25986\,
            in2 => \N__23608\,
            in3 => \N__17390\,
            lcout => \ScreenBuffer_1_2_RNIUP6F2FZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_0_1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24130\,
            in1 => \N__17300\,
            in2 => \_gnd_net_\,
            in3 => \N__17291\,
            lcout => \N_4566_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_RNIVS9G2F_4_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110100101"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__25984\,
            in2 => \N__23606\,
            in3 => \N__17333\,
            lcout => \ScreenBuffer_1_3_RNIVS9G2FZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \g1_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23585\,
            in2 => \_gnd_net_\,
            in3 => \N__23528\,
            lcout => OPEN,
            ltout => \g1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_22_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19385\,
            in1 => \N__25546\,
            in2 => \N__17309\,
            in3 => \N__19379\,
            lcout => OPEN,
            ltout => \N_1428_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g1_1_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__25395\,
            in1 => \N__23870\,
            in2 => \N__17306\,
            in3 => \N__23972\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_21_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011101100"
        )
    port map (
            in0 => \N__24514\,
            in1 => \N__24777\,
            in2 => \N__17303\,
            in3 => \N__17339\,
            lcout => \N_1300_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_24_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25136\,
            in1 => \N__25028\,
            in2 => \_gnd_net_\,
            in3 => \N__24513\,
            lcout => OPEN,
            ltout => \un112_pixel_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_1_2_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__25029\,
            in1 => \N__24776\,
            in2 => \N__17294\,
            in3 => \N__25211\,
            lcout => \N_1293_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m10_0_x1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__25991\,
            in1 => \N__25405\,
            in2 => \N__23030\,
            in3 => \N__21526\,
            lcout => m10_0_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_2_4_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__19318\,
            in1 => \N__17399\,
            in2 => \_gnd_net_\,
            in3 => \N__17389\,
            lcout => \ScreenBuffer_1_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_1_2_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001011110"
        )
    port map (
            in0 => \N__25738\,
            in1 => \N__17375\,
            in2 => \N__25538\,
            in3 => \N__17369\,
            lcout => OPEN,
            ltout => \un113_pixel_3_0_11__currentchar_1_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_1_4_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25403\,
            in1 => \N__25989\,
            in2 => \N__17354\,
            in3 => \N__22874\,
            lcout => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2\,
            ltout => \un113_pixel_3_0_11__currentchar_1_4Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un112_pixel_1_2_x1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001111"
        )
    port map (
            in0 => \N__25990\,
            in1 => \N__22994\,
            in2 => \N__17351\,
            in3 => \N__25404\,
            lcout => un112_pixel_1_2_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m10_0_ns_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__21527\,
            in1 => \N__17348\,
            in2 => \N__23018\,
            in3 => \N__19511\,
            lcout => un112_pixel_2_2,
            ltout => \un112_pixel_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIHMH43T2_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111000"
        )
    port map (
            in0 => \N__23433\,
            in1 => \N__25007\,
            in2 => \N__17342\,
            in3 => \N__24504\,
            lcout => \ScreenBuffer_0_7_RNIHMH43T2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_0_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__21528\,
            in1 => \N__23015\,
            in2 => \N__25068\,
            in3 => \N__23886\,
            lcout => \un113_pixel_3_0_11__g0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_4_am_7_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__23421\,
            in1 => \N__25017\,
            in2 => \_gnd_net_\,
            in3 => \N__24476\,
            lcout => un115_pixel_4_am_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDQUNU91_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__24477\,
            in1 => \N__25026\,
            in2 => \N__24860\,
            in3 => \N__23424\,
            lcout => OPEN,
            ltout => \beamY_RNIDQUNU91Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7RM4IF_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__17429\,
            in1 => \_gnd_net_\,
            in2 => \N__17423\,
            in3 => \N__24138\,
            lcout => \beamY_RNI7RM4IFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC0GLNQ_0_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__25016\,
            in1 => \N__23423\,
            in2 => \N__24861\,
            in3 => \N__25133\,
            lcout => OPEN,
            ltout => \un115_pixel_2_sn_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPQEDM42_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17414\,
            in2 => \N__17420\,
            in3 => \N__24479\,
            lcout => \beamY_RNIPQEDM42Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un112_pixel_7_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24478\,
            in1 => \N__25027\,
            in2 => \_gnd_net_\,
            in3 => \N__25134\,
            lcout => OPEN,
            ltout => \un112_pixel_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_1_4_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__24760\,
            in1 => \N__25018\,
            in2 => \N__17417\,
            in3 => \N__25207\,
            lcout => \N_1293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIINK7J73_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__25015\,
            in1 => \N__24759\,
            in2 => \_gnd_net_\,
            in3 => \N__23422\,
            lcout => \beamY_RNIINK7J73Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17903\,
            in2 => \N__18742\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17859\,
            in2 => \_gnd_net_\,
            in3 => \N__17408\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17828\,
            in2 => \_gnd_net_\,
            in3 => \N__17405\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__17762\,
            in2 => \_gnd_net_\,
            in3 => \N__17402\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17712\,
            in2 => \_gnd_net_\,
            in3 => \N__17561\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17661\,
            in2 => \_gnd_net_\,
            in3 => \N__17558\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17596\,
            in2 => \_gnd_net_\,
            in3 => \N__17555\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18359\,
            in2 => \_gnd_net_\,
            in3 => \N__17552\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__21062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18326\,
            in2 => \_gnd_net_\,
            in3 => \N__17549\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__21061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17462\,
            in1 => \N__17540\,
            in2 => \_gnd_net_\,
            in3 => \N__17471\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__22141\,
            in1 => \N__22254\,
            in2 => \_gnd_net_\,
            in3 => \N__22072\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22143\,
            lcout => if_generate_plus_mult1_un47_sum_0_cry_3_ma,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__N_1184_0_i_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22147\,
            in2 => \_gnd_net_\,
            in3 => \N__22075\,
            lcout => \N_1184_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111011000"
        )
    port map (
            in0 => \N__22073\,
            in1 => \N__22142\,
            in2 => \N__22157\,
            in3 => \N__22188\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18700\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17891\,
            in2 => \_gnd_net_\,
            in3 => \N__17870\,
            lcout => charx_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17860\,
            in2 => \_gnd_net_\,
            in3 => \N__17837\,
            lcout => charx_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17819\,
            in2 => \N__21870\,
            in3 => \N__17795\,
            lcout => chessboardpixel_un151_pixel_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17763\,
            in2 => \_gnd_net_\,
            in3 => \N__17732\,
            lcout => charx_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17713\,
            in2 => \_gnd_net_\,
            in3 => \N__17690\,
            lcout => charx_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21844\,
            in2 => \N__17679\,
            in3 => \N__17624\,
            lcout => charx_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17597\,
            in2 => \_gnd_net_\,
            in3 => \N__17564\,
            lcout => charx_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18360\,
            in2 => \N__21900\,
            in3 => \N__18338\,
            lcout => \un5_visiblex_cry_7_c_RNIVZ0Z952\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18327\,
            in2 => \_gnd_net_\,
            in3 => \N__18305\,
            lcout => \CO3_0\,
            ltout => \CO3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18302\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un26_sum_s_2_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un4_row_1_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__18293\,
            in1 => \N__18170\,
            in2 => \N__18050\,
            in3 => \N__20348\,
            lcout => \un113_pixel_4_0_15__un4_rowZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22310\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \voltage_0_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__18026\,
            in1 => \N__18008\,
            in2 => \_gnd_net_\,
            in3 => \N__17990\,
            lcout => \voltage_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19980\,
            ce => 'H',
            sr => \N__18548\
        );

    \voltage_0_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__17989\,
            in1 => \N__17957\,
            in2 => \_gnd_net_\,
            in3 => \N__17945\,
            lcout => \voltage_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19980\,
            ce => 'H',
            sr => \N__18548\
        );

    \nCS1_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__18578\,
            in1 => \N__19113\,
            in2 => \_gnd_net_\,
            in3 => \N__17914\,
            lcout => \nCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19980\,
            ce => 'H',
            sr => \N__18548\
        );

    \slaveselect_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__19114\,
            in1 => \N__18577\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \slaveselectZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19980\,
            ce => 'H',
            sr => \N__18548\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22817\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_e_0_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19110\,
            in1 => \N__18518\,
            in2 => \_gnd_net_\,
            in3 => \N__18456\,
            lcout => \ScreenBuffer_1_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19976\,
            ce => \N__18434\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_e_0_3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19111\,
            in1 => \N__19463\,
            in2 => \_gnd_net_\,
            in3 => \N__19433\,
            lcout => \ScreenBuffer_1_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19976\,
            ce => \N__18434\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_e_0_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19030\,
            in1 => \N__19373\,
            in2 => \_gnd_net_\,
            in3 => \N__19112\,
            lcout => \ScreenBuffer_1_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19976\,
            ce => \N__18434\,
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22769\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24347\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18628\,
            in2 => \N__18599\,
            in3 => \N__18386\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPME1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20381\,
            in2 => \N__20441\,
            in3 => \N__18371\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI5QPMEZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18629\,
            in2 => \N__20420\,
            in3 => \N__20379\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHR1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20399\,
            in2 => \_gnd_net_\,
            in3 => \N__18620\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNINBIHRZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22665\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23080\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20473\,
            in2 => \N__18851\,
            in3 => \N__18590\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25871\,
            in2 => \N__20588\,
            in3 => \N__18587\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25310\,
            in1 => \N__20474\,
            in2 => \N__20537\,
            in3 => \N__18584\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20495\,
            in2 => \_gnd_net_\,
            in3 => \N__18581\,
            lcout => column_1_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9A68G8_2_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101100110"
        )
    port map (
            in0 => \N__20983\,
            in1 => \N__20933\,
            in2 => \N__20894\,
            in3 => \N__20672\,
            lcout => chary_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_i_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22619\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFBK6ED_0_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100001"
        )
    port map (
            in0 => \N__20689\,
            in1 => \N__23300\,
            in2 => \N__18842\,
            in3 => \N__20892\,
            lcout => font_un64_pixel_ac0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_0_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21625\,
            in1 => \N__18740\,
            in2 => \N__18827\,
            in3 => \N__18637\,
            lcout => \un113_pixel_4_0_15__g0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un57_pixel_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18815\,
            in1 => \N__21624\,
            in2 => \N__18743\,
            in3 => \N__21289\,
            lcout => OPEN,
            ltout => \font_un57_pixel_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un125_pixel_m_6_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18803\,
            in2 => \N__18797\,
            in3 => \N__18794\,
            lcout => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3\,
            ltout => \un113_pixel_4_0_15__font_un125_pixel_m_6Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un125_pixel_m_6_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18788\,
            in1 => \N__18779\,
            in2 => \N__18773\,
            in3 => \N__21258\,
            lcout => \un113_pixel_4_0_15__font_un125_pixel_mZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21259\,
            in1 => \N__18770\,
            in2 => \N__18758\,
            in3 => \N__21235\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__g0_iZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_1_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__23348\,
            in1 => \N__18905\,
            in2 => \N__18746\,
            in3 => \N__21587\,
            lcout => g0_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__Pixel_6_iv_a3_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18741\,
            in2 => \_gnd_net_\,
            in3 => \N__18638\,
            lcout => \un113_pixel_4_0_15__Pixel_6_iv_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un112_pixel_7_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21325\,
            in1 => \N__25360\,
            in2 => \_gnd_net_\,
            in3 => \N__25585\,
            lcout => un112_pixel_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIOEPPEK1_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__25364\,
            in1 => \_gnd_net_\,
            in2 => \N__24852\,
            in3 => \N__21324\,
            lcout => OPEN,
            ltout => \beamY_RNIOEPPEK1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1G38U63_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__23879\,
            in1 => \N__23998\,
            in2 => \N__18920\,
            in3 => \N__24542\,
            lcout => OPEN,
            ltout => \N_3461_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_19_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__24800\,
            in1 => \N__18917\,
            in2 => \N__18911\,
            in3 => \N__23443\,
            lcout => OPEN,
            ltout => \N_4568_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_18_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__21443\,
            in1 => \_gnd_net_\,
            in2 => \N__18908\,
            in3 => \N__24168\,
            lcout => \N_1305_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__18899\,
            in1 => \N__24242\,
            in2 => \N__23349\,
            in3 => \N__19808\,
            lcout => OPEN,
            ltout => \N_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__18893\,
            in1 => \N__18881\,
            in2 => \N__18875\,
            in3 => \N__21206\,
            lcout => \un113_pixel_4_0_15__g0_i_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un71_pixellto5_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__23999\,
            in1 => \N__21326\,
            in2 => \N__25399\,
            in3 => \N__23880\,
            lcout => font_un71_pixellt7_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_m7_0_m3_ns_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__25736\,
            in1 => \N__18872\,
            in2 => \N__25540\,
            in3 => \N__18863\,
            lcout => OPEN,
            ltout => \un113_pixel_3_0_11__currentchar_m7_0_m3_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_m7_0_m3_ns_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__25525\,
            in1 => \N__19478\,
            in2 => \N__19469\,
            in3 => \N__19391\,
            lcout => \un113_pixel_3_0_11__currentchar_N_13\,
            ltout => \un113_pixel_3_0_11__currentchar_N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_m7_0_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__25937\,
            in1 => \_gnd_net_\,
            in2 => \N__19466\,
            in3 => \N__25394\,
            lcout => \un113_pixel_3_0_11__currentchar_m7_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19462\,
            in1 => \N__19177\,
            in2 => \_gnd_net_\,
            in3 => \N__19432\,
            lcout => \ScreenBuffer_1_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19979\,
            ce => \N__18998\,
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_1_0_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25739\,
            in1 => \N__21404\,
            in2 => \N__25988\,
            in3 => \N__21386\,
            lcout => \un113_pixel_4_0_15__g0_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_3_0_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25737\,
            in1 => \N__21437\,
            in2 => \N__25972\,
            in3 => \N__21422\,
            lcout => \un113_pixel_4_0_15__g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19368\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__19046\,
            lcout => \ScreenBuffer_1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19979\,
            ce => \N__18998\,
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_12_RNIE3Q33F_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__18974\,
            in2 => \N__23016\,
            in3 => \N__18959\,
            lcout => OPEN,
            ltout => \ScreenBuffer_0_12_RNIE3Q33FZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_6_RNIVTBDB12_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__25735\,
            in1 => \N__22990\,
            in2 => \N__18944\,
            in3 => \N__18941\,
            lcout => \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0\,
            ltout => \ScreenBuffer_0_6_RNIVTBDB12Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNII0GVLQ_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25541\,
            in2 => \N__19553\,
            in3 => \N__25246\,
            lcout => \ScreenBuffer_0_7_RNII0GVLQZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_m7_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__25386\,
            in1 => \N__25971\,
            in2 => \N__22986\,
            in3 => \N__19503\,
            lcout => currentchar_m7_0,
            ltout => \currentchar_m7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25387\,
            in1 => \N__19598\,
            in2 => \N__19550\,
            in3 => \N__25586\,
            lcout => \un113_pixel_4_0_15__N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIN5F98I1_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25734\,
            in1 => \N__19546\,
            in2 => \N__22985\,
            in3 => \N__19526\,
            lcout => \ScreenBuffer_0_7_RNIN5F98I1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__un115_pixel_5_bm_7_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__24484\,
            in1 => \N__23425\,
            in2 => \_gnd_net_\,
            in3 => \N__25141\,
            lcout => un115_pixel_5_bm_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIHMH43T2_0_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111011101"
        )
    port map (
            in0 => \N__25140\,
            in1 => \N__25006\,
            in2 => \N__23439\,
            in3 => \N__24483\,
            lcout => \ScreenBuffer_0_7_RNIHMH43T2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_1_12_1_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__25406\,
            in1 => \N__21359\,
            in2 => \N__25547\,
            in3 => \N__21341\,
            lcout => currentchar_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un112_pixel_1_2_ns_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__19510\,
            in1 => \N__21523\,
            in2 => \N__23031\,
            in3 => \N__19487\,
            lcout => un112_pixel_2_8,
            ltout => \un112_pixel_2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__m8_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19600\,
            in1 => \N__25417\,
            in2 => \N__19481\,
            in3 => \N__25591\,
            lcout => \un113_pixel_7_1_7__N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_1_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23019\,
            in2 => \_gnd_net_\,
            in3 => \N__21524\,
            lcout => currentchar_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_4_ns_7_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23322\,
            in1 => \N__19610\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => OPEN,
            ltout => \N_1287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_6_ns_7_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__24154\,
            in1 => \_gnd_net_\,
            in2 => \N__19616\,
            in3 => \N__21539\,
            lcout => \N_1289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIR2AGB22_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19599\,
            in1 => \N__25418\,
            in2 => \_gnd_net_\,
            in3 => \N__25590\,
            lcout => currentchar_1_0,
            ltout => \currentchar_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__m10_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010100000"
        )
    port map (
            in0 => \N__23791\,
            in1 => \N__23020\,
            in2 => \N__19613\,
            in3 => \N__21525\,
            lcout => \un113_pixel_7_1_7__N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_4_bm_7_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__23958\,
            in1 => \N__25021\,
            in2 => \N__23881\,
            in3 => \N__24480\,
            lcout => un115_pixel_4_bm_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__m21_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__25135\,
            in1 => \N__19604\,
            in2 => \N__25416\,
            in3 => \N__25592\,
            lcout => \un113_pixel_1_0_3__N_10_mux\,
            ltout => \un113_pixel_1_0_3__N_10_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_9_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__23852\,
            in1 => \N__24153\,
            in2 => \N__19580\,
            in3 => \N__19658\,
            lcout => OPEN,
            ltout => \N_1285_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_i_m2_0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011010001"
        )
    port map (
            in0 => \N__19559\,
            in1 => \N__23346\,
            in2 => \N__19577\,
            in3 => \N__19574\,
            lcout => \N_1286_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__m14_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__23959\,
            in1 => \N__25019\,
            in2 => \N__23882\,
            in3 => \N__24481\,
            lcout => m14,
            ltout => \m14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICJUESD2_1_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__25020\,
            in1 => \N__24837\,
            in2 => \N__19667\,
            in3 => \N__25205\,
            lcout => \beamY_RNICJUESD2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_4_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25206\,
            in1 => \N__25025\,
            in2 => \N__21014\,
            in3 => \N__19664\,
            lcout => \N_1327_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g0_6_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__24482\,
            in1 => \N__23017\,
            in2 => \N__25069\,
            in3 => \N__21529\,
            lcout => \un113_pixel_3_0_11__g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_3_5_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24169\,
            in1 => \N__19652\,
            in2 => \_gnd_net_\,
            in3 => \N__19646\,
            lcout => OPEN,
            ltout => \N_1306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23347\,
            in2 => \N__19640\,
            in3 => \N__19637\,
            lcout => \N_4561_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m11_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__25145\,
            in1 => \N__25065\,
            in2 => \_gnd_net_\,
            in3 => \N__24525\,
            lcout => OPEN,
            ltout => \m11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_5_ns_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24838\,
            in2 => \N__19631\,
            in3 => \N__19628\,
            lcout => \N_1322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m16_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__23987\,
            in1 => \N__25064\,
            in2 => \N__23883\,
            in3 => \N__24524\,
            lcout => \un113_pixel_4_0_15__N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_6_bm_2_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25067\,
            in1 => \N__21650\,
            in2 => \N__24862\,
            in3 => \N__21944\,
            lcout => OPEN,
            ltout => \un115_pixel_6_bm_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_6_ns_2_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24170\,
            in1 => \_gnd_net_\,
            in2 => \N__19811\,
            in3 => \N__19799\,
            lcout => \N_1330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_6_am_2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__25066\,
            in1 => \N__24839\,
            in2 => \_gnd_net_\,
            in3 => \N__25214\,
            lcout => un115_pixel_6_am_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__SUM4_3_i_a2_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22257\,
            in2 => \_gnd_net_\,
            in3 => \N__22319\,
            lcout => \N_56\,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DC_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19793\,
            in2 => \N__21746\,
            in3 => \N__19760\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIG3DCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDE_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21926\,
            in2 => \N__19682\,
            in3 => \N__19739\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRTDEZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS72T_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19716\,
            in1 => \N__19688\,
            in2 => \N__21776\,
            in3 => \N__19724\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IE_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19681\,
            in1 => \N__21761\,
            in2 => \N__22094\,
            in3 => \N__19721\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIV5IEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19677\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBR12_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21742\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIBRZ0Z12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22720\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19871\,
            in2 => \N__19832\,
            in3 => \N__19865\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19862\,
            in2 => \N__19856\,
            in3 => \N__19847\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19844\,
            in2 => \N__20234\,
            in3 => \N__19838\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19835\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_2_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22251\,
            lcout => un5_visiblex_i_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_2110_i_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__22023\,
            in1 => \N__22271\,
            in2 => \_gnd_net_\,
            in3 => \N__19820\,
            lcout => \N_2110_i\,
            ltout => \N_2110_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19823\,
            in3 => \N__20246\,
            lcout => if_generate_plus_mult1_un54_sum_axb_2_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_m_5_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22022\,
            in1 => \N__22270\,
            in2 => \_gnd_net_\,
            in3 => \N__19819\,
            lcout => if_generate_plus_mult1_un47_sum_m_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100101101100"
        )
    port map (
            in0 => \N__22067\,
            in1 => \N__20337\,
            in2 => \N__22745\,
            in3 => \N__22730\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101001011"
        )
    port map (
            in0 => \N__22024\,
            in1 => \N__22373\,
            in2 => \N__20349\,
            in3 => \N__20240\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111111010"
        )
    port map (
            in0 => \N__22252\,
            in1 => \N__22162\,
            in2 => \N__22320\,
            in3 => \N__22021\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22025\,
            in1 => \N__20225\,
            in2 => \N__20350\,
            in3 => \N__22385\,
            lcout => if_generate_plus_mult1_un54_sum_axb_3_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_9_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20216\,
            in1 => \N__20084\,
            in2 => \N__20039\,
            in3 => \N__20011\,
            lcout => \ScreenBuffer_0_9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19983\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20278\,
            in2 => \_gnd_net_\,
            in3 => \N__19886\,
            lcout => if_generate_plus_mult1_un54_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111000011"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__20344\,
            in2 => \N__22349\,
            in3 => \N__22032\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22449\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20363\,
            in2 => \N__20290\,
            in3 => \N__20354\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20351\,
            in2 => \N__20312\,
            in3 => \N__20300\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20565\,
            in1 => \N__20297\,
            in2 => \N__20291\,
            in3 => \N__20267\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_s_5_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20264\,
            in2 => \_gnd_net_\,
            in3 => \N__20258\,
            lcout => if_generate_plus_mult1_un54_sum_s_5,
            ltout => \if_generate_plus_mult1_un54_sum_s_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20255\,
            in3 => \_gnd_net_\,
            lcout => column_1_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22492\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23081\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PU8_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20464\,
            in2 => \N__20450\,
            in3 => \N__20252\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIM1PUZ0Z8\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSC_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22496\,
            in2 => \N__22562\,
            in3 => \N__20249\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI34KSCZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIU5ODU_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20620\,
            in1 => \N__20465\,
            in2 => \N__22544\,
            in3 => \N__20456\,
            lcout => charx_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22514\,
            in2 => \_gnd_net_\,
            in3 => \N__20453\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22607\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22664\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RF_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20602\,
            in2 => \N__20630\,
            in3 => \N__20432\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNIRT1RFZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNO_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20621\,
            in2 => \N__20429\,
            in3 => \N__20411\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIT6SNOZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI1QD7R1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20380\,
            in1 => \N__20603\,
            in2 => \N__20408\,
            in3 => \N__20393\,
            lcout => charx_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHU_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20390\,
            in2 => \_gnd_net_\,
            in3 => \N__20384\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMELHUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_2096_i_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22461\,
            lcout => \N_2096_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23089\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIH08LF_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20619\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22618\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20594\,
            in2 => \N__20525\,
            in3 => \N__20579\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20572\,
            in2 => \N__20549\,
            in3 => \N__20528\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25870\,
            in1 => \N__20524\,
            in2 => \N__20507\,
            in3 => \N__20489\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_s_5_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20486\,
            in2 => \_gnd_net_\,
            in3 => \N__20477\,
            lcout => column_1_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_i_sbtinv_3_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25869\,
            lcout => column_1_i_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010101"
        )
    port map (
            in0 => \N__21095\,
            in1 => \N__21083\,
            in2 => \N__21278\,
            in3 => \N__21077\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_5_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000000000"
        )
    port map (
            in0 => \N__21023\,
            in1 => \N__20691\,
            in2 => \N__20884\,
            in3 => \N__24725\,
            lcout => \N_3078_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_i_sbtinv_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25285\,
            lcout => column_1_i_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_12_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001111"
        )
    port map (
            in0 => \N__23877\,
            in1 => \N__21482\,
            in2 => \N__24853\,
            in3 => \N__21494\,
            lcout => OPEN,
            ltout => \N_1297_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_1_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__24117\,
            in1 => \_gnd_net_\,
            in2 => \N__20999\,
            in3 => \N__21458\,
            lcout => \N_4564_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_14_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__20900\,
            in1 => \N__20692\,
            in2 => \N__20885\,
            in3 => \N__23335\,
            lcout => font_un67_pixel_ac0_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_4_0_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__20984\,
            in1 => \N__20939\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un113_pixel_4_0_15__g0_4_0Z0Z_0\,
            ltout => \un113_pixel_4_0_15__g0_4_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_13_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101101"
        )
    port map (
            in0 => \N__20865\,
            in1 => \N__20693\,
            in2 => \N__20633\,
            in3 => \N__23336\,
            lcout => font_un64_pixel_ac0_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJIDRG11_0_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25035\,
            in1 => \N__24229\,
            in2 => \N__24804\,
            in3 => \N__25759\,
            lcout => \beamY_RNIJIDRG11_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_4_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21296\,
            in2 => \N__21104\,
            in3 => \N__21602\,
            lcout => \N_1342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_5_4_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21269\,
            in1 => \N__21260\,
            in2 => \N__21245\,
            in3 => \N__21236\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__g0_5Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_11_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__21221\,
            in1 => \N__21185\,
            in2 => \N__21209\,
            in3 => \N__21173\,
            lcout => \N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g2_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__25036\,
            in1 => \N__24752\,
            in2 => \_gnd_net_\,
            in3 => \N__25225\,
            lcout => OPEN,
            ltout => \un113_pixel_4_0_15__g2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_20_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__21410\,
            in1 => \N__23343\,
            in2 => \N__21200\,
            in3 => \N__21197\,
            lcout => un115_pixel_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_0_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23344\,
            in1 => \N__21692\,
            in2 => \_gnd_net_\,
            in3 => \N__21179\,
            lcout => \N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_10_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__21167\,
            in1 => \N__21134\,
            in2 => \N__21122\,
            in3 => \N__24251\,
            lcout => \N_2075\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_2_s_6_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__25398\,
            in1 => \N__24748\,
            in2 => \_gnd_net_\,
            in3 => \N__21316\,
            lcout => OPEN,
            ltout => \un115_pixel_2_s_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_2_d_0_6_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110010"
        )
    port map (
            in0 => \N__23878\,
            in1 => \N__23994\,
            in2 => \N__21449\,
            in3 => \N__24540\,
            lcout => OPEN,
            ltout => \un115_pixel_2_d_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_3_bm_6_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21365\,
            in2 => \N__21446\,
            in3 => \N__25042\,
            lcout => un115_pixel_3_bm_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_RNIF16BSN1_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25742\,
            in1 => \N__21436\,
            in2 => \N__23464\,
            in3 => \N__21421\,
            lcout => \ScreenBuffer_1_0_e_0_RNIF16BSN1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_23_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__21302\,
            in1 => \N__24146\,
            in2 => \N__24827\,
            in3 => \N__23844\,
            lcout => \N_1_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_RNIHFGISN1_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__25741\,
            in1 => \N__21403\,
            in2 => \N__23465\,
            in3 => \N__21385\,
            lcout => \ScreenBuffer_1_1_e_0_RNIHFGISN1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__m8_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111101111"
        )
    port map (
            in0 => \N__24474\,
            in1 => \N__23790\,
            in2 => \N__24833\,
            in3 => \N__23956\,
            lcout => m8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_RNISDB6RM_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25518\,
            in1 => \N__21355\,
            in2 => \_gnd_net_\,
            in3 => \N__21340\,
            lcout => \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1\,
            ltout => \ScreenBuffer_1_0_e_0_RNISDB6RMZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__un115_pixel_5_s_7_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23302\,
            in2 => \N__21305\,
            in3 => \N__25415\,
            lcout => un115_pixel_5_s_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__g1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23957\,
            in1 => \N__24996\,
            in2 => \_gnd_net_\,
            in3 => \N__24475\,
            lcout => \un113_pixel_3_0_11__gZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVDIFFI1_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111000111"
        )
    port map (
            in0 => \N__24473\,
            in1 => \N__23789\,
            in2 => \N__24832\,
            in3 => \N__23955\,
            lcout => \beamY_RNIVDIFFI1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIB3R6U63_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001010000"
        )
    port map (
            in0 => \N__23954\,
            in1 => \N__24995\,
            in2 => \N__23845\,
            in3 => \N__24471\,
            lcout => \ScreenBuffer_0_7_RNIB3R6U63Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__un115_pixel_5_am_7_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111110010"
        )
    port map (
            in0 => \N__24472\,
            in1 => \N__23788\,
            in2 => \N__23345\,
            in3 => \N__23429\,
            lcout => OPEN,
            ltout => \un115_pixel_5_am_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__un115_pixel_5_ns_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21554\,
            in2 => \N__21548\,
            in3 => \N__21545\,
            lcout => \N_1288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g1_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100100000100"
        )
    port map (
            in0 => \N__25057\,
            in1 => \N__21533\,
            in2 => \N__23033\,
            in3 => \N__24510\,
            lcout => \un113_pixel_4_0_15__g1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__m9_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001100000"
        )
    port map (
            in0 => \N__24511\,
            in1 => \N__25056\,
            in2 => \N__23866\,
            in3 => \N__23971\,
            lcout => m9,
            ltout => \m9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICJUESD2_0_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__24826\,
            in1 => \_gnd_net_\,
            in2 => \N__21470\,
            in3 => \N__21467\,
            lcout => \beamY_RNICJUESD2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m6_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000100000"
        )
    port map (
            in0 => \N__24512\,
            in1 => \N__25058\,
            in2 => \N__23865\,
            in3 => \N__23970\,
            lcout => m6,
            ltout => \m6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICJUESD2_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__24825\,
            in1 => \_gnd_net_\,
            in2 => \N__21461\,
            in3 => \N__21719\,
            lcout => \beamY_RNICJUESD2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24828\,
            in1 => \N__21644\,
            in2 => \_gnd_net_\,
            in3 => \N__21638\,
            lcout => OPEN,
            ltout => \N_4562_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21632\,
            in2 => \N__21605\,
            in3 => \N__21575\,
            lcout => \N_1340_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1H36941_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21560\,
            in1 => \_gnd_net_\,
            in2 => \N__24162\,
            in3 => \N__21593\,
            lcout => \beamY_RNI1H36941Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_5_ns_x0_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__24506\,
            in1 => \N__23434\,
            in2 => \N__24855\,
            in3 => \N__25030\,
            lcout => un115_pixel_5_ns_x0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_5_ns_x1_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__23435\,
            in1 => \N__25013\,
            in2 => \N__24856\,
            in3 => \N__24507\,
            lcout => un115_pixel_5_ns_x1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__font_un125_pixel_1_bm_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23353\,
            in1 => \N__21656\,
            in2 => \_gnd_net_\,
            in3 => \N__21671\,
            lcout => font_un125_pixel_1_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_2_0_3__m7_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__23968\,
            in1 => \N__25014\,
            in2 => \_gnd_net_\,
            in3 => \N__24508\,
            lcout => \un113_pixel_2_0_3__N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_6_1_5__m10_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__24509\,
            in1 => \N__23969\,
            in2 => \N__23885\,
            in3 => \N__25031\,
            lcout => OPEN,
            ltout => \un113_pixel_6_1_5__N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICJUESD2_2_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001001110"
        )
    port map (
            in0 => \N__24816\,
            in1 => \N__23864\,
            in2 => \N__21569\,
            in3 => \N__21566\,
            lcout => \beamY_RNICJUESD2_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__m12_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__25012\,
            in1 => \N__23859\,
            in2 => \_gnd_net_\,
            in3 => \N__23967\,
            lcout => m12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__m17_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010010000"
        )
    port map (
            in0 => \N__23966\,
            in1 => \N__25011\,
            in2 => \N__23884\,
            in3 => \N__24505\,
            lcout => m17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_5_ns_ns_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21713\,
            in1 => \N__21707\,
            in2 => \_gnd_net_\,
            in3 => \N__21701\,
            lcout => OPEN,
            ltout => \N_1325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_7_bm_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24161\,
            in2 => \N__21695\,
            in3 => \N__21932\,
            lcout => un115_pixel_7_bm_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_4_3_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001010101"
        )
    port map (
            in0 => \N__24821\,
            in1 => \N__25074\,
            in2 => \_gnd_net_\,
            in3 => \N__25212\,
            lcout => OPEN,
            ltout => \N_1315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_6_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24160\,
            in2 => \N__21680\,
            in3 => \N__21677\,
            lcout => \N_1329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_1_3_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000010110000"
        )
    port map (
            in0 => \N__25070\,
            in1 => \N__25151\,
            in2 => \N__24857\,
            in3 => \N__24535\,
            lcout => OPEN,
            ltout => \N_1294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_3_ns_3_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24159\,
            in2 => \N__21665\,
            in3 => \N__21662\,
            lcout => \N_1308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_5_d_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000010"
        )
    port map (
            in0 => \N__23860\,
            in1 => \N__24002\,
            in2 => \N__24858\,
            in3 => \N__24536\,
            lcout => un115_pixel_5_d_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMR86ES2_0_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111000100"
        )
    port map (
            in0 => \N__25213\,
            in1 => \N__24817\,
            in2 => \N__25082\,
            in3 => \N__21943\,
            lcout => \beamY_RNIMR86ES2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22330\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9254_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21731\,
            in2 => \_gnd_net_\,
            in3 => \N__21917\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z9254\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIA464_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21725\,
            in2 => \N__21904\,
            in3 => \N__21764\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAZ0Z464\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22088\,
            in2 => \_gnd_net_\,
            in3 => \N__21752\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21749\,
            lcout => \chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_3_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22086\,
            lcout => chessboardpixel_un151_pixel_if_generate_plus_mult1_un47_sum_s_5_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_2_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__22193\,
            in1 => \N__22163\,
            in2 => \_gnd_net_\,
            in3 => \N__22071\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22736\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22202\,
            in2 => \N__22092\,
            in3 => \N__22376\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22100\,
            in2 => \N__21953\,
            in3 => \N__22361\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22358\,
            in2 => \N__22093\,
            in3 => \N__22334\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__22084\,
            in2 => \N__22331\,
            in3 => \N__22274\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_3_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22258\,
            lcout => un5_visiblex_i_0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__22192\,
            in1 => \N__22158\,
            in2 => \_gnd_net_\,
            in3 => \N__22077\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_charx_if_generate_plus_mult1_un26_sum_axb_3_i_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22085\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un26_sum_axb_3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22620\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22525\,
            in2 => \N__22472\,
            in3 => \N__22547\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22813\,
            in2 => \N__22397\,
            in3 => \N__22529\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI0CRJF_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22491\,
            in1 => \N__22526\,
            in2 => \N__22850\,
            in3 => \N__22502\,
            lcout => charx_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLER8_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22838\,
            in2 => \_gnd_net_\,
            in3 => \N__22499\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIHLERZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22463\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22460\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22406\,
            in2 => \N__22682\,
            in3 => \N__22388\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22778\,
            in2 => \N__22862\,
            in3 => \N__22841\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNIU99G8_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22812\,
            in1 => \N__22751\,
            in2 => \N__22793\,
            in3 => \N__22832\,
            lcout => charx_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22829\,
            in2 => \_gnd_net_\,
            in3 => \N__22820\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINP73_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__22792\,
            in1 => \N__22777\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIINPZ0Z73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22744\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23146\,
            in2 => \_gnd_net_\,
            in3 => \N__25321\,
            lcout => if_generate_plus_mult1_un75_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22673\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22672\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22634\,
            in2 => \N__23042\,
            in3 => \N__22625\,
            lcout => if_generate_plus_mult1_un75_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25400\,
            in2 => \N__23174\,
            in3 => \N__23159\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25688\,
            in1 => \N__23156\,
            in2 => \N__23150\,
            in3 => \N__23126\,
            lcout => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23123\,
            in2 => \_gnd_net_\,
            in3 => \N__23111\,
            lcout => un6_rowlto1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un6_rowlto3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__25401\,
            in1 => \N__25983\,
            in2 => \N__25512\,
            in3 => \N__25709\,
            lcout => un6_rowlt7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_i_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23093\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPPD7L31_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24834\,
            in1 => \N__23032\,
            in2 => \_gnd_net_\,
            in3 => \N__22919\,
            lcout => OPEN,
            ltout => \d_N_3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2RNL4M2_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__24001\,
            in1 => \N__23887\,
            in2 => \N__22907\,
            in3 => \N__24545\,
            lcout => \beamY_RNI2RNL4M2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__currentchar_1_4_1_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100101"
        )
    port map (
            in0 => \N__25708\,
            in1 => \N__22904\,
            in2 => \N__25517\,
            in3 => \N__22889\,
            lcout => \un113_pixel_3_0_11__currentchar_1_4_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_10_RNIGDGIE9_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__23612\,
            in1 => \N__23529\,
            in2 => \_gnd_net_\,
            in3 => \N__23717\,
            lcout => \ScreenBuffer_0_10_RNIGDGIE9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_11_RNI9RVK2F_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101111"
        )
    port map (
            in0 => \N__23530\,
            in1 => \N__23613\,
            in2 => \N__25987\,
            in3 => \N__23693\,
            lcout => OPEN,
            ltout => \currentchar_1_5_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_3_e_0_RNIR8DINK_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__25968\,
            in1 => \N__23672\,
            in2 => \N__23660\,
            in3 => \N__23657\,
            lcout => \ScreenBuffer_1_3_e_0_RNIR8DINKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_3_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25078\,
            in1 => \N__23633\,
            in2 => \_gnd_net_\,
            in3 => \N__23621\,
            lcout => \N_1303_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \currentchar_1_5_0_a2_0_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23614\,
            in2 => \N__23534\,
            in3 => \N__25969\,
            lcout => \N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_i_m2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__25150\,
            in1 => \N__25080\,
            in2 => \N__23447\,
            in3 => \N__24544\,
            lcout => OPEN,
            ltout => \N_4581_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110011"
        )
    port map (
            in0 => \N__25081\,
            in1 => \N__24835\,
            in2 => \N__23375\,
            in3 => \N__25226\,
            lcout => \N_1296_0\,
            ltout => \N_1296_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_16_x1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__24136\,
            in1 => \N__23359\,
            in2 => \N__23372\,
            in3 => \N__24010\,
            lcout => g0_16_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_16_x0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__24011\,
            in1 => \N__23369\,
            in2 => \N__23363\,
            in3 => \N__24137\,
            lcout => OPEN,
            ltout => \g0_16_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_16_ns_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24266\,
            in2 => \N__24260\,
            in3 => \N__24257\,
            lcout => \N_4560_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_2_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24135\,
            in1 => \N__24368\,
            in2 => \_gnd_net_\,
            in3 => \N__25157\,
            lcout => \N_1309_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJIDRG11_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__25075\,
            in1 => \N__24230\,
            in2 => \N__24854\,
            in3 => \N__25760\,
            lcout => OPEN,
            ltout => \beamY_RNIJIDRG11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRG0LHO1_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24212\,
            in2 => \N__24200\,
            in3 => \N__24197\,
            lcout => \beamY_RNIRG0LHO1Z0Z_0\,
            ltout => \beamY_RNIRG0LHO1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_2_x0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__24808\,
            in1 => \N__24131\,
            in2 => \N__24185\,
            in3 => \N__24181\,
            lcout => g0_2_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_2_x1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__24182\,
            in1 => \N__24809\,
            in2 => \N__24158\,
            in3 => \N__24035\,
            lcout => OPEN,
            ltout => \g0_2_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_7_1_7__g0_2_ns_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24029\,
            in2 => \N__24020\,
            in3 => \N__24017\,
            lcout => \N_1331_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_3_0_11__m15_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001010000"
        )
    port map (
            in0 => \N__24000\,
            in1 => \N__25076\,
            in2 => \N__23891\,
            in3 => \N__24543\,
            lcout => OPEN,
            ltout => \un113_pixel_3_0_11__N_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__g0_3_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__25077\,
            in1 => \N__24836\,
            in2 => \N__25229\,
            in3 => \N__25224\,
            lcout => \N_4573_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un113_pixel_4_0_15__un115_pixel_3_am_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011010000"
        )
    port map (
            in0 => \N__25149\,
            in1 => \N__25079\,
            in2 => \N__24863\,
            in3 => \N__24541\,
            lcout => un115_pixel_3_am_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24362\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24305\,
            in2 => \N__24314\,
            in3 => \N__25686\,
            lcout => \G_673\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25689\,
            in2 => \N__24299\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24281\,
            in2 => \N__24290\,
            in3 => \N__25687\,
            lcout => \G_674\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_s_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24275\,
            in2 => \_gnd_net_\,
            in3 => \N__24269\,
            lcout => un6_rowlto0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_10_RNIB0Q4B12_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111101010"
        )
    port map (
            in0 => \N__25690\,
            in1 => \N__25966\,
            in2 => \N__25811\,
            in3 => \N__25819\,
            lcout => \ScreenBuffer_0_10_RNIB0Q4B12Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_10_RNIB0Q4B12_0_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__25967\,
            in1 => \N__25691\,
            in2 => \N__25823\,
            in3 => \N__25807\,
            lcout => OPEN,
            ltout => \ScreenBuffer_0_10_RNIB0Q4B12_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_RNI1J74DN_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25790\,
            in2 => \N__25781\,
            in3 => \N__25778\,
            lcout => \ScreenBuffer_1_0_e_0_RNI1J74DNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_6_RNITJ4B17_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__25397\,
            in1 => \N__25772\,
            in2 => \N__25513\,
            in3 => \N__25235\,
            lcout => \ScreenBuffer_0_6_RNITJ4B17Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__25692\,
            in1 => \N__25478\,
            in2 => \N__25625\,
            in3 => \N__25633\,
            lcout => \ScreenBuffer_1_1_e_0_RNIHD6DAP3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_1_e_0_RNIHD6DAP3_0_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__25477\,
            in1 => \N__25693\,
            in2 => \N__25637\,
            in3 => \N__25621\,
            lcout => OPEN,
            ltout => \ScreenBuffer_1_1_e_0_RNIHD6DAP3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_1_0_e_0_RNI3EKU1A_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25607\,
            in2 => \N__25601\,
            in3 => \N__25598\,
            lcout => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0\,
            ltout => \ScreenBuffer_1_0_e_0_RNI3EKU1AZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ScreenBuffer_0_7_RNIS4U201_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__25479\,
            in1 => \N__25402\,
            in2 => \N__25256\,
            in3 => \N__25253\,
            lcout => un115_pixel_5_am_sx_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
