// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 16:21:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSync,
    Pixel,
    HSync,
    Clock12MHz);

    output VSync;
    output Pixel;
    output HSync;
    input Clock12MHz;

    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4753;
    wire N__4752;
    wire N__4751;
    wire N__4744;
    wire N__4743;
    wire N__4742;
    wire N__4735;
    wire N__4734;
    wire N__4733;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4709;
    wire N__4708;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4676;
    wire N__4671;
    wire N__4666;
    wire N__4663;
    wire N__4662;
    wire N__4659;
    wire N__4654;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4637;
    wire N__4632;
    wire N__4627;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4584;
    wire N__4581;
    wire N__4580;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4568;
    wire N__4567;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4540;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4478;
    wire N__4477;
    wire N__4476;
    wire N__4475;
    wire N__4474;
    wire N__4473;
    wire N__4472;
    wire N__4471;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4435;
    wire N__4434;
    wire N__4433;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4353;
    wire N__4350;
    wire N__4349;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4277;
    wire N__4276;
    wire N__4275;
    wire N__4274;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4257;
    wire N__4252;
    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4230;
    wire N__4225;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4202;
    wire N__4199;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4179;
    wire N__4176;
    wire N__4175;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4159;
    wire N__4158;
    wire N__4157;
    wire N__4156;
    wire N__4151;
    wire N__4144;
    wire N__4135;
    wire N__4134;
    wire N__4133;
    wire N__4130;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4089;
    wire N__4088;
    wire N__4087;
    wire N__4086;
    wire N__4085;
    wire N__4084;
    wire N__4081;
    wire N__4072;
    wire N__4069;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4005;
    wire N__4002;
    wire N__4001;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3962;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3864;
    wire N__3863;
    wire N__3860;
    wire N__3859;
    wire N__3856;
    wire N__3851;
    wire N__3846;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3834;
    wire N__3833;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3788;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3764;
    wire N__3763;
    wire N__3762;
    wire N__3759;
    wire N__3752;
    wire N__3747;
    wire N__3744;
    wire N__3743;
    wire N__3742;
    wire N__3739;
    wire N__3734;
    wire N__3729;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3707;
    wire N__3706;
    wire N__3705;
    wire N__3704;
    wire N__3703;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3664;
    wire N__3657;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3645;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3581;
    wire N__3580;
    wire N__3579;
    wire N__3576;
    wire N__3569;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3531;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3519;
    wire N__3516;
    wire N__3515;
    wire N__3514;
    wire N__3513;
    wire N__3512;
    wire N__3511;
    wire N__3510;
    wire N__3509;
    wire N__3508;
    wire N__3507;
    wire N__3506;
    wire N__3505;
    wire N__3504;
    wire N__3503;
    wire N__3502;
    wire N__3495;
    wire N__3486;
    wire N__3477;
    wire N__3468;
    wire N__3459;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3447;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3435;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3423;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3411;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3399;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3360;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3348;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3323;
    wire N__3322;
    wire N__3319;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3304;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3284;
    wire N__3281;
    wire N__3280;
    wire N__3277;
    wire N__3276;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3226;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3213;
    wire N__3208;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3194;
    wire N__3193;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3165;
    wire N__3162;
    wire N__3161;
    wire N__3160;
    wire N__3159;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3131;
    wire N__3130;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3105;
    wire N__3102;
    wire N__3101;
    wire N__3100;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3088;
    wire N__3081;
    wire N__3078;
    wire N__3077;
    wire N__3076;
    wire N__3073;
    wire N__3068;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3056;
    wire N__3055;
    wire N__3052;
    wire N__3051;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3036;
    wire N__3031;
    wire N__3024;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3012;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3000;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2966;
    wire N__2965;
    wire N__2960;
    wire N__2957;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2939;
    wire N__2936;
    wire N__2935;
    wire N__2934;
    wire N__2927;
    wire N__2924;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2882;
    wire N__2881;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2864;
    wire N__2861;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2828;
    wire N__2825;
    wire N__2824;
    wire N__2823;
    wire N__2816;
    wire N__2813;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2756;
    wire N__2753;
    wire N__2752;
    wire N__2751;
    wire N__2744;
    wire N__2741;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2666;
    wire N__2663;
    wire N__2662;
    wire N__2661;
    wire N__2654;
    wire N__2651;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2613;
    wire N__2612;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2593;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2581;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2565;
    wire N__2562;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2543;
    wire N__2542;
    wire N__2539;
    wire N__2538;
    wire N__2535;
    wire N__2534;
    wire N__2531;
    wire N__2522;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2508;
    wire N__2505;
    wire N__2502;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2421;
    wire N__2418;
    wire N__2415;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2397;
    wire N__2394;
    wire N__2391;
    wire N__2388;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2373;
    wire N__2370;
    wire N__2367;
    wire N__2364;
    wire N__2361;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2349;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2331;
    wire N__2328;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2313;
    wire N__2310;
    wire N__2309;
    wire N__2308;
    wire N__2305;
    wire N__2304;
    wire N__2301;
    wire N__2294;
    wire N__2291;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2265;
    wire N__2262;
    wire N__2259;
    wire N__2256;
    wire N__2253;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_1_0_;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un61_sum_i_0;
    wire bfn_1_2_0_;
    wire un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_;
    wire un2_y_if_generate_plus_mult1_un61_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_i_0;
    wire bfn_1_3_0_;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_;
    wire bfn_1_4_0_;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un40_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_i_0;
    wire un13_x_i_i_a2_1;
    wire N_130_cascade_;
    wire y_RNIA5P7Z0Z_9;
    wire un13_x_i_i_a2_0_3_cascade_;
    wire bfn_1_6_0_;
    wire Counter_cry_0;
    wire Counter_cry_1;
    wire Counter_cry_2;
    wire Counter_cry_3;
    wire Counter_cry_4;
    wire Counter_cry_5;
    wire Counter_cry_6;
    wire Counter_cry_7;
    wire bfn_1_7_0_;
    wire Counter_cry_8;
    wire Counter_cry_9;
    wire Counter_cry_10;
    wire Counter_cry_11;
    wire Counter_cry_12;
    wire ClockVGAZ0;
    wire Clock12MHz_c_g;
    wire G_167;
    wire bfn_2_1_0_;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un75_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un68_sum_i_0;
    wire bfn_2_2_0_;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un61_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_;
    wire un2_y_if_generate_plus_mult1_un54_sum_i_7;
    wire bfn_2_3_0_;
    wire un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81;
    wire un2_y_if_generate_plus_mult1_un40_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un47_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_;
    wire un2_y_if_generate_plus_mult1_un47_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un47_sum_i_0;
    wire bfn_2_4_0_;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_;
    wire un2_y_if_generate_plus_mult1_un33_sum_i_7;
    wire N_140;
    wire un2_y_if_generate_plus_mult1_un40_sum_i_0;
    wire yZ0Z_0;
    wire bfn_2_5_0_;
    wire un3_y_cry_1_THRU_CO;
    wire un3_y_cry_1;
    wire yZ0Z_3;
    wire un3_y_cry_2_THRU_CO;
    wire un3_y_cry_2;
    wire yZ0Z_4;
    wire un3_y_cry_3;
    wire yZ0Z_5;
    wire un3_y_cry_4;
    wire yZ0Z_6;
    wire un3_y_cry_5;
    wire yZ0Z_7;
    wire un3_y_cry_6;
    wire yZ0Z_8;
    wire un3_y_cry_7;
    wire un3_y_cry_8;
    wire N_130;
    wire bfn_2_6_0_;
    wire yZ0Z_9;
    wire CounterZ0Z_7;
    wire CounterZ0Z_6;
    wire CounterZ0Z_8;
    wire CounterZ0Z_13;
    wire CounterZ0Z_12;
    wire un2_counterlt11_cascade_;
    wire un2_counter_0;
    wire CounterZ0Z_4;
    wire CounterZ0Z_0;
    wire CounterZ0Z_3;
    wire CounterZ0Z_2;
    wire CounterZ0Z_1;
    wire CounterZ0Z_5;
    wire un2_counterlto4_2;
    wire un2_counterlt7;
    wire CounterZ0Z_11;
    wire CounterZ0Z_9;
    wire CounterZ0Z_10;
    wire un2_counterlto11_1;
    wire N_83_cascade_;
    wire N_85;
    wire un13lto4_i_1_cascade_;
    wire CONSTANT_ONE_NET_cascade_;
    wire yZ0Z_2;
    wire un2_y_if_generate_plus_mult1_un75_sum_i_0;
    wire bfn_5_1_0_;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0;
    wire un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO;
    wire un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1;
    wire un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO;
    wire un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3;
    wire Pixel_RNOZ0Z_4;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1;
    wire N_49;
    wire un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4;
    wire bfn_5_2_0_;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un68_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_;
    wire un2_x_if_generate_plus_mult1_un68_sum_i;
    wire xZ0Z_0;
    wire xZ0Z_1;
    wire bfn_5_4_0_;
    wire xZ0Z_2;
    wire un16_x_cry_1;
    wire N_89;
    wire un16_x_cry_2;
    wire un16_x_cry_3;
    wire un16_x_cry_4;
    wire un16_x_cry_5;
    wire un16_x_cry_6;
    wire un16_x_cry_7;
    wire un16_x_cry_8;
    wire bfn_5_5_0_;
    wire bfn_6_1_0_;
    wire un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4;
    wire Pixel_RNOZ0Z_6;
    wire un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0;
    wire un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO;
    wire N_57;
    wire N_59;
    wire N_55;
    wire N_47;
    wire Pixel_c;
    wire bfn_6_2_0_;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un75_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5;
    wire un2_x_if_generate_plus_mult1_un75_sum_i_0;
    wire bfn_6_3_0_;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un68_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_;
    wire un2_x_if_generate_plus_mult1_un61_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un61_sum_i;
    wire un2_x_if_generate_plus_mult1_un54_sum_i;
    wire Pixel_0_sqmuxa_i_1;
    wire Pixel_0_sqmuxa_i_0;
    wire HSync_c;
    wire N_90;
    wire xZ0Z_5;
    wire xZ0Z_6;
    wire xZ0Z_4;
    wire un11_x_0_a2_2_2;
    wire un11_x_0_a2_1_cascade_;
    wire x_RNID8R22Z0Z_9;
    wire xZ0Z_9;
    wire un1_xlto9_i_0;
    wire bfn_6_5_0_;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_;
    wire xZ0Z_7;
    wire bfn_7_3_0_;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un61_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_;
    wire un2_x_if_generate_plus_mult1_un54_sum_i_8;
    wire bfn_7_4_0_;
    wire un2_x_if_generate_plus_mult1_un40_sum_i;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8;
    wire CONSTANT_ONE_NET;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un54_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_;
    wire un2_x_if_generate_plus_mult1_un47_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0;
    wire xZ0Z_8;
    wire un2_x_if_generate_plus_mult1_un47_sum_i;
    wire y_RNIMA162Z0Z_9;
    wire VSync_c;
    wire ClockVGA_g;
    wire _gnd_net_;

    PRE_IO_GBUF Clock12MHz_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__4762),
            .GLOBALBUFFEROUTPUT(Clock12MHz_c_g));
    defparam Clock12MHz_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_gb_io_iopad (
            .OE(N__4764),
            .DIN(N__4763),
            .DOUT(N__4762),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_gb_io_preio (
            .PADOEN(N__4764),
            .PADOUT(N__4763),
            .PADIN(N__4762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__4753),
            .DIN(N__4752),
            .DOUT(N__4751),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__4753),
            .PADOUT(N__4752),
            .PADIN(N__4751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__4744),
            .DIN(N__4743),
            .DOUT(N__4742),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__4744),
            .PADOUT(N__4743),
            .PADIN(N__4742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4302),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__4735),
            .DIN(N__4734),
            .DOUT(N__4733),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__4735),
            .PADOUT(N__4734),
            .PADIN(N__4733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1021 (
            .O(N__4716),
            .I(N__4713));
    LocalMux I__1020 (
            .O(N__4713),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8));
    CascadeMux I__1019 (
            .O(N__4710),
            .I(N__4703));
    CascadeMux I__1018 (
            .O(N__4709),
            .I(N__4700));
    CascadeMux I__1017 (
            .O(N__4708),
            .I(N__4696));
    CascadeMux I__1016 (
            .O(N__4707),
            .I(N__4693));
    CascadeMux I__1015 (
            .O(N__4706),
            .I(N__4690));
    InMux I__1014 (
            .O(N__4703),
            .I(N__4684));
    InMux I__1013 (
            .O(N__4700),
            .I(N__4681));
    InMux I__1012 (
            .O(N__4699),
            .I(N__4676));
    InMux I__1011 (
            .O(N__4696),
            .I(N__4676));
    InMux I__1010 (
            .O(N__4693),
            .I(N__4671));
    InMux I__1009 (
            .O(N__4690),
            .I(N__4671));
    InMux I__1008 (
            .O(N__4689),
            .I(N__4666));
    InMux I__1007 (
            .O(N__4688),
            .I(N__4666));
    InMux I__1006 (
            .O(N__4687),
            .I(N__4663));
    LocalMux I__1005 (
            .O(N__4684),
            .I(N__4659));
    LocalMux I__1004 (
            .O(N__4681),
            .I(N__4654));
    LocalMux I__1003 (
            .O(N__4676),
            .I(N__4654));
    LocalMux I__1002 (
            .O(N__4671),
            .I(N__4649));
    LocalMux I__1001 (
            .O(N__4666),
            .I(N__4649));
    LocalMux I__1000 (
            .O(N__4663),
            .I(N__4646));
    CascadeMux I__999 (
            .O(N__4662),
            .I(N__4643));
    Span4Mux_h I__998 (
            .O(N__4659),
            .I(N__4637));
    Span4Mux_s3_h I__997 (
            .O(N__4654),
            .I(N__4637));
    Span4Mux_v I__996 (
            .O(N__4649),
            .I(N__4632));
    Span4Mux_v I__995 (
            .O(N__4646),
            .I(N__4632));
    InMux I__994 (
            .O(N__4643),
            .I(N__4627));
    InMux I__993 (
            .O(N__4642),
            .I(N__4627));
    Odrv4 I__992 (
            .O(N__4637),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__991 (
            .O(N__4632),
            .I(CONSTANT_ONE_NET));
    LocalMux I__990 (
            .O(N__4627),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__989 (
            .O(N__4620),
            .I(N__4617));
    InMux I__988 (
            .O(N__4617),
            .I(N__4614));
    LocalMux I__987 (
            .O(N__4614),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0));
    InMux I__986 (
            .O(N__4611),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__985 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__984 (
            .O(N__4605),
            .I(un2_x_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__983 (
            .O(N__4602),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__982 (
            .O(N__4599),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__981 (
            .O(N__4596),
            .I(N__4592));
    InMux I__980 (
            .O(N__4595),
            .I(N__4589));
    LocalMux I__979 (
            .O(N__4592),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0));
    LocalMux I__978 (
            .O(N__4589),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0));
    CascadeMux I__977 (
            .O(N__4584),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_));
    InMux I__976 (
            .O(N__4581),
            .I(N__4575));
    InMux I__975 (
            .O(N__4580),
            .I(N__4575));
    LocalMux I__974 (
            .O(N__4575),
            .I(un2_x_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__973 (
            .O(N__4572),
            .I(N__4569));
    InMux I__972 (
            .O(N__4569),
            .I(N__4560));
    InMux I__971 (
            .O(N__4568),
            .I(N__4560));
    InMux I__970 (
            .O(N__4567),
            .I(N__4560));
    LocalMux I__969 (
            .O(N__4560),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__968 (
            .O(N__4557),
            .I(N__4554));
    LocalMux I__967 (
            .O(N__4554),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0));
    InMux I__966 (
            .O(N__4551),
            .I(N__4540));
    InMux I__965 (
            .O(N__4550),
            .I(N__4540));
    InMux I__964 (
            .O(N__4549),
            .I(N__4535));
    InMux I__963 (
            .O(N__4548),
            .I(N__4535));
    InMux I__962 (
            .O(N__4547),
            .I(N__4532));
    InMux I__961 (
            .O(N__4546),
            .I(N__4529));
    InMux I__960 (
            .O(N__4545),
            .I(N__4526));
    LocalMux I__959 (
            .O(N__4540),
            .I(N__4521));
    LocalMux I__958 (
            .O(N__4535),
            .I(N__4521));
    LocalMux I__957 (
            .O(N__4532),
            .I(xZ0Z_8));
    LocalMux I__956 (
            .O(N__4529),
            .I(xZ0Z_8));
    LocalMux I__955 (
            .O(N__4526),
            .I(xZ0Z_8));
    Odrv4 I__954 (
            .O(N__4521),
            .I(xZ0Z_8));
    CascadeMux I__953 (
            .O(N__4512),
            .I(N__4509));
    InMux I__952 (
            .O(N__4509),
            .I(N__4506));
    LocalMux I__951 (
            .O(N__4506),
            .I(un2_x_if_generate_plus_mult1_un47_sum_i));
    InMux I__950 (
            .O(N__4503),
            .I(N__4499));
    InMux I__949 (
            .O(N__4502),
            .I(N__4496));
    LocalMux I__948 (
            .O(N__4499),
            .I(N__4491));
    LocalMux I__947 (
            .O(N__4496),
            .I(N__4491));
    Odrv12 I__946 (
            .O(N__4491),
            .I(y_RNIMA162Z0Z_9));
    IoInMux I__945 (
            .O(N__4488),
            .I(N__4485));
    LocalMux I__944 (
            .O(N__4485),
            .I(N__4482));
    Odrv12 I__943 (
            .O(N__4482),
            .I(VSync_c));
    ClkMux I__942 (
            .O(N__4479),
            .I(N__4452));
    ClkMux I__941 (
            .O(N__4478),
            .I(N__4452));
    ClkMux I__940 (
            .O(N__4477),
            .I(N__4452));
    ClkMux I__939 (
            .O(N__4476),
            .I(N__4452));
    ClkMux I__938 (
            .O(N__4475),
            .I(N__4452));
    ClkMux I__937 (
            .O(N__4474),
            .I(N__4452));
    ClkMux I__936 (
            .O(N__4473),
            .I(N__4452));
    ClkMux I__935 (
            .O(N__4472),
            .I(N__4452));
    ClkMux I__934 (
            .O(N__4471),
            .I(N__4452));
    GlobalMux I__933 (
            .O(N__4452),
            .I(N__4449));
    gio2CtrlBuf I__932 (
            .O(N__4449),
            .I(ClockVGA_g));
    CascadeMux I__931 (
            .O(N__4446),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_));
    InMux I__930 (
            .O(N__4443),
            .I(N__4439));
    CascadeMux I__929 (
            .O(N__4442),
            .I(N__4436));
    LocalMux I__928 (
            .O(N__4439),
            .I(N__4429));
    InMux I__927 (
            .O(N__4436),
            .I(N__4426));
    InMux I__926 (
            .O(N__4435),
            .I(N__4423));
    InMux I__925 (
            .O(N__4434),
            .I(N__4418));
    InMux I__924 (
            .O(N__4433),
            .I(N__4418));
    InMux I__923 (
            .O(N__4432),
            .I(N__4415));
    Span4Mux_h I__922 (
            .O(N__4429),
            .I(N__4412));
    LocalMux I__921 (
            .O(N__4426),
            .I(xZ0Z_7));
    LocalMux I__920 (
            .O(N__4423),
            .I(xZ0Z_7));
    LocalMux I__919 (
            .O(N__4418),
            .I(xZ0Z_7));
    LocalMux I__918 (
            .O(N__4415),
            .I(xZ0Z_7));
    Odrv4 I__917 (
            .O(N__4412),
            .I(xZ0Z_7));
    CascadeMux I__916 (
            .O(N__4401),
            .I(N__4398));
    InMux I__915 (
            .O(N__4398),
            .I(N__4395));
    LocalMux I__914 (
            .O(N__4395),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0));
    InMux I__913 (
            .O(N__4392),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__912 (
            .O(N__4389),
            .I(N__4386));
    InMux I__911 (
            .O(N__4386),
            .I(N__4383));
    LocalMux I__910 (
            .O(N__4383),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0));
    InMux I__909 (
            .O(N__4380),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__908 (
            .O(N__4377),
            .I(N__4374));
    LocalMux I__907 (
            .O(N__4374),
            .I(un2_x_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__906 (
            .O(N__4371),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__905 (
            .O(N__4368),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__904 (
            .O(N__4365),
            .I(N__4361));
    InMux I__903 (
            .O(N__4364),
            .I(N__4358));
    LocalMux I__902 (
            .O(N__4361),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1));
    LocalMux I__901 (
            .O(N__4358),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1));
    CascadeMux I__900 (
            .O(N__4353),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_));
    InMux I__899 (
            .O(N__4350),
            .I(N__4344));
    InMux I__898 (
            .O(N__4349),
            .I(N__4344));
    LocalMux I__897 (
            .O(N__4344),
            .I(un2_x_if_generate_plus_mult1_un54_sum_i_8));
    InMux I__896 (
            .O(N__4341),
            .I(N__4338));
    LocalMux I__895 (
            .O(N__4338),
            .I(un2_x_if_generate_plus_mult1_un40_sum_i));
    CascadeMux I__894 (
            .O(N__4335),
            .I(N__4332));
    InMux I__893 (
            .O(N__4332),
            .I(N__4329));
    LocalMux I__892 (
            .O(N__4329),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0));
    InMux I__891 (
            .O(N__4326),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__890 (
            .O(N__4323),
            .I(N__4320));
    InMux I__889 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__888 (
            .O(N__4317),
            .I(N__4314));
    Odrv4 I__887 (
            .O(N__4314),
            .I(Pixel_0_sqmuxa_i_1));
    InMux I__886 (
            .O(N__4311),
            .I(N__4308));
    LocalMux I__885 (
            .O(N__4308),
            .I(N__4305));
    Odrv4 I__884 (
            .O(N__4305),
            .I(Pixel_0_sqmuxa_i_0));
    IoInMux I__883 (
            .O(N__4302),
            .I(N__4299));
    LocalMux I__882 (
            .O(N__4299),
            .I(N__4296));
    IoSpan4Mux I__881 (
            .O(N__4296),
            .I(N__4293));
    Span4Mux_s2_v I__880 (
            .O(N__4293),
            .I(N__4290));
    Odrv4 I__879 (
            .O(N__4290),
            .I(HSync_c));
    CascadeMux I__878 (
            .O(N__4287),
            .I(N__4284));
    InMux I__877 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__876 (
            .O(N__4281),
            .I(N_90));
    InMux I__875 (
            .O(N__4278),
            .I(N__4270));
    InMux I__874 (
            .O(N__4277),
            .I(N__4267));
    InMux I__873 (
            .O(N__4276),
            .I(N__4264));
    InMux I__872 (
            .O(N__4275),
            .I(N__4257));
    InMux I__871 (
            .O(N__4274),
            .I(N__4257));
    InMux I__870 (
            .O(N__4273),
            .I(N__4257));
    LocalMux I__869 (
            .O(N__4270),
            .I(N__4252));
    LocalMux I__868 (
            .O(N__4267),
            .I(N__4252));
    LocalMux I__867 (
            .O(N__4264),
            .I(xZ0Z_5));
    LocalMux I__866 (
            .O(N__4257),
            .I(xZ0Z_5));
    Odrv4 I__865 (
            .O(N__4252),
            .I(xZ0Z_5));
    InMux I__864 (
            .O(N__4245),
            .I(N__4237));
    InMux I__863 (
            .O(N__4244),
            .I(N__4230));
    InMux I__862 (
            .O(N__4243),
            .I(N__4230));
    InMux I__861 (
            .O(N__4242),
            .I(N__4230));
    InMux I__860 (
            .O(N__4241),
            .I(N__4225));
    InMux I__859 (
            .O(N__4240),
            .I(N__4225));
    LocalMux I__858 (
            .O(N__4237),
            .I(xZ0Z_6));
    LocalMux I__857 (
            .O(N__4230),
            .I(xZ0Z_6));
    LocalMux I__856 (
            .O(N__4225),
            .I(xZ0Z_6));
    CascadeMux I__855 (
            .O(N__4218),
            .I(N__4210));
    InMux I__854 (
            .O(N__4217),
            .I(N__4207));
    InMux I__853 (
            .O(N__4216),
            .I(N__4202));
    InMux I__852 (
            .O(N__4215),
            .I(N__4202));
    InMux I__851 (
            .O(N__4214),
            .I(N__4199));
    InMux I__850 (
            .O(N__4213),
            .I(N__4194));
    InMux I__849 (
            .O(N__4210),
            .I(N__4194));
    LocalMux I__848 (
            .O(N__4207),
            .I(N__4191));
    LocalMux I__847 (
            .O(N__4202),
            .I(N__4188));
    LocalMux I__846 (
            .O(N__4199),
            .I(xZ0Z_4));
    LocalMux I__845 (
            .O(N__4194),
            .I(xZ0Z_4));
    Odrv4 I__844 (
            .O(N__4191),
            .I(xZ0Z_4));
    Odrv4 I__843 (
            .O(N__4188),
            .I(xZ0Z_4));
    CascadeMux I__842 (
            .O(N__4179),
            .I(N__4176));
    InMux I__841 (
            .O(N__4176),
            .I(N__4170));
    InMux I__840 (
            .O(N__4175),
            .I(N__4170));
    LocalMux I__839 (
            .O(N__4170),
            .I(un11_x_0_a2_2_2));
    CascadeMux I__838 (
            .O(N__4167),
            .I(un11_x_0_a2_1_cascade_));
    InMux I__837 (
            .O(N__4164),
            .I(N__4151));
    InMux I__836 (
            .O(N__4163),
            .I(N__4151));
    InMux I__835 (
            .O(N__4162),
            .I(N__4144));
    InMux I__834 (
            .O(N__4161),
            .I(N__4144));
    InMux I__833 (
            .O(N__4160),
            .I(N__4144));
    InMux I__832 (
            .O(N__4159),
            .I(N__4135));
    InMux I__831 (
            .O(N__4158),
            .I(N__4135));
    InMux I__830 (
            .O(N__4157),
            .I(N__4135));
    InMux I__829 (
            .O(N__4156),
            .I(N__4135));
    LocalMux I__828 (
            .O(N__4151),
            .I(N__4130));
    LocalMux I__827 (
            .O(N__4144),
            .I(N__4125));
    LocalMux I__826 (
            .O(N__4135),
            .I(N__4125));
    InMux I__825 (
            .O(N__4134),
            .I(N__4122));
    InMux I__824 (
            .O(N__4133),
            .I(N__4119));
    Span4Mux_v I__823 (
            .O(N__4130),
            .I(N__4110));
    Span4Mux_v I__822 (
            .O(N__4125),
            .I(N__4110));
    LocalMux I__821 (
            .O(N__4122),
            .I(N__4110));
    LocalMux I__820 (
            .O(N__4119),
            .I(N__4107));
    InMux I__819 (
            .O(N__4118),
            .I(N__4104));
    InMux I__818 (
            .O(N__4117),
            .I(N__4101));
    Span4Mux_h I__817 (
            .O(N__4110),
            .I(N__4098));
    Odrv4 I__816 (
            .O(N__4107),
            .I(x_RNID8R22Z0Z_9));
    LocalMux I__815 (
            .O(N__4104),
            .I(x_RNID8R22Z0Z_9));
    LocalMux I__814 (
            .O(N__4101),
            .I(x_RNID8R22Z0Z_9));
    Odrv4 I__813 (
            .O(N__4098),
            .I(x_RNID8R22Z0Z_9));
    InMux I__812 (
            .O(N__4089),
            .I(N__4081));
    InMux I__811 (
            .O(N__4088),
            .I(N__4072));
    InMux I__810 (
            .O(N__4087),
            .I(N__4072));
    InMux I__809 (
            .O(N__4086),
            .I(N__4072));
    InMux I__808 (
            .O(N__4085),
            .I(N__4072));
    InMux I__807 (
            .O(N__4084),
            .I(N__4069));
    LocalMux I__806 (
            .O(N__4081),
            .I(xZ0Z_9));
    LocalMux I__805 (
            .O(N__4072),
            .I(xZ0Z_9));
    LocalMux I__804 (
            .O(N__4069),
            .I(xZ0Z_9));
    InMux I__803 (
            .O(N__4062),
            .I(N__4059));
    LocalMux I__802 (
            .O(N__4059),
            .I(un1_xlto9_i_0));
    InMux I__801 (
            .O(N__4056),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5));
    CascadeMux I__800 (
            .O(N__4053),
            .I(N__4050));
    InMux I__799 (
            .O(N__4050),
            .I(N__4047));
    LocalMux I__798 (
            .O(N__4047),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02));
    InMux I__797 (
            .O(N__4044),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__796 (
            .O(N__4041),
            .I(N__4038));
    InMux I__795 (
            .O(N__4038),
            .I(N__4035));
    LocalMux I__794 (
            .O(N__4035),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2));
    InMux I__793 (
            .O(N__4032),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__792 (
            .O(N__4029),
            .I(N__4026));
    LocalMux I__791 (
            .O(N__4026),
            .I(un2_x_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__790 (
            .O(N__4023),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__789 (
            .O(N__4020),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__788 (
            .O(N__4017),
            .I(N__4013));
    InMux I__787 (
            .O(N__4016),
            .I(N__4010));
    LocalMux I__786 (
            .O(N__4013),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2));
    LocalMux I__785 (
            .O(N__4010),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2));
    CascadeMux I__784 (
            .O(N__4005),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_));
    InMux I__783 (
            .O(N__4002),
            .I(N__3996));
    InMux I__782 (
            .O(N__4001),
            .I(N__3996));
    LocalMux I__781 (
            .O(N__3996),
            .I(un2_x_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__780 (
            .O(N__3993),
            .I(N__3990));
    InMux I__779 (
            .O(N__3990),
            .I(N__3987));
    LocalMux I__778 (
            .O(N__3987),
            .I(un2_x_if_generate_plus_mult1_un61_sum_i));
    CascadeMux I__777 (
            .O(N__3984),
            .I(N__3981));
    InMux I__776 (
            .O(N__3981),
            .I(N__3978));
    LocalMux I__775 (
            .O(N__3978),
            .I(un2_x_if_generate_plus_mult1_un54_sum_i));
    InMux I__774 (
            .O(N__3975),
            .I(N__3972));
    LocalMux I__773 (
            .O(N__3972),
            .I(Pixel_RNOZ0Z_6));
    InMux I__772 (
            .O(N__3969),
            .I(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5));
    CascadeMux I__771 (
            .O(N__3966),
            .I(N__3963));
    InMux I__770 (
            .O(N__3963),
            .I(N__3957));
    InMux I__769 (
            .O(N__3962),
            .I(N__3957));
    LocalMux I__768 (
            .O(N__3957),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747));
    InMux I__767 (
            .O(N__3954),
            .I(N__3948));
    InMux I__766 (
            .O(N__3953),
            .I(N__3948));
    LocalMux I__765 (
            .O(N__3948),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0));
    CascadeMux I__764 (
            .O(N__3945),
            .I(N__3942));
    InMux I__763 (
            .O(N__3942),
            .I(N__3939));
    LocalMux I__762 (
            .O(N__3939),
            .I(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO));
    InMux I__761 (
            .O(N__3936),
            .I(N__3933));
    LocalMux I__760 (
            .O(N__3933),
            .I(N_57));
    CascadeMux I__759 (
            .O(N__3930),
            .I(N__3927));
    InMux I__758 (
            .O(N__3927),
            .I(N__3924));
    LocalMux I__757 (
            .O(N__3924),
            .I(N_59));
    InMux I__756 (
            .O(N__3921),
            .I(N__3918));
    LocalMux I__755 (
            .O(N__3918),
            .I(N_55));
    InMux I__754 (
            .O(N__3915),
            .I(N__3912));
    LocalMux I__753 (
            .O(N__3912),
            .I(N_47));
    IoInMux I__752 (
            .O(N__3909),
            .I(N__3906));
    LocalMux I__751 (
            .O(N__3906),
            .I(N__3903));
    Span4Mux_s0_v I__750 (
            .O(N__3903),
            .I(N__3900));
    Odrv4 I__749 (
            .O(N__3900),
            .I(Pixel_c));
    InMux I__748 (
            .O(N__3897),
            .I(N__3894));
    LocalMux I__747 (
            .O(N__3894),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3));
    InMux I__746 (
            .O(N__3891),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__745 (
            .O(N__3888),
            .I(N__3885));
    InMux I__744 (
            .O(N__3885),
            .I(N__3882));
    LocalMux I__743 (
            .O(N__3882),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465));
    InMux I__742 (
            .O(N__3879),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__741 (
            .O(N__3876),
            .I(N__3873));
    LocalMux I__740 (
            .O(N__3873),
            .I(un2_x_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__739 (
            .O(N__3870),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__738 (
            .O(N__3867),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__737 (
            .O(N__3864),
            .I(N__3860));
    InMux I__736 (
            .O(N__3863),
            .I(N__3856));
    InMux I__735 (
            .O(N__3860),
            .I(N__3851));
    InMux I__734 (
            .O(N__3859),
            .I(N__3851));
    LocalMux I__733 (
            .O(N__3856),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5));
    LocalMux I__732 (
            .O(N__3851),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5));
    InMux I__731 (
            .O(N__3846),
            .I(N__3842));
    InMux I__730 (
            .O(N__3845),
            .I(N__3839));
    LocalMux I__729 (
            .O(N__3842),
            .I(un2_x_if_generate_plus_mult1_un75_sum_i_0));
    LocalMux I__728 (
            .O(N__3839),
            .I(un2_x_if_generate_plus_mult1_un75_sum_i_0));
    InMux I__727 (
            .O(N__3834),
            .I(N__3829));
    InMux I__726 (
            .O(N__3833),
            .I(N__3826));
    InMux I__725 (
            .O(N__3832),
            .I(N__3823));
    LocalMux I__724 (
            .O(N__3829),
            .I(N__3820));
    LocalMux I__723 (
            .O(N__3826),
            .I(N_89));
    LocalMux I__722 (
            .O(N__3823),
            .I(N_89));
    Odrv4 I__721 (
            .O(N__3820),
            .I(N_89));
    InMux I__720 (
            .O(N__3813),
            .I(un16_x_cry_2));
    InMux I__719 (
            .O(N__3810),
            .I(un16_x_cry_3));
    InMux I__718 (
            .O(N__3807),
            .I(un16_x_cry_4));
    InMux I__717 (
            .O(N__3804),
            .I(un16_x_cry_5));
    InMux I__716 (
            .O(N__3801),
            .I(un16_x_cry_6));
    InMux I__715 (
            .O(N__3798),
            .I(un16_x_cry_7));
    InMux I__714 (
            .O(N__3795),
            .I(bfn_5_5_0_));
    InMux I__713 (
            .O(N__3792),
            .I(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4));
    InMux I__712 (
            .O(N__3789),
            .I(N__3783));
    InMux I__711 (
            .O(N__3788),
            .I(N__3783));
    LocalMux I__710 (
            .O(N__3783),
            .I(un2_x_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__709 (
            .O(N__3780),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__708 (
            .O(N__3777),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_));
    CascadeMux I__707 (
            .O(N__3774),
            .I(N__3771));
    InMux I__706 (
            .O(N__3771),
            .I(N__3768));
    LocalMux I__705 (
            .O(N__3768),
            .I(un2_x_if_generate_plus_mult1_un68_sum_i));
    InMux I__704 (
            .O(N__3765),
            .I(N__3759));
    InMux I__703 (
            .O(N__3764),
            .I(N__3752));
    InMux I__702 (
            .O(N__3763),
            .I(N__3752));
    InMux I__701 (
            .O(N__3762),
            .I(N__3752));
    LocalMux I__700 (
            .O(N__3759),
            .I(xZ0Z_0));
    LocalMux I__699 (
            .O(N__3752),
            .I(xZ0Z_0));
    CascadeMux I__698 (
            .O(N__3747),
            .I(N__3744));
    InMux I__697 (
            .O(N__3744),
            .I(N__3739));
    InMux I__696 (
            .O(N__3743),
            .I(N__3734));
    InMux I__695 (
            .O(N__3742),
            .I(N__3734));
    LocalMux I__694 (
            .O(N__3739),
            .I(xZ0Z_1));
    LocalMux I__693 (
            .O(N__3734),
            .I(xZ0Z_1));
    CascadeMux I__692 (
            .O(N__3729),
            .I(N__3725));
    InMux I__691 (
            .O(N__3728),
            .I(N__3722));
    InMux I__690 (
            .O(N__3725),
            .I(N__3719));
    LocalMux I__689 (
            .O(N__3722),
            .I(xZ0Z_2));
    LocalMux I__688 (
            .O(N__3719),
            .I(xZ0Z_2));
    InMux I__687 (
            .O(N__3714),
            .I(un16_x_cry_1));
    CascadeMux I__686 (
            .O(N__3711),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__685 (
            .O(N__3708),
            .I(N__3698));
    InMux I__684 (
            .O(N__3707),
            .I(N__3698));
    InMux I__683 (
            .O(N__3706),
            .I(N__3695));
    InMux I__682 (
            .O(N__3705),
            .I(N__3692));
    CascadeMux I__681 (
            .O(N__3704),
            .I(N__3689));
    InMux I__680 (
            .O(N__3703),
            .I(N__3685));
    LocalMux I__679 (
            .O(N__3698),
            .I(N__3682));
    LocalMux I__678 (
            .O(N__3695),
            .I(N__3677));
    LocalMux I__677 (
            .O(N__3692),
            .I(N__3677));
    InMux I__676 (
            .O(N__3689),
            .I(N__3674));
    InMux I__675 (
            .O(N__3688),
            .I(N__3671));
    LocalMux I__674 (
            .O(N__3685),
            .I(N__3664));
    Span4Mux_h I__673 (
            .O(N__3682),
            .I(N__3664));
    Span4Mux_s0_v I__672 (
            .O(N__3677),
            .I(N__3664));
    LocalMux I__671 (
            .O(N__3674),
            .I(yZ0Z_2));
    LocalMux I__670 (
            .O(N__3671),
            .I(yZ0Z_2));
    Odrv4 I__669 (
            .O(N__3664),
            .I(yZ0Z_2));
    InMux I__668 (
            .O(N__3657),
            .I(N__3653));
    InMux I__667 (
            .O(N__3656),
            .I(N__3650));
    LocalMux I__666 (
            .O(N__3653),
            .I(un2_y_if_generate_plus_mult1_un75_sum_i_0));
    LocalMux I__665 (
            .O(N__3650),
            .I(un2_y_if_generate_plus_mult1_un75_sum_i_0));
    CascadeMux I__664 (
            .O(N__3645),
            .I(N__3641));
    InMux I__663 (
            .O(N__3644),
            .I(N__3638));
    InMux I__662 (
            .O(N__3641),
            .I(N__3635));
    LocalMux I__661 (
            .O(N__3638),
            .I(N__3630));
    LocalMux I__660 (
            .O(N__3635),
            .I(N__3630));
    Odrv4 I__659 (
            .O(N__3630),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0));
    InMux I__658 (
            .O(N__3627),
            .I(N__3624));
    LocalMux I__657 (
            .O(N__3624),
            .I(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO));
    InMux I__656 (
            .O(N__3621),
            .I(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2));
    InMux I__655 (
            .O(N__3618),
            .I(N__3615));
    LocalMux I__654 (
            .O(N__3615),
            .I(N__3611));
    InMux I__653 (
            .O(N__3614),
            .I(N__3608));
    Span4Mux_s0_v I__652 (
            .O(N__3611),
            .I(N__3603));
    LocalMux I__651 (
            .O(N__3608),
            .I(N__3603));
    Odrv4 I__650 (
            .O(N__3603),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1));
    InMux I__649 (
            .O(N__3600),
            .I(N__3597));
    LocalMux I__648 (
            .O(N__3597),
            .I(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO));
    InMux I__647 (
            .O(N__3594),
            .I(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3));
    InMux I__646 (
            .O(N__3591),
            .I(N__3588));
    LocalMux I__645 (
            .O(N__3588),
            .I(N__3585));
    Odrv4 I__644 (
            .O(N__3585),
            .I(Pixel_RNOZ0Z_4));
    InMux I__643 (
            .O(N__3582),
            .I(N__3576));
    InMux I__642 (
            .O(N__3581),
            .I(N__3569));
    InMux I__641 (
            .O(N__3580),
            .I(N__3569));
    InMux I__640 (
            .O(N__3579),
            .I(N__3569));
    LocalMux I__639 (
            .O(N__3576),
            .I(N__3564));
    LocalMux I__638 (
            .O(N__3569),
            .I(N__3564));
    Odrv12 I__637 (
            .O(N__3564),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1));
    CascadeMux I__636 (
            .O(N__3561),
            .I(N__3558));
    InMux I__635 (
            .O(N__3558),
            .I(N__3555));
    LocalMux I__634 (
            .O(N__3555),
            .I(N_49));
    InMux I__633 (
            .O(N__3552),
            .I(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4));
    InMux I__632 (
            .O(N__3549),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__631 (
            .O(N__3546),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__630 (
            .O(N__3543),
            .I(N__3539));
    InMux I__629 (
            .O(N__3542),
            .I(N__3536));
    LocalMux I__628 (
            .O(N__3539),
            .I(CounterZ0Z_13));
    LocalMux I__627 (
            .O(N__3536),
            .I(CounterZ0Z_13));
    InMux I__626 (
            .O(N__3531),
            .I(N__3527));
    InMux I__625 (
            .O(N__3530),
            .I(N__3524));
    LocalMux I__624 (
            .O(N__3527),
            .I(CounterZ0Z_12));
    LocalMux I__623 (
            .O(N__3524),
            .I(CounterZ0Z_12));
    CascadeMux I__622 (
            .O(N__3519),
            .I(un2_counterlt11_cascade_));
    InMux I__621 (
            .O(N__3516),
            .I(N__3495));
    InMux I__620 (
            .O(N__3515),
            .I(N__3495));
    InMux I__619 (
            .O(N__3514),
            .I(N__3495));
    InMux I__618 (
            .O(N__3513),
            .I(N__3486));
    InMux I__617 (
            .O(N__3512),
            .I(N__3486));
    InMux I__616 (
            .O(N__3511),
            .I(N__3486));
    InMux I__615 (
            .O(N__3510),
            .I(N__3486));
    InMux I__614 (
            .O(N__3509),
            .I(N__3477));
    InMux I__613 (
            .O(N__3508),
            .I(N__3477));
    InMux I__612 (
            .O(N__3507),
            .I(N__3477));
    InMux I__611 (
            .O(N__3506),
            .I(N__3477));
    InMux I__610 (
            .O(N__3505),
            .I(N__3468));
    InMux I__609 (
            .O(N__3504),
            .I(N__3468));
    InMux I__608 (
            .O(N__3503),
            .I(N__3468));
    InMux I__607 (
            .O(N__3502),
            .I(N__3468));
    LocalMux I__606 (
            .O(N__3495),
            .I(un2_counter_0));
    LocalMux I__605 (
            .O(N__3486),
            .I(un2_counter_0));
    LocalMux I__604 (
            .O(N__3477),
            .I(un2_counter_0));
    LocalMux I__603 (
            .O(N__3468),
            .I(un2_counter_0));
    InMux I__602 (
            .O(N__3459),
            .I(N__3455));
    InMux I__601 (
            .O(N__3458),
            .I(N__3452));
    LocalMux I__600 (
            .O(N__3455),
            .I(CounterZ0Z_4));
    LocalMux I__599 (
            .O(N__3452),
            .I(CounterZ0Z_4));
    InMux I__598 (
            .O(N__3447),
            .I(N__3443));
    InMux I__597 (
            .O(N__3446),
            .I(N__3440));
    LocalMux I__596 (
            .O(N__3443),
            .I(CounterZ0Z_0));
    LocalMux I__595 (
            .O(N__3440),
            .I(CounterZ0Z_0));
    InMux I__594 (
            .O(N__3435),
            .I(N__3431));
    InMux I__593 (
            .O(N__3434),
            .I(N__3428));
    LocalMux I__592 (
            .O(N__3431),
            .I(CounterZ0Z_3));
    LocalMux I__591 (
            .O(N__3428),
            .I(CounterZ0Z_3));
    InMux I__590 (
            .O(N__3423),
            .I(N__3419));
    InMux I__589 (
            .O(N__3422),
            .I(N__3416));
    LocalMux I__588 (
            .O(N__3419),
            .I(CounterZ0Z_2));
    LocalMux I__587 (
            .O(N__3416),
            .I(CounterZ0Z_2));
    InMux I__586 (
            .O(N__3411),
            .I(N__3407));
    InMux I__585 (
            .O(N__3410),
            .I(N__3404));
    LocalMux I__584 (
            .O(N__3407),
            .I(CounterZ0Z_1));
    LocalMux I__583 (
            .O(N__3404),
            .I(CounterZ0Z_1));
    CascadeMux I__582 (
            .O(N__3399),
            .I(N__3395));
    InMux I__581 (
            .O(N__3398),
            .I(N__3392));
    InMux I__580 (
            .O(N__3395),
            .I(N__3389));
    LocalMux I__579 (
            .O(N__3392),
            .I(CounterZ0Z_5));
    LocalMux I__578 (
            .O(N__3389),
            .I(CounterZ0Z_5));
    InMux I__577 (
            .O(N__3384),
            .I(N__3381));
    LocalMux I__576 (
            .O(N__3381),
            .I(un2_counterlto4_2));
    InMux I__575 (
            .O(N__3378),
            .I(N__3375));
    LocalMux I__574 (
            .O(N__3375),
            .I(un2_counterlt7));
    InMux I__573 (
            .O(N__3372),
            .I(N__3368));
    InMux I__572 (
            .O(N__3371),
            .I(N__3365));
    LocalMux I__571 (
            .O(N__3368),
            .I(CounterZ0Z_11));
    LocalMux I__570 (
            .O(N__3365),
            .I(CounterZ0Z_11));
    InMux I__569 (
            .O(N__3360),
            .I(N__3356));
    InMux I__568 (
            .O(N__3359),
            .I(N__3353));
    LocalMux I__567 (
            .O(N__3356),
            .I(CounterZ0Z_9));
    LocalMux I__566 (
            .O(N__3353),
            .I(CounterZ0Z_9));
    InMux I__565 (
            .O(N__3348),
            .I(N__3344));
    InMux I__564 (
            .O(N__3347),
            .I(N__3341));
    LocalMux I__563 (
            .O(N__3344),
            .I(CounterZ0Z_10));
    LocalMux I__562 (
            .O(N__3341),
            .I(CounterZ0Z_10));
    InMux I__561 (
            .O(N__3336),
            .I(N__3333));
    LocalMux I__560 (
            .O(N__3333),
            .I(un2_counterlto11_1));
    CascadeMux I__559 (
            .O(N__3330),
            .I(N_83_cascade_));
    InMux I__558 (
            .O(N__3327),
            .I(N__3324));
    LocalMux I__557 (
            .O(N__3324),
            .I(N__3319));
    CascadeMux I__556 (
            .O(N__3323),
            .I(N__3315));
    InMux I__555 (
            .O(N__3322),
            .I(N__3312));
    Span4Mux_h I__554 (
            .O(N__3319),
            .I(N__3309));
    InMux I__553 (
            .O(N__3318),
            .I(N__3304));
    InMux I__552 (
            .O(N__3315),
            .I(N__3304));
    LocalMux I__551 (
            .O(N__3312),
            .I(N_85));
    Odrv4 I__550 (
            .O(N__3309),
            .I(N_85));
    LocalMux I__549 (
            .O(N__3304),
            .I(N_85));
    CascadeMux I__548 (
            .O(N__3297),
            .I(un13lto4_i_1_cascade_));
    InMux I__547 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__546 (
            .O(N__3291),
            .I(un3_y_cry_1_THRU_CO));
    InMux I__545 (
            .O(N__3288),
            .I(un3_y_cry_1));
    InMux I__544 (
            .O(N__3285),
            .I(N__3281));
    CascadeMux I__543 (
            .O(N__3284),
            .I(N__3277));
    LocalMux I__542 (
            .O(N__3281),
            .I(N__3272));
    InMux I__541 (
            .O(N__3280),
            .I(N__3269));
    InMux I__540 (
            .O(N__3277),
            .I(N__3266));
    InMux I__539 (
            .O(N__3276),
            .I(N__3263));
    InMux I__538 (
            .O(N__3275),
            .I(N__3260));
    Span4Mux_s1_v I__537 (
            .O(N__3272),
            .I(N__3257));
    LocalMux I__536 (
            .O(N__3269),
            .I(N__3254));
    LocalMux I__535 (
            .O(N__3266),
            .I(yZ0Z_3));
    LocalMux I__534 (
            .O(N__3263),
            .I(yZ0Z_3));
    LocalMux I__533 (
            .O(N__3260),
            .I(yZ0Z_3));
    Odrv4 I__532 (
            .O(N__3257),
            .I(yZ0Z_3));
    Odrv12 I__531 (
            .O(N__3254),
            .I(yZ0Z_3));
    InMux I__530 (
            .O(N__3243),
            .I(N__3240));
    LocalMux I__529 (
            .O(N__3240),
            .I(un3_y_cry_2_THRU_CO));
    InMux I__528 (
            .O(N__3237),
            .I(un3_y_cry_2));
    InMux I__527 (
            .O(N__3234),
            .I(N__3230));
    CascadeMux I__526 (
            .O(N__3233),
            .I(N__3227));
    LocalMux I__525 (
            .O(N__3230),
            .I(N__3222));
    InMux I__524 (
            .O(N__3227),
            .I(N__3219));
    InMux I__523 (
            .O(N__3226),
            .I(N__3216));
    InMux I__522 (
            .O(N__3225),
            .I(N__3213));
    Span4Mux_s1_h I__521 (
            .O(N__3222),
            .I(N__3208));
    LocalMux I__520 (
            .O(N__3219),
            .I(N__3208));
    LocalMux I__519 (
            .O(N__3216),
            .I(yZ0Z_4));
    LocalMux I__518 (
            .O(N__3213),
            .I(yZ0Z_4));
    Odrv4 I__517 (
            .O(N__3208),
            .I(yZ0Z_4));
    InMux I__516 (
            .O(N__3201),
            .I(un3_y_cry_3));
    InMux I__515 (
            .O(N__3198),
            .I(N__3195));
    LocalMux I__514 (
            .O(N__3195),
            .I(N__3189));
    InMux I__513 (
            .O(N__3194),
            .I(N__3186));
    InMux I__512 (
            .O(N__3193),
            .I(N__3183));
    InMux I__511 (
            .O(N__3192),
            .I(N__3180));
    Span4Mux_s3_v I__510 (
            .O(N__3189),
            .I(N__3177));
    LocalMux I__509 (
            .O(N__3186),
            .I(N__3174));
    LocalMux I__508 (
            .O(N__3183),
            .I(yZ0Z_5));
    LocalMux I__507 (
            .O(N__3180),
            .I(yZ0Z_5));
    Odrv4 I__506 (
            .O(N__3177),
            .I(yZ0Z_5));
    Odrv4 I__505 (
            .O(N__3174),
            .I(yZ0Z_5));
    InMux I__504 (
            .O(N__3165),
            .I(un3_y_cry_4));
    InMux I__503 (
            .O(N__3162),
            .I(N__3154));
    InMux I__502 (
            .O(N__3161),
            .I(N__3154));
    InMux I__501 (
            .O(N__3160),
            .I(N__3151));
    InMux I__500 (
            .O(N__3159),
            .I(N__3148));
    LocalMux I__499 (
            .O(N__3154),
            .I(N__3145));
    LocalMux I__498 (
            .O(N__3151),
            .I(yZ0Z_6));
    LocalMux I__497 (
            .O(N__3148),
            .I(yZ0Z_6));
    Odrv4 I__496 (
            .O(N__3145),
            .I(yZ0Z_6));
    InMux I__495 (
            .O(N__3138),
            .I(un3_y_cry_5));
    InMux I__494 (
            .O(N__3135),
            .I(N__3132));
    LocalMux I__493 (
            .O(N__3132),
            .I(N__3126));
    InMux I__492 (
            .O(N__3131),
            .I(N__3123));
    InMux I__491 (
            .O(N__3130),
            .I(N__3120));
    InMux I__490 (
            .O(N__3129),
            .I(N__3117));
    Span4Mux_s1_h I__489 (
            .O(N__3126),
            .I(N__3114));
    LocalMux I__488 (
            .O(N__3123),
            .I(yZ0Z_7));
    LocalMux I__487 (
            .O(N__3120),
            .I(yZ0Z_7));
    LocalMux I__486 (
            .O(N__3117),
            .I(yZ0Z_7));
    Odrv4 I__485 (
            .O(N__3114),
            .I(yZ0Z_7));
    InMux I__484 (
            .O(N__3105),
            .I(un3_y_cry_6));
    InMux I__483 (
            .O(N__3102),
            .I(N__3096));
    InMux I__482 (
            .O(N__3101),
            .I(N__3093));
    InMux I__481 (
            .O(N__3100),
            .I(N__3088));
    InMux I__480 (
            .O(N__3099),
            .I(N__3088));
    LocalMux I__479 (
            .O(N__3096),
            .I(yZ0Z_8));
    LocalMux I__478 (
            .O(N__3093),
            .I(yZ0Z_8));
    LocalMux I__477 (
            .O(N__3088),
            .I(yZ0Z_8));
    InMux I__476 (
            .O(N__3081),
            .I(un3_y_cry_7));
    InMux I__475 (
            .O(N__3078),
            .I(N__3073));
    InMux I__474 (
            .O(N__3077),
            .I(N__3068));
    InMux I__473 (
            .O(N__3076),
            .I(N__3068));
    LocalMux I__472 (
            .O(N__3073),
            .I(N_130));
    LocalMux I__471 (
            .O(N__3068),
            .I(N_130));
    InMux I__470 (
            .O(N__3063),
            .I(bfn_2_6_0_));
    CascadeMux I__469 (
            .O(N__3060),
            .I(N__3057));
    InMux I__468 (
            .O(N__3057),
            .I(N__3052));
    InMux I__467 (
            .O(N__3056),
            .I(N__3047));
    InMux I__466 (
            .O(N__3055),
            .I(N__3044));
    LocalMux I__465 (
            .O(N__3052),
            .I(N__3041));
    InMux I__464 (
            .O(N__3051),
            .I(N__3036));
    InMux I__463 (
            .O(N__3050),
            .I(N__3036));
    LocalMux I__462 (
            .O(N__3047),
            .I(N__3031));
    LocalMux I__461 (
            .O(N__3044),
            .I(N__3031));
    Odrv4 I__460 (
            .O(N__3041),
            .I(yZ0Z_9));
    LocalMux I__459 (
            .O(N__3036),
            .I(yZ0Z_9));
    Odrv4 I__458 (
            .O(N__3031),
            .I(yZ0Z_9));
    InMux I__457 (
            .O(N__3024),
            .I(N__3020));
    InMux I__456 (
            .O(N__3023),
            .I(N__3017));
    LocalMux I__455 (
            .O(N__3020),
            .I(CounterZ0Z_7));
    LocalMux I__454 (
            .O(N__3017),
            .I(CounterZ0Z_7));
    InMux I__453 (
            .O(N__3012),
            .I(N__3008));
    InMux I__452 (
            .O(N__3011),
            .I(N__3005));
    LocalMux I__451 (
            .O(N__3008),
            .I(CounterZ0Z_6));
    LocalMux I__450 (
            .O(N__3005),
            .I(CounterZ0Z_6));
    CascadeMux I__449 (
            .O(N__3000),
            .I(N__2996));
    InMux I__448 (
            .O(N__2999),
            .I(N__2993));
    InMux I__447 (
            .O(N__2996),
            .I(N__2990));
    LocalMux I__446 (
            .O(N__2993),
            .I(CounterZ0Z_8));
    LocalMux I__445 (
            .O(N__2990),
            .I(CounterZ0Z_8));
    InMux I__444 (
            .O(N__2985),
            .I(N__2982));
    LocalMux I__443 (
            .O(N__2982),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0));
    InMux I__442 (
            .O(N__2979),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__441 (
            .O(N__2976),
            .I(N__2973));
    LocalMux I__440 (
            .O(N__2973),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0));
    InMux I__439 (
            .O(N__2970),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__438 (
            .O(N__2967),
            .I(N__2960));
    InMux I__437 (
            .O(N__2966),
            .I(N__2960));
    InMux I__436 (
            .O(N__2965),
            .I(N__2957));
    LocalMux I__435 (
            .O(N__2960),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0));
    LocalMux I__434 (
            .O(N__2957),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0));
    InMux I__433 (
            .O(N__2952),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_4));
    InMux I__432 (
            .O(N__2949),
            .I(N__2946));
    LocalMux I__431 (
            .O(N__2946),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO));
    InMux I__430 (
            .O(N__2943),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_5));
    CascadeMux I__429 (
            .O(N__2940),
            .I(N__2936));
    InMux I__428 (
            .O(N__2939),
            .I(N__2927));
    InMux I__427 (
            .O(N__2936),
            .I(N__2927));
    InMux I__426 (
            .O(N__2935),
            .I(N__2927));
    InMux I__425 (
            .O(N__2934),
            .I(N__2924));
    LocalMux I__424 (
            .O(N__2927),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0));
    LocalMux I__423 (
            .O(N__2924),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0));
    CascadeMux I__422 (
            .O(N__2919),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_));
    CascadeMux I__421 (
            .O(N__2916),
            .I(N__2913));
    InMux I__420 (
            .O(N__2913),
            .I(N__2910));
    LocalMux I__419 (
            .O(N__2910),
            .I(un2_y_if_generate_plus_mult1_un33_sum_i_7));
    CascadeMux I__418 (
            .O(N__2907),
            .I(N__2903));
    InMux I__417 (
            .O(N__2906),
            .I(N__2900));
    InMux I__416 (
            .O(N__2903),
            .I(N__2897));
    LocalMux I__415 (
            .O(N__2900),
            .I(N_140));
    LocalMux I__414 (
            .O(N__2897),
            .I(N_140));
    CascadeMux I__413 (
            .O(N__2892),
            .I(N__2889));
    InMux I__412 (
            .O(N__2889),
            .I(N__2886));
    LocalMux I__411 (
            .O(N__2886),
            .I(un2_y_if_generate_plus_mult1_un40_sum_i_0));
    CascadeMux I__410 (
            .O(N__2883),
            .I(N__2877));
    CascadeMux I__409 (
            .O(N__2882),
            .I(N__2874));
    CascadeMux I__408 (
            .O(N__2881),
            .I(N__2871));
    InMux I__407 (
            .O(N__2880),
            .I(N__2864));
    InMux I__406 (
            .O(N__2877),
            .I(N__2864));
    InMux I__405 (
            .O(N__2874),
            .I(N__2864));
    InMux I__404 (
            .O(N__2871),
            .I(N__2861));
    LocalMux I__403 (
            .O(N__2864),
            .I(yZ0Z_0));
    LocalMux I__402 (
            .O(N__2861),
            .I(yZ0Z_0));
    InMux I__401 (
            .O(N__2856),
            .I(N__2853));
    LocalMux I__400 (
            .O(N__2853),
            .I(un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2));
    InMux I__399 (
            .O(N__2850),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__398 (
            .O(N__2847),
            .I(N__2844));
    LocalMux I__397 (
            .O(N__2844),
            .I(un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0));
    CascadeMux I__396 (
            .O(N__2841),
            .I(N__2838));
    InMux I__395 (
            .O(N__2838),
            .I(N__2835));
    LocalMux I__394 (
            .O(N__2835),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573));
    InMux I__393 (
            .O(N__2832),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_3));
    CascadeMux I__392 (
            .O(N__2829),
            .I(N__2825));
    InMux I__391 (
            .O(N__2828),
            .I(N__2816));
    InMux I__390 (
            .O(N__2825),
            .I(N__2816));
    InMux I__389 (
            .O(N__2824),
            .I(N__2816));
    InMux I__388 (
            .O(N__2823),
            .I(N__2813));
    LocalMux I__387 (
            .O(N__2816),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12));
    LocalMux I__386 (
            .O(N__2813),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12));
    CascadeMux I__385 (
            .O(N__2808),
            .I(N__2805));
    InMux I__384 (
            .O(N__2805),
            .I(N__2802));
    LocalMux I__383 (
            .O(N__2802),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31));
    InMux I__382 (
            .O(N__2799),
            .I(N__2796));
    LocalMux I__381 (
            .O(N__2796),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3));
    InMux I__380 (
            .O(N__2793),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__379 (
            .O(N__2790),
            .I(N__2787));
    LocalMux I__378 (
            .O(N__2787),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81));
    CascadeMux I__377 (
            .O(N__2784),
            .I(N__2781));
    InMux I__376 (
            .O(N__2781),
            .I(N__2778));
    LocalMux I__375 (
            .O(N__2778),
            .I(un2_y_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__374 (
            .O(N__2775),
            .I(N__2772));
    LocalMux I__373 (
            .O(N__2772),
            .I(un2_y_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__372 (
            .O(N__2769),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__371 (
            .O(N__2766),
            .I(N__2763));
    LocalMux I__370 (
            .O(N__2763),
            .I(un2_y_if_generate_plus_mult1_un47_sum_axb_7));
    InMux I__369 (
            .O(N__2760),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__368 (
            .O(N__2757),
            .I(N__2753));
    InMux I__367 (
            .O(N__2756),
            .I(N__2744));
    InMux I__366 (
            .O(N__2753),
            .I(N__2744));
    InMux I__365 (
            .O(N__2752),
            .I(N__2744));
    InMux I__364 (
            .O(N__2751),
            .I(N__2741));
    LocalMux I__363 (
            .O(N__2744),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3));
    LocalMux I__362 (
            .O(N__2741),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3));
    CascadeMux I__361 (
            .O(N__2736),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_));
    CascadeMux I__360 (
            .O(N__2733),
            .I(N__2730));
    InMux I__359 (
            .O(N__2730),
            .I(N__2727));
    LocalMux I__358 (
            .O(N__2727),
            .I(un2_y_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__357 (
            .O(N__2724),
            .I(N__2721));
    InMux I__356 (
            .O(N__2721),
            .I(N__2718));
    LocalMux I__355 (
            .O(N__2718),
            .I(un2_y_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__354 (
            .O(N__2715),
            .I(N__2712));
    LocalMux I__353 (
            .O(N__2712),
            .I(un2_y_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__352 (
            .O(N__2709),
            .I(N__2706));
    LocalMux I__351 (
            .O(N__2706),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14));
    InMux I__350 (
            .O(N__2703),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__349 (
            .O(N__2700),
            .I(N__2697));
    InMux I__348 (
            .O(N__2697),
            .I(N__2694));
    LocalMux I__347 (
            .O(N__2694),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6));
    InMux I__346 (
            .O(N__2691),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__345 (
            .O(N__2688),
            .I(N__2685));
    LocalMux I__344 (
            .O(N__2685),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6));
    InMux I__343 (
            .O(N__2682),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__342 (
            .O(N__2679),
            .I(N__2676));
    LocalMux I__341 (
            .O(N__2676),
            .I(un2_y_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__340 (
            .O(N__2673),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__339 (
            .O(N__2670),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__338 (
            .O(N__2667),
            .I(N__2663));
    InMux I__337 (
            .O(N__2666),
            .I(N__2654));
    InMux I__336 (
            .O(N__2663),
            .I(N__2654));
    InMux I__335 (
            .O(N__2662),
            .I(N__2654));
    InMux I__334 (
            .O(N__2661),
            .I(N__2651));
    LocalMux I__333 (
            .O(N__2654),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7));
    LocalMux I__332 (
            .O(N__2651),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7));
    CascadeMux I__331 (
            .O(N__2646),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_));
    CascadeMux I__330 (
            .O(N__2643),
            .I(N__2640));
    InMux I__329 (
            .O(N__2640),
            .I(N__2637));
    LocalMux I__328 (
            .O(N__2637),
            .I(un2_y_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__327 (
            .O(N__2634),
            .I(Counter_cry_12));
    IoInMux I__326 (
            .O(N__2631),
            .I(N__2628));
    LocalMux I__325 (
            .O(N__2628),
            .I(N__2625));
    IoSpan4Mux I__324 (
            .O(N__2625),
            .I(N__2621));
    InMux I__323 (
            .O(N__2624),
            .I(N__2618));
    Odrv4 I__322 (
            .O(N__2621),
            .I(ClockVGAZ0));
    LocalMux I__321 (
            .O(N__2618),
            .I(ClockVGAZ0));
    ClkMux I__320 (
            .O(N__2613),
            .I(N__2607));
    ClkMux I__319 (
            .O(N__2612),
            .I(N__2607));
    GlobalMux I__318 (
            .O(N__2607),
            .I(N__2604));
    gio2CtrlBuf I__317 (
            .O(N__2604),
            .I(Clock12MHz_c_g));
    SRMux I__316 (
            .O(N__2601),
            .I(N__2597));
    SRMux I__315 (
            .O(N__2600),
            .I(N__2594));
    LocalMux I__314 (
            .O(N__2597),
            .I(N__2589));
    LocalMux I__313 (
            .O(N__2594),
            .I(N__2586));
    InMux I__312 (
            .O(N__2593),
            .I(N__2581));
    InMux I__311 (
            .O(N__2592),
            .I(N__2581));
    Odrv12 I__310 (
            .O(N__2589),
            .I(G_167));
    Odrv4 I__309 (
            .O(N__2586),
            .I(G_167));
    LocalMux I__308 (
            .O(N__2581),
            .I(G_167));
    InMux I__307 (
            .O(N__2574),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__306 (
            .O(N__2571),
            .I(N__2568));
    InMux I__305 (
            .O(N__2568),
            .I(N__2565));
    LocalMux I__304 (
            .O(N__2565),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0));
    InMux I__303 (
            .O(N__2562),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__302 (
            .O(N__2559),
            .I(N__2556));
    LocalMux I__301 (
            .O(N__2556),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0));
    InMux I__300 (
            .O(N__2553),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__299 (
            .O(N__2550),
            .I(N__2547));
    LocalMux I__298 (
            .O(N__2547),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0));
    CascadeMux I__297 (
            .O(N__2544),
            .I(N__2539));
    CascadeMux I__296 (
            .O(N__2543),
            .I(N__2535));
    InMux I__295 (
            .O(N__2542),
            .I(N__2531));
    InMux I__294 (
            .O(N__2539),
            .I(N__2522));
    InMux I__293 (
            .O(N__2538),
            .I(N__2522));
    InMux I__292 (
            .O(N__2535),
            .I(N__2522));
    InMux I__291 (
            .O(N__2534),
            .I(N__2522));
    LocalMux I__290 (
            .O(N__2531),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0));
    LocalMux I__289 (
            .O(N__2522),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0));
    CascadeMux I__288 (
            .O(N__2517),
            .I(N__2514));
    InMux I__287 (
            .O(N__2514),
            .I(N__2511));
    LocalMux I__286 (
            .O(N__2511),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0));
    InMux I__285 (
            .O(N__2508),
            .I(N__2505));
    LocalMux I__284 (
            .O(N__2505),
            .I(un2_y_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__283 (
            .O(N__2502),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__282 (
            .O(N__2499),
            .I(Counter_cry_3));
    InMux I__281 (
            .O(N__2496),
            .I(Counter_cry_4));
    InMux I__280 (
            .O(N__2493),
            .I(Counter_cry_5));
    InMux I__279 (
            .O(N__2490),
            .I(Counter_cry_6));
    InMux I__278 (
            .O(N__2487),
            .I(bfn_1_7_0_));
    InMux I__277 (
            .O(N__2484),
            .I(Counter_cry_8));
    InMux I__276 (
            .O(N__2481),
            .I(Counter_cry_9));
    InMux I__275 (
            .O(N__2478),
            .I(Counter_cry_10));
    InMux I__274 (
            .O(N__2475),
            .I(Counter_cry_11));
    CascadeMux I__273 (
            .O(N__2472),
            .I(un13_x_i_i_a2_0_3_cascade_));
    InMux I__272 (
            .O(N__2469),
            .I(bfn_1_6_0_));
    InMux I__271 (
            .O(N__2466),
            .I(Counter_cry_0));
    InMux I__270 (
            .O(N__2463),
            .I(Counter_cry_1));
    InMux I__269 (
            .O(N__2460),
            .I(Counter_cry_2));
    CascadeMux I__268 (
            .O(N__2457),
            .I(N__2454));
    InMux I__267 (
            .O(N__2454),
            .I(N__2451));
    LocalMux I__266 (
            .O(N__2451),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0));
    InMux I__265 (
            .O(N__2448),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__264 (
            .O(N__2445),
            .I(N__2442));
    LocalMux I__263 (
            .O(N__2442),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0));
    InMux I__262 (
            .O(N__2439),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4));
    InMux I__261 (
            .O(N__2436),
            .I(N__2433));
    LocalMux I__260 (
            .O(N__2433),
            .I(un2_y_if_generate_plus_mult1_un40_sum_axb_7));
    InMux I__259 (
            .O(N__2430),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__258 (
            .O(N__2427),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_6));
    CascadeMux I__257 (
            .O(N__2424),
            .I(N__2421));
    InMux I__256 (
            .O(N__2421),
            .I(N__2418));
    LocalMux I__255 (
            .O(N__2418),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0));
    CascadeMux I__254 (
            .O(N__2415),
            .I(N__2412));
    InMux I__253 (
            .O(N__2412),
            .I(N__2409));
    LocalMux I__252 (
            .O(N__2409),
            .I(un2_y_if_generate_plus_mult1_un33_sum_i_0));
    InMux I__251 (
            .O(N__2406),
            .I(N__2403));
    LocalMux I__250 (
            .O(N__2403),
            .I(N__2400));
    Odrv12 I__249 (
            .O(N__2400),
            .I(un13_x_i_i_a2_1));
    CascadeMux I__248 (
            .O(N__2397),
            .I(N_130_cascade_));
    InMux I__247 (
            .O(N__2394),
            .I(N__2391));
    LocalMux I__246 (
            .O(N__2391),
            .I(y_RNIA5P7Z0Z_9));
    InMux I__245 (
            .O(N__2388),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__244 (
            .O(N__2385),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__243 (
            .O(N__2382),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__242 (
            .O(N__2379),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__241 (
            .O(N__2376),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__240 (
            .O(N__2373),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_));
    InMux I__239 (
            .O(N__2370),
            .I(N__2367));
    LocalMux I__238 (
            .O(N__2367),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0));
    InMux I__237 (
            .O(N__2364),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_2));
    CascadeMux I__236 (
            .O(N__2361),
            .I(N__2358));
    InMux I__235 (
            .O(N__2358),
            .I(N__2355));
    LocalMux I__234 (
            .O(N__2355),
            .I(un2_y_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__233 (
            .O(N__2352),
            .I(N__2349));
    LocalMux I__232 (
            .O(N__2349),
            .I(un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7));
    InMux I__231 (
            .O(N__2346),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__230 (
            .O(N__2343),
            .I(N__2340));
    InMux I__229 (
            .O(N__2340),
            .I(N__2337));
    LocalMux I__228 (
            .O(N__2337),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0));
    InMux I__227 (
            .O(N__2334),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__226 (
            .O(N__2331),
            .I(N__2328));
    LocalMux I__225 (
            .O(N__2328),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0));
    InMux I__224 (
            .O(N__2325),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__223 (
            .O(N__2322),
            .I(N__2319));
    LocalMux I__222 (
            .O(N__2319),
            .I(un2_y_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__221 (
            .O(N__2316),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__220 (
            .O(N__2313),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__219 (
            .O(N__2310),
            .I(N__2305));
    InMux I__218 (
            .O(N__2309),
            .I(N__2301));
    InMux I__217 (
            .O(N__2308),
            .I(N__2294));
    InMux I__216 (
            .O(N__2305),
            .I(N__2294));
    InMux I__215 (
            .O(N__2304),
            .I(N__2294));
    LocalMux I__214 (
            .O(N__2301),
            .I(N__2291));
    LocalMux I__213 (
            .O(N__2294),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0));
    Odrv4 I__212 (
            .O(N__2291),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0));
    CascadeMux I__211 (
            .O(N__2286),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_));
    CascadeMux I__210 (
            .O(N__2283),
            .I(N__2280));
    InMux I__209 (
            .O(N__2280),
            .I(N__2277));
    LocalMux I__208 (
            .O(N__2277),
            .I(un2_y_if_generate_plus_mult1_un61_sum_i_7));
    CascadeMux I__207 (
            .O(N__2274),
            .I(N__2271));
    InMux I__206 (
            .O(N__2271),
            .I(N__2268));
    LocalMux I__205 (
            .O(N__2268),
            .I(un2_y_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__204 (
            .O(N__2265),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__203 (
            .O(N__2262),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__202 (
            .O(N__2259),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__201 (
            .O(N__2256),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__200 (
            .O(N__2253),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(un3_y_cry_8),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_1_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_5_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_1_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_6_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_1_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(un16_x_cry_8),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_1_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_1_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(Counter_cry_7),
            .carryinitout(bfn_1_7_0_));
    ICE_GB ClockVGA_derived_clock_RNIND52 (
            .USERSIGNALTOGLOBALBUFFER(N__2631),
            .GLOBALBUFFEROUTPUT(ClockVGA_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam y_RNI7THF_3_LC_1_1_0.C_ON=1'b1;
    defparam y_RNI7THF_3_LC_1_1_0.SEQ_MODE=4'b0000;
    defparam y_RNI7THF_3_LC_1_1_0.LUT_INIT=16'b1000100010001000;
    LogicCell40 y_RNI7THF_3_LC_1_1_0 (
            .in0(N__3706),
            .in1(N__3280),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un13_x_i_i_a2_1),
            .ltout(),
            .carryin(bfn_1_1_0_),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NF_LC_1_1_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NF_LC_1_1_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NF_LC_1_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NF_LC_1_1_1 (
            .in0(_gnd_net_),
            .in1(N__2304),
            .in2(N__2361),
            .in3(N__2265),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNIDS8NFZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3N_LC_1_1_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3N_LC_1_1_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3N_LC_1_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3N_LC_1_1_2 (
            .in0(_gnd_net_),
            .in1(N__2352),
            .in2(N__2310),
            .in3(N__2262),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4IC3NZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1R_LC_1_1_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1R_LC_1_1_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1R_LC_1_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1R_LC_1_1_3 (
            .in0(_gnd_net_),
            .in1(N__2308),
            .in2(N__2343),
            .in3(N__2259),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNI36E1RZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8LRER1_LC_1_1_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8LRER1_LC_1_1_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8LRER1_LC_1_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8LRER1_LC_1_1_4 (
            .in0(N__2542),
            .in1(N__2331),
            .in2(N__2283),
            .in3(N__2256),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUT_LC_1_1_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUT_LC_1_1_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUT_LC_1_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUT_LC_1_1_5 (
            .in0(_gnd_net_),
            .in1(N__2322),
            .in2(_gnd_net_),
            .in3(N__2253),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI22UUTZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_1_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_1_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3234),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_2_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_2_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3233),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNP7_LC_1_2_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNP7_LC_1_2_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNP7_LC_1_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNP7_LC_1_2_1 (
            .in0(_gnd_net_),
            .in1(N__2662),
            .in2(N__2274),
            .in3(N__2346),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNIHHNPZ0Z7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONB_LC_1_2_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONB_LC_1_2_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONB_LC_1_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONB_LC_1_2_2 (
            .in0(_gnd_net_),
            .in1(N__2709),
            .in2(N__2667),
            .in3(N__2334),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIF3ONBZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66E_LC_1_2_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66E_LC_1_2_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66E_LC_1_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66E_LC_1_2_3 (
            .in0(_gnd_net_),
            .in1(N__2666),
            .in2(N__2700),
            .in3(N__2325),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIHE66EZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHL7KT_LC_1_2_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHL7KT_LC_1_2_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHL7KT_LC_1_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHL7KT_LC_1_2_4 (
            .in0(N__2309),
            .in1(N__2688),
            .in2(N__2643),
            .in3(N__2316),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_LC_1_2_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_LC_1_2_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_LC_1_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_LC_1_2_5 (
            .in0(_gnd_net_),
            .in1(N__2679),
            .in2(_gnd_net_),
            .in3(N__2313),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0),
            .ltout(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VEZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_0_LC_1_2_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_0_LC_1_2_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_0_LC_1_2_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5Q1VE_0_LC_1_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2286),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_2_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_2_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3198),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_3_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_3_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_3_0 (
            .in0(_gnd_net_),
            .in1(N__3135),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LP_LC_1_3_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LP_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LP_LC_1_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LP_LC_1_3_1 (
            .in0(_gnd_net_),
            .in1(N__2935),
            .in2(N__2415),
            .in3(N__2388),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_sbtinv_RNIG1LPZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QD31_LC_1_3_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QD31_LC_1_3_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QD31_LC_1_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QD31_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(N__2370),
            .in2(N__2940),
            .in3(N__2385),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6QDZ0Z31),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HA81_LC_1_3_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HA81_LC_1_3_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HA81_LC_1_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HA81_LC_1_3_3 (
            .in0(_gnd_net_),
            .in1(N__2939),
            .in2(N__2457),
            .in3(N__2382),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNI5HAZ0Z81),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNI5DAA3_LC_1_3_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNI5DAA3_LC_1_3_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNI5DAA3_LC_1_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNI5DAA3_LC_1_3_4 (
            .in0(N__2823),
            .in1(N__2445),
            .in2(N__2916),
            .in3(N__2379),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_LC_1_3_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_LC_1_3_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_LC_1_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_LC_1_3_5 (
            .in0(_gnd_net_),
            .in1(N__2436),
            .in2(_gnd_net_),
            .in3(N__2376),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12),
            .ltout(un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLSZ0Z12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_0_LC_1_3_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_0_LC_1_3_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_0_LC_1_3_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_6_c_RNITLS12_0_LC_1_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2373),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_4_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(N__3099),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_4_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_4_1 (
            .in0(_gnd_net_),
            .in1(N__2394),
            .in2(N__4706),
            .in3(N__2364),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_4_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_4_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_4_2 (
            .in0(_gnd_net_),
            .in1(N__2985),
            .in2(N__4709),
            .in3(N__2448),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHF_LC_1_4_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHF_LC_1_4_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHF_LC_1_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHF_LC_1_4_3 (
            .in0(_gnd_net_),
            .in1(N__2976),
            .in2(N__4707),
            .in3(N__2439),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIFVHFZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIM3MO1_LC_1_4_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIM3MO1_LC_1_4_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIM3MO1_LC_1_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIM3MO1_LC_1_4_4 (
            .in0(N__2934),
            .in1(N__2967),
            .in2(N__2424),
            .in3(N__2430),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_1_4_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_1_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2427),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBP_LC_1_4_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBP_LC_1_4_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBP_LC_1_4_6.LUT_INIT=16'b0110011001100110;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBP_LC_1_4_6 (
            .in0(N__2965),
            .in1(N__2966),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNIIOBPZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_LC_1_4_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_LC_1_4_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_sbtinv_LC_1_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_sbtinv_LC_1_4_7 (
            .in0(N__3100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIN6QD2_0_LC_1_5_0.C_ON=1'b0;
    defparam y_RNIN6QD2_0_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam y_RNIN6QD2_0_LC_1_5_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 y_RNIN6QD2_0_LC_1_5_0 (
            .in0(N__2406),
            .in1(N__2906),
            .in2(N__2882),
            .in3(N__3051),
            .lcout(N_130),
            .ltout(N_130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_0_LC_1_5_1.C_ON=1'b0;
    defparam y_0_LC_1_5_1.SEQ_MODE=4'b1000;
    defparam y_0_LC_1_5_1.LUT_INIT=16'b0000001111001100;
    LogicCell40 y_0_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__2880),
            .in2(N__2397),
            .in3(N__4157),
            .lcout(yZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4471),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIA5P7_9_LC_1_5_2.C_ON=1'b0;
    defparam y_RNIA5P7_9_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam y_RNIA5P7_9_LC_1_5_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 y_RNIA5P7_9_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3050),
            .lcout(y_RNIA5P7Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_2_LC_1_5_3.C_ON=1'b0;
    defparam y_2_LC_1_5_3.SEQ_MODE=4'b1000;
    defparam y_2_LC_1_5_3.LUT_INIT=16'b0001001011110000;
    LogicCell40 y_2_LC_1_5_3 (
            .in0(N__3294),
            .in1(N__3076),
            .in2(N__3704),
            .in3(N__4158),
            .lcout(yZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4471),
            .ce(),
            .sr(_gnd_net_));
    defparam y_1_LC_1_5_4.C_ON=1'b0;
    defparam y_1_LC_1_5_4.SEQ_MODE=4'b1000;
    defparam y_1_LC_1_5_4.LUT_INIT=16'b0101111110100000;
    LogicCell40 y_1_LC_1_5_4 (
            .in0(N__4156),
            .in1(_gnd_net_),
            .in2(N__2883),
            .in3(N__3318),
            .lcout(N_85),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4471),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIO44V_1_LC_1_5_5.C_ON=1'b0;
    defparam y_RNIO44V_1_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam y_RNIO44V_1_LC_1_5_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 y_RNIO44V_1_LC_1_5_5 (
            .in0(N__3192),
            .in1(N__3159),
            .in2(N__3323),
            .in3(N__3101),
            .lcout(),
            .ltout(un13_x_i_i_a2_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNI58ME1_4_LC_1_5_6.C_ON=1'b0;
    defparam y_RNI58ME1_4_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam y_RNI58ME1_4_LC_1_5_6.LUT_INIT=16'b0000000000110000;
    LogicCell40 y_RNI58ME1_4_LC_1_5_6 (
            .in0(_gnd_net_),
            .in1(N__3225),
            .in2(N__2472),
            .in3(N__3130),
            .lcout(N_140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_3_LC_1_5_7.C_ON=1'b0;
    defparam y_3_LC_1_5_7.SEQ_MODE=4'b1000;
    defparam y_3_LC_1_5_7.LUT_INIT=16'b0001001011110000;
    LogicCell40 y_3_LC_1_5_7 (
            .in0(N__3243),
            .in1(N__3077),
            .in2(N__3284),
            .in3(N__4159),
            .lcout(yZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4471),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_0_LC_1_6_0.C_ON=1'b1;
    defparam Counter_0_LC_1_6_0.SEQ_MODE=4'b1010;
    defparam Counter_0_LC_1_6_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_0_LC_1_6_0 (
            .in0(N__3510),
            .in1(N__3447),
            .in2(_gnd_net_),
            .in3(N__2469),
            .lcout(CounterZ0Z_0),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(Counter_cry_0),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_1_LC_1_6_1.C_ON=1'b1;
    defparam Counter_1_LC_1_6_1.SEQ_MODE=4'b1010;
    defparam Counter_1_LC_1_6_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_1_LC_1_6_1 (
            .in0(N__3502),
            .in1(N__3411),
            .in2(_gnd_net_),
            .in3(N__2466),
            .lcout(CounterZ0Z_1),
            .ltout(),
            .carryin(Counter_cry_0),
            .carryout(Counter_cry_1),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_2_LC_1_6_2.C_ON=1'b1;
    defparam Counter_2_LC_1_6_2.SEQ_MODE=4'b1010;
    defparam Counter_2_LC_1_6_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_2_LC_1_6_2 (
            .in0(N__3511),
            .in1(N__3423),
            .in2(_gnd_net_),
            .in3(N__2463),
            .lcout(CounterZ0Z_2),
            .ltout(),
            .carryin(Counter_cry_1),
            .carryout(Counter_cry_2),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_3_LC_1_6_3.C_ON=1'b1;
    defparam Counter_3_LC_1_6_3.SEQ_MODE=4'b1010;
    defparam Counter_3_LC_1_6_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_3_LC_1_6_3 (
            .in0(N__3503),
            .in1(N__3435),
            .in2(_gnd_net_),
            .in3(N__2460),
            .lcout(CounterZ0Z_3),
            .ltout(),
            .carryin(Counter_cry_2),
            .carryout(Counter_cry_3),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_4_LC_1_6_4.C_ON=1'b1;
    defparam Counter_4_LC_1_6_4.SEQ_MODE=4'b1010;
    defparam Counter_4_LC_1_6_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_4_LC_1_6_4 (
            .in0(N__3512),
            .in1(N__3459),
            .in2(_gnd_net_),
            .in3(N__2499),
            .lcout(CounterZ0Z_4),
            .ltout(),
            .carryin(Counter_cry_3),
            .carryout(Counter_cry_4),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_5_LC_1_6_5.C_ON=1'b1;
    defparam Counter_5_LC_1_6_5.SEQ_MODE=4'b1010;
    defparam Counter_5_LC_1_6_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_5_LC_1_6_5 (
            .in0(N__3504),
            .in1(N__3398),
            .in2(_gnd_net_),
            .in3(N__2496),
            .lcout(CounterZ0Z_5),
            .ltout(),
            .carryin(Counter_cry_4),
            .carryout(Counter_cry_5),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_6_LC_1_6_6.C_ON=1'b1;
    defparam Counter_6_LC_1_6_6.SEQ_MODE=4'b1010;
    defparam Counter_6_LC_1_6_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_6_LC_1_6_6 (
            .in0(N__3513),
            .in1(N__3012),
            .in2(_gnd_net_),
            .in3(N__2493),
            .lcout(CounterZ0Z_6),
            .ltout(),
            .carryin(Counter_cry_5),
            .carryout(Counter_cry_6),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_7_LC_1_6_7.C_ON=1'b1;
    defparam Counter_7_LC_1_6_7.SEQ_MODE=4'b1010;
    defparam Counter_7_LC_1_6_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_7_LC_1_6_7 (
            .in0(N__3505),
            .in1(N__3024),
            .in2(_gnd_net_),
            .in3(N__2490),
            .lcout(CounterZ0Z_7),
            .ltout(),
            .carryin(Counter_cry_6),
            .carryout(Counter_cry_7),
            .clk(N__2613),
            .ce(),
            .sr(N__2601));
    defparam Counter_8_LC_1_7_0.C_ON=1'b1;
    defparam Counter_8_LC_1_7_0.SEQ_MODE=4'b1010;
    defparam Counter_8_LC_1_7_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_8_LC_1_7_0 (
            .in0(N__3516),
            .in1(N__2999),
            .in2(_gnd_net_),
            .in3(N__2487),
            .lcout(CounterZ0Z_8),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(Counter_cry_8),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Counter_9_LC_1_7_1.C_ON=1'b1;
    defparam Counter_9_LC_1_7_1.SEQ_MODE=4'b1010;
    defparam Counter_9_LC_1_7_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_9_LC_1_7_1 (
            .in0(N__3507),
            .in1(N__3360),
            .in2(_gnd_net_),
            .in3(N__2484),
            .lcout(CounterZ0Z_9),
            .ltout(),
            .carryin(Counter_cry_8),
            .carryout(Counter_cry_9),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Counter_10_LC_1_7_2.C_ON=1'b1;
    defparam Counter_10_LC_1_7_2.SEQ_MODE=4'b1010;
    defparam Counter_10_LC_1_7_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_10_LC_1_7_2 (
            .in0(N__3514),
            .in1(N__3348),
            .in2(_gnd_net_),
            .in3(N__2481),
            .lcout(CounterZ0Z_10),
            .ltout(),
            .carryin(Counter_cry_9),
            .carryout(Counter_cry_10),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Counter_11_LC_1_7_3.C_ON=1'b1;
    defparam Counter_11_LC_1_7_3.SEQ_MODE=4'b1010;
    defparam Counter_11_LC_1_7_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_11_LC_1_7_3 (
            .in0(N__3506),
            .in1(N__3372),
            .in2(_gnd_net_),
            .in3(N__2478),
            .lcout(CounterZ0Z_11),
            .ltout(),
            .carryin(Counter_cry_10),
            .carryout(Counter_cry_11),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Counter_12_LC_1_7_4.C_ON=1'b1;
    defparam Counter_12_LC_1_7_4.SEQ_MODE=4'b1010;
    defparam Counter_12_LC_1_7_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_12_LC_1_7_4 (
            .in0(N__3515),
            .in1(N__3531),
            .in2(_gnd_net_),
            .in3(N__2475),
            .lcout(CounterZ0Z_12),
            .ltout(),
            .carryin(Counter_cry_11),
            .carryout(Counter_cry_12),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Counter_13_LC_1_7_5.C_ON=1'b0;
    defparam Counter_13_LC_1_7_5.SEQ_MODE=4'b1010;
    defparam Counter_13_LC_1_7_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 Counter_13_LC_1_7_5 (
            .in0(N__3508),
            .in1(N__3543),
            .in2(_gnd_net_),
            .in3(N__2634),
            .lcout(CounterZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam ClockVGA_LC_1_7_6.C_ON=1'b0;
    defparam ClockVGA_LC_1_7_6.SEQ_MODE=4'b1010;
    defparam ClockVGA_LC_1_7_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 ClockVGA_LC_1_7_6 (
            .in0(_gnd_net_),
            .in1(N__2624),
            .in2(_gnd_net_),
            .in3(N__3509),
            .lcout(ClockVGAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2612),
            .ce(),
            .sr(N__2600));
    defparam Reset_latch_LC_1_8_0.C_ON=1'b0;
    defparam Reset_latch_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam Reset_latch_LC_1_8_0.LUT_INIT=16'b0000000011100100;
    LogicCell40 Reset_latch_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(N__2592),
            .in2(_gnd_net_),
            .in3(N__2593),
            .lcout(G_167),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_1_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_1_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_1_0 (
            .in0(_gnd_net_),
            .in1(N__3705),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_1_0_),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCU_LC_2_1_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCU_LC_2_1_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCU_LC_2_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCU_LC_2_1_1 (
            .in0(_gnd_net_),
            .in1(N__2715),
            .in2(N__2543),
            .in3(N__2574),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIFQFCUZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1ND1_LC_2_1_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1ND1_LC_2_1_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1ND1_LC_2_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1ND1_LC_2_1_2 (
            .in0(_gnd_net_),
            .in1(N__2538),
            .in2(N__2571),
            .in3(N__2562),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNIRD1NDZ0Z1),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_4_LC_2_1_3.C_ON=1'b1;
    defparam Pixel_RNO_4_LC_2_1_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_4_LC_2_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_4_LC_2_1_3 (
            .in0(_gnd_net_),
            .in1(N__2559),
            .in2(N__2544),
            .in3(N__2553),
            .lcout(Pixel_RNOZ0Z_4),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_1_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_1_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_1_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_1_4 (
            .in0(_gnd_net_),
            .in1(N__2550),
            .in2(N__2517),
            .in3(N__2534),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFR1_LC_2_1_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFR1_LC_2_1_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFR1_LC_2_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFR1_LC_2_1_5 (
            .in0(_gnd_net_),
            .in1(N__2508),
            .in2(_gnd_net_),
            .in3(N__2502),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNINAPFRZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_1_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_1_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3285),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_2_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_2_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_2_2_0 (
            .in0(_gnd_net_),
            .in1(N__3194),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2O14_LC_2_2_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2O14_LC_2_2_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2O14_LC_2_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2O14_LC_2_2_1 (
            .in0(_gnd_net_),
            .in1(N__2752),
            .in2(N__2724),
            .in3(N__2703),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIQ2OZ0Z14),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5G6_LC_2_2_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5G6_LC_2_2_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5G6_LC_2_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5G6_LC_2_2_2 (
            .in0(_gnd_net_),
            .in1(N__2856),
            .in2(N__2757),
            .in3(N__2691),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIRB5GZ0Z6),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3V6_LC_2_2_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3V6_LC_2_2_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3V6_LC_2_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3V6_LC_2_2_3 (
            .in0(_gnd_net_),
            .in1(N__2756),
            .in2(N__2841),
            .in3(N__2682),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNILM3VZ0Z6),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNIR1SME_LC_2_2_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNIR1SME_LC_2_2_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNIR1SME_LC_2_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNIR1SME_LC_2_2_4 (
            .in0(N__2661),
            .in1(N__2799),
            .in2(N__2733),
            .in3(N__2673),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_LC_2_2_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_LC_2_2_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_LC_2_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_LC_2_2_5 (
            .in0(_gnd_net_),
            .in1(N__2775),
            .in2(_gnd_net_),
            .in3(N__2670),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7),
            .ltout(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETDZ0Z7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_0_LC_2_2_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_0_LC_2_2_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_0_LC_2_2_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIEETD7_0_LC_2_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2646),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_3_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_3_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_3_0 (
            .in0(_gnd_net_),
            .in1(N__3161),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8O2_LC_2_3_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8O2_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8O2_LC_2_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8O2_LC_2_3_1 (
            .in0(_gnd_net_),
            .in1(N__2824),
            .in2(N__2892),
            .in3(N__2850),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIVE8OZ0Z2),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNION573_LC_2_3_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNION573_LC_2_3_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNION573_LC_2_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNION573_LC_2_3_2 (
            .in0(_gnd_net_),
            .in1(N__2847),
            .in2(N__2829),
            .in3(N__2832),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNIONZ0Z573),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVG3_LC_2_3_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVG3_LC_2_3_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVG3_LC_2_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVG3_LC_2_3_3 (
            .in0(_gnd_net_),
            .in1(N__2828),
            .in2(N__2808),
            .in3(N__2793),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIFIVGZ0Z3),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI2VUB7_LC_2_3_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI2VUB7_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI2VUB7_LC_2_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI2VUB7_LC_2_3_4 (
            .in0(N__2751),
            .in1(N__2790),
            .in2(N__2784),
            .in3(N__2769),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_LC_2_3_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_LC_2_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_LC_2_3_5 (
            .in0(_gnd_net_),
            .in1(N__2766),
            .in2(_gnd_net_),
            .in3(N__2760),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3),
            .ltout(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1MZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_0_LC_2_3_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_0_LC_2_3_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_0_LC_2_3_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIJJ1M3_0_LC_2_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2736),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_3_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_3_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_3_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_3_7 (
            .in0(N__3162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_4_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_4_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_4_0 (
            .in0(_gnd_net_),
            .in1(N__3055),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(un2_y_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJC_LC_2_4_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJC_LC_2_4_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJC_LC_2_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJC_LC_2_4_1 (
            .in0(_gnd_net_),
            .in1(N__4688),
            .in2(N__4708),
            .in3(N__2979),
            .lcout(un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_RNI7OJCZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKC_LC_2_4_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKC_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKC_LC_2_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKC_LC_2_4_2 (
            .in0(_gnd_net_),
            .in1(N__4699),
            .in2(_gnd_net_),
            .in3(N__2970),
            .lcout(un2_y_if_generate_plus_mult1_un26_sum_cry_3_c_RNI8QKCZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLC_LC_2_4_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLC_LC_2_4_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLC_LC_2_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLC_LC_2_4_3 (
            .in0(_gnd_net_),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__2952),
            .lcout(un2_y_if_generate_plus_mult1_un26_sum_cry_4_c_RNI9SLCZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un26_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un26_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_LC_2_4_4.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_LC_2_4_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_LC_2_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_LC_2_4_4 (
            .in0(_gnd_net_),
            .in1(N__2949),
            .in2(_gnd_net_),
            .in3(N__2943),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0),
            .ltout(un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MFZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_0_LC_2_4_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_0_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_0_LC_2_4_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_6_c_RNIJ7MF_0_LC_2_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2919),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIMA162_9_LC_2_4_6.C_ON=1'b0;
    defparam y_RNIMA162_9_LC_2_4_6.SEQ_MODE=4'b0000;
    defparam y_RNIMA162_9_LC_2_4_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 y_RNIMA162_9_LC_2_4_6 (
            .in0(N__3056),
            .in1(N__3688),
            .in2(N__2907),
            .in3(N__3275),
            .lcout(y_RNIMA162Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_4_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_4_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3129),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un3_y_cry_1_c_LC_2_5_0.C_ON=1'b1;
    defparam un3_y_cry_1_c_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam un3_y_cry_1_c_LC_2_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un3_y_cry_1_c_LC_2_5_0 (
            .in0(_gnd_net_),
            .in1(N__3322),
            .in2(N__2881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(un3_y_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un3_y_cry_1_THRU_LUT4_0_LC_2_5_1.C_ON=1'b1;
    defparam un3_y_cry_1_THRU_LUT4_0_LC_2_5_1.SEQ_MODE=4'b0000;
    defparam un3_y_cry_1_THRU_LUT4_0_LC_2_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un3_y_cry_1_THRU_LUT4_0_LC_2_5_1 (
            .in0(_gnd_net_),
            .in1(N__3703),
            .in2(_gnd_net_),
            .in3(N__3288),
            .lcout(un3_y_cry_1_THRU_CO),
            .ltout(),
            .carryin(un3_y_cry_1),
            .carryout(un3_y_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un3_y_cry_2_THRU_LUT4_0_LC_2_5_2.C_ON=1'b1;
    defparam un3_y_cry_2_THRU_LUT4_0_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam un3_y_cry_2_THRU_LUT4_0_LC_2_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un3_y_cry_2_THRU_LUT4_0_LC_2_5_2 (
            .in0(_gnd_net_),
            .in1(N__3276),
            .in2(_gnd_net_),
            .in3(N__3237),
            .lcout(un3_y_cry_2_THRU_CO),
            .ltout(),
            .carryin(un3_y_cry_2),
            .carryout(un3_y_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_4_LC_2_5_3.C_ON=1'b1;
    defparam y_4_LC_2_5_3.SEQ_MODE=4'b1000;
    defparam y_4_LC_2_5_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_4_LC_2_5_3 (
            .in0(N__4160),
            .in1(N__3226),
            .in2(_gnd_net_),
            .in3(N__3201),
            .lcout(yZ0Z_4),
            .ltout(),
            .carryin(un3_y_cry_3),
            .carryout(un3_y_cry_4),
            .clk(N__4473),
            .ce(),
            .sr(_gnd_net_));
    defparam y_5_LC_2_5_4.C_ON=1'b1;
    defparam y_5_LC_2_5_4.SEQ_MODE=4'b1000;
    defparam y_5_LC_2_5_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_5_LC_2_5_4 (
            .in0(N__4163),
            .in1(N__3193),
            .in2(_gnd_net_),
            .in3(N__3165),
            .lcout(yZ0Z_5),
            .ltout(),
            .carryin(un3_y_cry_4),
            .carryout(un3_y_cry_5),
            .clk(N__4473),
            .ce(),
            .sr(_gnd_net_));
    defparam y_6_LC_2_5_5.C_ON=1'b1;
    defparam y_6_LC_2_5_5.SEQ_MODE=4'b1000;
    defparam y_6_LC_2_5_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_6_LC_2_5_5 (
            .in0(N__4161),
            .in1(N__3160),
            .in2(_gnd_net_),
            .in3(N__3138),
            .lcout(yZ0Z_6),
            .ltout(),
            .carryin(un3_y_cry_5),
            .carryout(un3_y_cry_6),
            .clk(N__4473),
            .ce(),
            .sr(_gnd_net_));
    defparam y_7_LC_2_5_6.C_ON=1'b1;
    defparam y_7_LC_2_5_6.SEQ_MODE=4'b1000;
    defparam y_7_LC_2_5_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_7_LC_2_5_6 (
            .in0(N__4164),
            .in1(N__3131),
            .in2(_gnd_net_),
            .in3(N__3105),
            .lcout(yZ0Z_7),
            .ltout(),
            .carryin(un3_y_cry_6),
            .carryout(un3_y_cry_7),
            .clk(N__4473),
            .ce(),
            .sr(_gnd_net_));
    defparam y_8_LC_2_5_7.C_ON=1'b1;
    defparam y_8_LC_2_5_7.SEQ_MODE=4'b1000;
    defparam y_8_LC_2_5_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_8_LC_2_5_7 (
            .in0(N__4162),
            .in1(N__3102),
            .in2(_gnd_net_),
            .in3(N__3081),
            .lcout(yZ0Z_8),
            .ltout(),
            .carryin(un3_y_cry_7),
            .carryout(un3_y_cry_8),
            .clk(N__4473),
            .ce(),
            .sr(_gnd_net_));
    defparam y_9_LC_2_6_0.C_ON=1'b0;
    defparam y_9_LC_2_6_0.SEQ_MODE=4'b1000;
    defparam y_9_LC_2_6_0.LUT_INIT=16'b0011010001110000;
    LogicCell40 y_9_LC_2_6_0 (
            .in0(N__3078),
            .in1(N__4134),
            .in2(N__3060),
            .in3(N__3063),
            .lcout(yZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4472),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_RNICJ474_6_LC_2_6_1.C_ON=1'b0;
    defparam Counter_RNICJ474_6_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam Counter_RNICJ474_6_LC_2_6_1.LUT_INIT=16'b0000111100000111;
    LogicCell40 Counter_RNICJ474_6_LC_2_6_1 (
            .in0(N__3023),
            .in1(N__3011),
            .in2(N__3000),
            .in3(N__3378),
            .lcout(),
            .ltout(un2_counterlt11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_RNI7QMJ6_13_LC_2_6_2.C_ON=1'b0;
    defparam Counter_RNI7QMJ6_13_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam Counter_RNI7QMJ6_13_LC_2_6_2.LUT_INIT=16'b1000101010001000;
    LogicCell40 Counter_RNI7QMJ6_13_LC_2_6_2 (
            .in0(N__3542),
            .in1(N__3530),
            .in2(N__3519),
            .in3(N__3336),
            .lcout(un2_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_RNIVB1D1_0_LC_2_6_3.C_ON=1'b0;
    defparam Counter_RNIVB1D1_0_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam Counter_RNIVB1D1_0_LC_2_6_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 Counter_RNIVB1D1_0_LC_2_6_3 (
            .in0(N__3458),
            .in1(N__3446),
            .in2(_gnd_net_),
            .in3(N__3434),
            .lcout(un2_counterlto4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_RNIVO2Q2_1_LC_2_6_4.C_ON=1'b0;
    defparam Counter_RNIVO2Q2_1_LC_2_6_4.SEQ_MODE=4'b0000;
    defparam Counter_RNIVO2Q2_1_LC_2_6_4.LUT_INIT=16'b0000011100001111;
    LogicCell40 Counter_RNIVO2Q2_1_LC_2_6_4 (
            .in0(N__3422),
            .in1(N__3410),
            .in2(N__3399),
            .in3(N__3384),
            .lcout(un2_counterlt7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Counter_RNI4CPD1_9_LC_2_7_2.C_ON=1'b0;
    defparam Counter_RNI4CPD1_9_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam Counter_RNI4CPD1_9_LC_2_7_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 Counter_RNI4CPD1_9_LC_2_7_2 (
            .in0(N__3371),
            .in1(N__3359),
            .in2(_gnd_net_),
            .in3(N__3347),
            .lcout(un2_counterlto11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_11_LC_4_1_1.C_ON=1'b0;
    defparam Pixel_RNO_11_LC_4_1_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_11_LC_4_1_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 Pixel_RNO_11_LC_4_1_1 (
            .in0(N__3627),
            .in1(N__3644),
            .in2(_gnd_net_),
            .in3(N__3579),
            .lcout(),
            .ltout(N_83_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_9_LC_4_1_2.C_ON=1'b0;
    defparam Pixel_RNO_9_LC_4_1_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_9_LC_4_1_2.LUT_INIT=16'b0011111110011111;
    LogicCell40 Pixel_RNO_9_LC_4_1_2 (
            .in0(N__3580),
            .in1(N__3614),
            .in2(N__3330),
            .in3(N__3600),
            .lcout(),
            .ltout(un13lto4_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_5_LC_4_1_3.C_ON=1'b0;
    defparam Pixel_RNO_5_LC_4_1_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_5_LC_4_1_3.LUT_INIT=16'b1111011111111101;
    LogicCell40 Pixel_RNO_5_LC_4_1_3 (
            .in0(N__3327),
            .in1(N__3708),
            .in2(N__3297),
            .in3(N__3581),
            .lcout(N_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_1_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_1_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_1_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_inv_LC_4_1_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_inv_LC_4_1_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_inv_LC_4_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_inv_LC_4_1_5 (
            .in0(_gnd_net_),
            .in1(N__3657),
            .in2(N__3711),
            .in3(N__3707),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_LC_5_1_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_LC_5_1_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_LC_5_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_c_LC_5_1_0 (
            .in0(_gnd_net_),
            .in1(N__3656),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_1_0_),
            .carryout(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_LUT4_0_LC_5_1_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_LUT4_0_LC_5_1_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_LUT4_0_LC_5_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_LUT4_0_LC_5_1_1 (
            .in0(_gnd_net_),
            .in1(N__4642),
            .in2(N__3645),
            .in3(N__3621),
            .lcout(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2_THRU_CO),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_LUT4_0_LC_5_1_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_LUT4_0_LC_5_1_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_LUT4_0_LC_5_1_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_LUT4_0_LC_5_1_2 (
            .in0(_gnd_net_),
            .in1(N__3618),
            .in2(N__4662),
            .in3(N__3594),
            .lcout(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3_THRU_CO),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un1_rem_adjust_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_0_LC_5_1_3.C_ON=1'b0;
    defparam Pixel_RNO_0_LC_5_1_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_0_LC_5_1_3.LUT_INIT=16'b1010111101101111;
    LogicCell40 Pixel_RNO_0_LC_5_1_3 (
            .in0(N__3591),
            .in1(N__3582),
            .in2(N__3561),
            .in3(N__3552),
            .lcout(N_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_2_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_2_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_2_0 (
            .in0(_gnd_net_),
            .in1(N__4215),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_5_2_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_5_2_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_5_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_5_2_1 (
            .in0(_gnd_net_),
            .in1(N__3788),
            .in2(N__3774),
            .in3(N__3549),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_6_LC_5_2_2.C_ON=1'b1;
    defparam Pixel_RNO_6_LC_5_2_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_6_LC_5_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_6_LC_5_2_2 (
            .in0(_gnd_net_),
            .in1(N__3897),
            .in2(N__3864),
            .in3(N__3546),
            .lcout(Pixel_RNOZ0Z_6),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_2_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_2_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_2_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_2_3 (
            .in0(_gnd_net_),
            .in1(N__3789),
            .in2(N__3888),
            .in3(N__3859),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_5_2_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_5_2_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_5_2_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_5_2_4 (
            .in0(_gnd_net_),
            .in1(N__3876),
            .in2(_gnd_net_),
            .in3(N__3780),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0),
            .ltout(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_10_LC_5_2_5.C_ON=1'b0;
    defparam Pixel_RNO_10_LC_5_2_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_10_LC_5_2_5.LUT_INIT=16'b1111111110100101;
    LogicCell40 Pixel_RNO_10_LC_5_2_5 (
            .in0(N__4216),
            .in1(_gnd_net_),
            .in2(N__3777),
            .in3(N__3834),
            .lcout(N_57),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI5UL6_5_LC_5_2_7.C_ON=1'b0;
    defparam x_RNI5UL6_5_LC_5_2_7.SEQ_MODE=4'b0000;
    defparam x_RNI5UL6_5_LC_5_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI5UL6_5_LC_5_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4278),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI6ANQ_1_LC_5_3_1.C_ON=1'b0;
    defparam x_RNI6ANQ_1_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam x_RNI6ANQ_1_LC_5_3_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 x_RNI6ANQ_1_LC_5_3_1 (
            .in0(N__3742),
            .in1(N__3762),
            .in2(N__3729),
            .in3(N__3832),
            .lcout(un11_x_0_a2_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_0_LC_5_3_5.C_ON=1'b0;
    defparam x_0_LC_5_3_5.SEQ_MODE=4'b1000;
    defparam x_0_LC_5_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_0_LC_5_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3763),
            .lcout(xZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4476),
            .ce(),
            .sr(_gnd_net_));
    defparam x_1_LC_5_3_6.C_ON=1'b0;
    defparam x_1_LC_5_3_6.SEQ_MODE=4'b1000;
    defparam x_1_LC_5_3_6.LUT_INIT=16'b1010010101011010;
    LogicCell40 x_1_LC_5_3_6 (
            .in0(N__3764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3743),
            .lcout(xZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4476),
            .ce(),
            .sr(_gnd_net_));
    defparam un16_x_cry_1_c_LC_5_4_0.C_ON=1'b1;
    defparam un16_x_cry_1_c_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam un16_x_cry_1_c_LC_5_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un16_x_cry_1_c_LC_5_4_0 (
            .in0(_gnd_net_),
            .in1(N__3765),
            .in2(N__3747),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(un16_x_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_2_LC_5_4_1.C_ON=1'b1;
    defparam x_2_LC_5_4_1.SEQ_MODE=4'b1000;
    defparam x_2_LC_5_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_2_LC_5_4_1 (
            .in0(_gnd_net_),
            .in1(N__3728),
            .in2(_gnd_net_),
            .in3(N__3714),
            .lcout(xZ0Z_2),
            .ltout(),
            .carryin(un16_x_cry_1),
            .carryout(un16_x_cry_2),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_3_LC_5_4_2.C_ON=1'b1;
    defparam x_3_LC_5_4_2.SEQ_MODE=4'b1000;
    defparam x_3_LC_5_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_3_LC_5_4_2 (
            .in0(_gnd_net_),
            .in1(N__3833),
            .in2(_gnd_net_),
            .in3(N__3813),
            .lcout(N_89),
            .ltout(),
            .carryin(un16_x_cry_2),
            .carryout(un16_x_cry_3),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_4_LC_5_4_3.C_ON=1'b1;
    defparam x_4_LC_5_4_3.SEQ_MODE=4'b1000;
    defparam x_4_LC_5_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_4_LC_5_4_3 (
            .in0(_gnd_net_),
            .in1(N__4214),
            .in2(_gnd_net_),
            .in3(N__3810),
            .lcout(xZ0Z_4),
            .ltout(),
            .carryin(un16_x_cry_3),
            .carryout(un16_x_cry_4),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_5_LC_5_4_4.C_ON=1'b1;
    defparam x_5_LC_5_4_4.SEQ_MODE=4'b1000;
    defparam x_5_LC_5_4_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 x_5_LC_5_4_4 (
            .in0(N__4133),
            .in1(N__4276),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(xZ0Z_5),
            .ltout(),
            .carryin(un16_x_cry_4),
            .carryout(un16_x_cry_5),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_6_LC_5_4_5.C_ON=1'b1;
    defparam x_6_LC_5_4_5.SEQ_MODE=4'b1000;
    defparam x_6_LC_5_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_6_LC_5_4_5 (
            .in0(_gnd_net_),
            .in1(N__4245),
            .in2(_gnd_net_),
            .in3(N__3804),
            .lcout(xZ0Z_6),
            .ltout(),
            .carryin(un16_x_cry_5),
            .carryout(un16_x_cry_6),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_7_LC_5_4_6.C_ON=1'b1;
    defparam x_7_LC_5_4_6.SEQ_MODE=4'b1000;
    defparam x_7_LC_5_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_7_LC_5_4_6 (
            .in0(_gnd_net_),
            .in1(N__4435),
            .in2(_gnd_net_),
            .in3(N__3801),
            .lcout(xZ0Z_7),
            .ltout(),
            .carryin(un16_x_cry_6),
            .carryout(un16_x_cry_7),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_8_LC_5_4_7.C_ON=1'b1;
    defparam x_8_LC_5_4_7.SEQ_MODE=4'b1000;
    defparam x_8_LC_5_4_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 x_8_LC_5_4_7 (
            .in0(N__4117),
            .in1(N__4546),
            .in2(_gnd_net_),
            .in3(N__3798),
            .lcout(xZ0Z_8),
            .ltout(),
            .carryin(un16_x_cry_7),
            .carryout(un16_x_cry_8),
            .clk(N__4475),
            .ce(),
            .sr(_gnd_net_));
    defparam x_9_LC_5_5_0.C_ON=1'b0;
    defparam x_9_LC_5_5_0.SEQ_MODE=4'b1000;
    defparam x_9_LC_5_5_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 x_9_LC_5_5_0 (
            .in0(N__4089),
            .in1(N__4118),
            .in2(_gnd_net_),
            .in3(N__3795),
            .lcout(xZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4474),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_LC_6_1_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_LC_6_1_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_LC_6_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_LC_6_1_0 (
            .in0(_gnd_net_),
            .in1(N__3845),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_1_0_),
            .carryout(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_LUT4_0_LC_6_1_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_LUT4_0_LC_6_1_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_LUT4_0_LC_6_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_LUT4_0_LC_6_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3966),
            .in3(N__3792),
            .lcout(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_THRU_CO),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_1_LC_6_1_2.C_ON=1'b0;
    defparam Pixel_RNO_1_LC_6_1_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_1_LC_6_1_2.LUT_INIT=16'b1100111101101111;
    LogicCell40 Pixel_RNO_1_LC_6_1_2 (
            .in0(N__3954),
            .in1(N__3975),
            .in2(N__3930),
            .in3(N__3969),
            .lcout(N_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_7_LC_6_1_3.C_ON=1'b0;
    defparam Pixel_RNO_7_LC_6_1_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_7_LC_6_1_3.LUT_INIT=16'b1001010111111111;
    LogicCell40 Pixel_RNO_7_LC_6_1_3 (
            .in0(N__3962),
            .in1(N__3953),
            .in2(N__3945),
            .in3(N__3936),
            .lcout(N_59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_6_1_7.C_ON=1'b0;
    defparam PixelZ0_LC_6_1_7.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_6_1_7.LUT_INIT=16'b0000000100000100;
    LogicCell40 PixelZ0_LC_6_1_7 (
            .in0(N__4311),
            .in1(N__3921),
            .in2(N__4323),
            .in3(N__3915),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4479),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_6_2_0 (
            .in0(_gnd_net_),
            .in1(N__4277),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_6_2_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_6_2_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_6_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_6_2_1 (
            .in0(_gnd_net_),
            .in1(N__4001),
            .in2(N__3993),
            .in3(N__3891),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_6_2_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_6_2_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_6_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_6_2_2 (
            .in0(_gnd_net_),
            .in1(N__4017),
            .in2(N__4053),
            .in3(N__3879),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_6_2_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_6_2_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_6_2_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_6_2_3 (
            .in0(N__3863),
            .in1(N__4002),
            .in2(N__4041),
            .in3(N__3870),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_6_2_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_6_2_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_6_2_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_6_2_4 (
            .in0(_gnd_net_),
            .in1(N__4029),
            .in2(_gnd_net_),
            .in3(N__3867),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_inv_LC_6_2_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_inv_LC_6_2_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_inv_LC_6_2_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_x_if_generate_plus_mult1_un1_rem_adjust_cry_4_c_inv_LC_6_2_5 (
            .in0(N__3846),
            .in1(N__4687),
            .in2(_gnd_net_),
            .in3(N__4217),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_3_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(N__4240),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_3_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_3_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_3_1 (
            .in0(_gnd_net_),
            .in1(N__4349),
            .in2(N__3984),
            .in3(N__4044),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_3_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(N__4365),
            .in2(N__4401),
            .in3(N__4032),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_3_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_3_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_3_3 (
            .in0(N__4016),
            .in1(N__4350),
            .in2(N__4389),
            .in3(N__4023),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_3_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_3_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_3_4 (
            .in0(_gnd_net_),
            .in1(N__4377),
            .in2(_gnd_net_),
            .in3(N__4020),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2),
            .ltout(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_3_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_3_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4005),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI6VL6_6_LC_6_3_6.C_ON=1'b0;
    defparam x_RNI6VL6_6_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam x_RNI6VL6_6_LC_6_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI6VL6_6_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI70M6_7_LC_6_3_7.C_ON=1'b0;
    defparam x_RNI70M6_7_LC_6_3_7.SEQ_MODE=4'b0000;
    defparam x_RNI70M6_7_LC_6_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI70M6_7_LC_6_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4432),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_3_LC_6_4_0.C_ON=1'b0;
    defparam Pixel_RNO_3_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_3_LC_6_4_0.LUT_INIT=16'b1010100000010101;
    LogicCell40 Pixel_RNO_3_LC_6_4_0 (
            .in0(N__4087),
            .in1(N__4434),
            .in2(N__4287),
            .in3(N__4547),
            .lcout(Pixel_0_sqmuxa_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI92M6_9_LC_6_4_1.C_ON=1'b0;
    defparam x_RNI92M6_9_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam x_RNI92M6_9_LC_6_4_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI92M6_9_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4085),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_2_LC_6_4_3.C_ON=1'b0;
    defparam Pixel_RNO_2_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_2_LC_6_4_3.LUT_INIT=16'b1110101010101010;
    LogicCell40 Pixel_RNO_2_LC_6_4_3 (
            .in0(N__4502),
            .in1(N__4551),
            .in2(N__4179),
            .in3(N__4088),
            .lcout(Pixel_0_sqmuxa_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSyncZ0_LC_6_4_4.C_ON=1'b0;
    defparam HSyncZ0_LC_6_4_4.SEQ_MODE=4'b1000;
    defparam HSyncZ0_LC_6_4_4.LUT_INIT=16'b1111111111111000;
    LogicCell40 HSyncZ0_LC_6_4_4 (
            .in0(N__4275),
            .in1(N__4244),
            .in2(N__4442),
            .in3(N__4062),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4477),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_8_LC_6_4_5.C_ON=1'b0;
    defparam Pixel_RNO_8_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_8_LC_6_4_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 Pixel_RNO_8_LC_6_4_5 (
            .in0(N__4243),
            .in1(N__4213),
            .in2(_gnd_net_),
            .in3(N__4274),
            .lcout(N_90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNIMQNQ_4_LC_6_4_6.C_ON=1'b0;
    defparam x_RNIMQNQ_4_LC_6_4_6.SEQ_MODE=4'b0000;
    defparam x_RNIMQNQ_4_LC_6_4_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 x_RNIMQNQ_4_LC_6_4_6 (
            .in0(N__4273),
            .in1(N__4242),
            .in2(N__4218),
            .in3(N__4433),
            .lcout(),
            .ltout(un11_x_0_a2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNID8R22_9_LC_6_4_7.C_ON=1'b0;
    defparam x_RNID8R22_9_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam x_RNID8R22_9_LC_6_4_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 x_RNID8R22_9_LC_6_4_7 (
            .in0(N__4175),
            .in1(N__4550),
            .in2(N__4167),
            .in3(N__4086),
            .lcout(x_RNID8R22Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_RNO_0_LC_6_5_0.C_ON=1'b1;
    defparam HSync_RNO_0_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam HSync_RNO_0_LC_6_5_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 HSync_RNO_0_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(N__4084),
            .in2(_gnd_net_),
            .in3(N__4545),
            .lcout(un1_xlto9_i_0),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(un2_x_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_6_5_1.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_6_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4056),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_6_5_2.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_6_5_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4446),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__4443),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_7_3_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_7_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__4580),
            .in2(N__4512),
            .in3(N__4392),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_7_3_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_7_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__4596),
            .in2(N__4335),
            .in3(N__4380),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_7_3_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_7_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_7_3_3 (
            .in0(N__4364),
            .in1(N__4581),
            .in2(N__4620),
            .in3(N__4371),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_7_3_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_7_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__4608),
            .in2(_gnd_net_),
            .in3(N__4368),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1),
            .ltout(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_7_3_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_7_3_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_7_3_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_7_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4353),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_4_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_7_4_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_7_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__4341),
            .in2(_gnd_net_),
            .in3(N__4326),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_7_4_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__4716),
            .in2(N__4710),
            .in3(N__4611),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_7_4_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_7_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_7_4_3 (
            .in0(N__4595),
            .in1(N__4557),
            .in2(N__4572),
            .in3(N__4602),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_7_4_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_7_4_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4599),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0),
            .ltout(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_7_4_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_7_4_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_7_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4584),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_7_4_6.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_7_4_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_7_4_6 (
            .in0(_gnd_net_),
            .in1(N__4567),
            .in2(_gnd_net_),
            .in3(N__4568),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI81M6_8_LC_7_4_7.C_ON=1'b0;
    defparam x_RNI81M6_8_LC_7_4_7.SEQ_MODE=4'b0000;
    defparam x_RNI81M6_8_LC_7_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 x_RNI81M6_8_LC_7_4_7 (
            .in0(N__4549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSyncZ0_LC_8_4_3.C_ON=1'b0;
    defparam VSyncZ0_LC_8_4_3.SEQ_MODE=4'b1000;
    defparam VSyncZ0_LC_8_4_3.LUT_INIT=16'b0011001100110011;
    LogicCell40 VSyncZ0_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(N__4503),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4478),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
