-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 24 2015 16:35:13

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSync : out std_logic;
    SCLK1 : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic;
    nCS2 : out std_logic;
    SDATA2 : out std_logic;
    SCLK2 : out std_logic;
    Clock12MHz : in std_logic;
    nCS1 : out std_logic;
    SDATA1 : in std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \font_un3_pixel_29_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_18_cascade_\ : std_logic;
signal \N_1214_0_cascade_\ : std_logic;
signal g1 : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\ : std_logic;
signal charx_i_24 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3\ : std_logic;
signal charx_i_23 : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal un18_beamylto9_2 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_axb_3_i : std_logic;
signal \g1_2_cascade_\ : std_logic;
signal \g2_3_0_cascade_\ : std_logic;
signal g2_2_0 : std_logic;
signal \g3_3_cascade_\ : std_logic;
signal \g0_0_2_cascade_\ : std_logic;
signal \g0_3_cascade_\ : std_logic;
signal \N_21_0\ : std_logic;
signal \Pixel_RNOZ0Z_37\ : std_logic;
signal \font_un126_pixel_m_2_1_1_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_71\ : std_logic;
signal g0_0_1 : std_logic;
signal font_un3_pixel_29 : std_logic;
signal \font_un126_pixel_m_2_1_cascade_\ : std_logic;
signal g2_2_0_1 : std_logic;
signal \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\ : std_logic;
signal font_un126_pixel_5_a0_2 : std_logic;
signal \G_19_i_a11_0_1_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_36\ : std_logic;
signal \g1_1_0_0_cascade_\ : std_logic;
signal g0_0 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \un13_beamylt7_0_cascade_\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un3_beamx_5 : std_logic;
signal un3_beamx_7 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_i_5 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7 : std_logic;
signal \g2_1_cascade_\ : std_logic;
signal \N_7_cascade_\ : std_logic;
signal g2_1 : std_logic;
signal \g0_1_0_cascade_\ : std_logic;
signal \g0_1_3_cascade_\ : std_logic;
signal \g3_2_2_cascade_\ : std_logic;
signal \N_20\ : std_logic;
signal \g0_4_cascade_\ : std_logic;
signal \G_21_i_2\ : std_logic;
signal \Pixel_c\ : std_logic;
signal g1_1_0 : std_logic;
signal g0_2_0 : std_logic;
signal \g1_1_cascade_\ : std_logic;
signal g3_1 : std_logic;
signal g0_5 : std_logic;
signal g1_0_0 : std_logic;
signal g0_0_a3_0 : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \N_35\ : std_logic;
signal \N_58_mux\ : std_logic;
signal charx_if_generate_plus_mult1_un1_sum_axb1 : std_logic;
signal \beamY_RNIDQG2Z0Z_0_cascade_\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\ : std_logic;
signal \beamY_RNINKIU27Z0Z_0\ : std_logic;
signal \beamY_RNINKIU27Z0Z_0_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_29_cascade_\ : std_logic;
signal \N_10\ : std_logic;
signal chessboardpixel_un152_pixel_27 : std_logic;
signal chessboardpixel_un174_pixellt10 : std_logic;
signal chessboardpixel_un175_pixel : std_logic;
signal g1_2_1 : std_logic;
signal \chessboardpixel_un175_pixel_cascade_\ : std_logic;
signal g2_3_0_0 : std_logic;
signal un13_beamylt7 : std_logic;
signal un15_beamy : std_logic;
signal un18_beamylt10_0 : std_logic;
signal un15_beamy_2 : std_logic;
signal \Pixel_RNOZ0Z_44_cascade_\ : std_logic;
signal \N_10_0_0\ : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un1_beamx_2 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \HSync_c\ : std_logic;
signal un4_row : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_3_l_ofx : std_logic;
signal \column_1_if_generate_plus_mult1_un47_sum_c5_iZ0\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_4_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal un5_visiblex_i_26 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \un4_row_9_2_cascade_\ : std_logic;
signal un4_row_9_5 : std_logic;
signal un4_row_9_0 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \column_1_if_generate_plus_mult1_un47_sum_cZ0Z5\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_axb_3 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8 : std_logic;
signal \Pixel_RNOZ0Z_14\ : std_logic;
signal font_un126_pixel_5_a0_1 : std_logic;
signal \N_1740_0\ : std_logic;
signal \font_un28_pixel_29_cascade_\ : std_logic;
signal \beamY_RNIDA2GGA3Z0Z_0\ : std_logic;
signal g0_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\ : std_logic;
signal \beamY_RNIDA2GGA3Z0Z_0_cascade_\ : std_logic;
signal \N_19_0_0\ : std_logic;
signal font_un28_pixel_30 : std_logic;
signal font_un28_pixel_29 : std_logic;
signal \N_15_i\ : std_logic;
signal \Pixel_RNOZ0Z_28_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_9\ : std_logic;
signal chary_24 : std_logic;
signal \chary_1_24_cascade_\ : std_logic;
signal \N_1737_0\ : std_logic;
signal \chary_1_0_24_cascade_\ : std_logic;
signal \g2_3_cascade_\ : std_logic;
signal g1_1_1 : std_logic;
signal un116_pixel_0_0_0 : std_logic;
signal \N_5_1\ : std_logic;
signal g0_0_a3_4 : std_logic;
signal \un8_beamylto9_1_cascade_\ : std_logic;
signal un8_beamy : std_logic;
signal \N_134_0\ : std_logic;
signal g4_1 : std_logic;
signal g0_0_a3_5 : std_logic;
signal \m4_rn_1_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_40\ : std_logic;
signal \content_content_ram0__RNIR1C2R81Z0Z_0_cascade_\ : std_logic;
signal \N_331_i\ : std_logic;
signal \un4_row_m7_ns_1_cascade_\ : std_logic;
signal \beamY_RNIPAQ91Z0Z_6\ : std_logic;
signal un4_beamy_0 : std_logic;
signal m4_sn : std_logic;
signal \content_content_ram0__RNIR1C2R81_0Z0Z_0\ : std_logic;
signal un6_rowlt7_0 : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal un5_visiblex_i_27 : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \if_generate_plus_mult1_un61_sum_s_5_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal chary_2_24 : std_logic;
signal \beamY_RNI539IG9Z0Z_3\ : std_logic;
signal \beamY_RNI539IG9Z0Z_3_cascade_\ : std_logic;
signal g4 : std_logic;
signal chary_0_24 : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_axbxc5_1 : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_\ : std_logic;
signal g1_2_0 : std_logic;
signal \beamY_RNIMSO1N7_0Z0Z_2_cascade_\ : std_logic;
signal g4_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0 : std_logic;
signal \g2_1_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_0_5 : std_logic;
signal \Pixel_RNOZ0Z_66\ : std_logic;
signal un5_visibley_0_28 : std_logic;
signal g2 : std_logic;
signal un5_visibley_0_29 : std_logic;
signal \Pixel_RNOZ0Z_67\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal un4_beamylt8_0 : std_logic;
signal \GB_BUFFER_Clock12MHz_c_g_THRU_CO\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal \G_383\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal un6_rowlto0 : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_iZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal content_column_1_i_2_i_2 : std_logic;
signal un6_rowlto1 : std_logic;
signal \content_N_25\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \content_column_1_i_2_2_cascade_\ : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal if_generate_plus_mult1_un75_sum_axb_4_l_fx : std_logic;
signal chessboardpixel_un152_pixel_24 : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal \content_m7_ns_1_cascade_\ : std_logic;
signal \content_N_8\ : std_logic;
signal \content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_\ : std_logic;
signal \content_content_ram7__RNI6B0NG3Z0Z_0\ : std_logic;
signal \content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0\ : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_2_5 : std_logic;
signal un5_visibley_2_29 : std_logic;
signal g2_0_0 : std_logic;
signal \beamY_RNIMSO1N7Z0Z_2\ : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_1_0_5 : std_logic;
signal g2_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1 : std_logic;
signal \g2_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_1_5 : std_logic;
signal \VSync_c\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3 : std_logic;
signal un5_visibley_3_28 : std_logic;
signal \un5_visibley_3_28_cascade_\ : std_logic;
signal \g1_3_cascade_\ : std_logic;
signal g2_0_1 : std_logic;
signal un1_beamylto9_2 : std_logic;
signal un5_visibley_1_28 : std_logic;
signal \chessboardpixel_un200_pixellto4_1_cascade_\ : std_logic;
signal chessboardpixel_un200_pixellt10 : std_logic;
signal un8_beamy_3 : std_logic;
signal \beamY_i_2_cascade_\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0\ : std_logic;
signal chessboardpixel_un178_pixel_26 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_cZ0Z5\ : std_logic;
signal \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axbxc5 : std_logic;
signal \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\ : std_logic;
signal \content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_\ : std_logic;
signal \content_content_ram9__e_0_RNIFBHPN1Z0Z_0\ : std_logic;
signal \content_content_ram5__RNIEM2QF3Z0Z_0\ : std_logic;
signal content_ram9_0 : std_logic;
signal content_ram11_0 : std_logic;
signal \nCS1_c\ : std_logic;
signal un5_visibley_2_28 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0 : std_logic;
signal \beamY_RNIVMI9D5Z0Z_3\ : std_logic;
signal un5_visibley_1_29 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c4 : std_logic;
signal \beamY_RNI8325Z0Z_6_cascade_\ : std_logic;
signal \un5_visibley_c5_cascade_\ : std_logic;
signal un1_beamylto9_1 : std_logic;
signal \un5_visibley_c3_cascade_\ : std_logic;
signal \un5_beamx_2_0_cascade_\ : std_logic;
signal un5_beamx_3 : std_logic;
signal \un5_visibley_ac0_11_0_1_cascade_\ : std_logic;
signal \beamY_RNI8325_0Z0Z_6\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \CO4_1\ : std_logic;
signal \row_1_if_generate_plus_mult1_un47_sum_cZ0Z5\ : std_logic;
signal content_ram8_0 : std_logic;
signal \content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_\ : std_logic;
signal \content_N_19\ : std_logic;
signal content_column_1_i_2_2 : std_logic;
signal if_generate_plus_mult1_un61_sum_s_5 : std_logic;
signal \content_content_ram10__e_0_RNIOLNMN1Z0Z_0\ : std_logic;
signal content_ram3_0 : std_logic;
signal content_awe9 : std_logic;
signal content_ram0_0 : std_logic;
signal content_awe8 : std_logic;
signal content_awe11 : std_logic;
signal content_ram5_0 : std_logic;
signal content_ram12_0 : std_logic;
signal content_awe0_0_a2_0 : std_logic;
signal \content_awe0_0_a2_0_cascade_\ : std_logic;
signal content_ram4_0 : std_logic;
signal \content_N_36\ : std_logic;
signal \content_N_36_cascade_\ : std_logic;
signal \content_awe7_1_cascade_\ : std_logic;
signal content_ram6_0 : std_logic;
signal content_awe7_1 : std_logic;
signal content_ram7_0 : std_logic;
signal \nCS1_0_sqmuxa\ : std_logic;
signal \un19_slaveselectlt5_0_cascade_\ : std_logic;
signal un19_slaveselectlt5_0 : std_logic;
signal \counter_RNI4HQB1Z0Z_5_cascade_\ : std_logic;
signal \beamY_RNI4FVGVZ0Z_4_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal \N_596_2\ : std_logic;
signal \un5_visibley_4_28_cascade_\ : std_logic;
signal un5_visibley_3_29 : std_logic;
signal \g1_8_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axb4_i : std_logic;
signal g1_3_0 : std_logic;
signal un5_visibley_1_0_28 : std_logic;
signal \beamY_RNIJ0H2Z0Z_4_cascade_\ : std_logic;
signal un5_visibley_c5 : std_logic;
signal un5_visibley_c6_0_0_0 : std_logic;
signal \un5_visibley_c6_0_0_0_cascade_\ : std_logic;
signal un5_visibley_c3 : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal g2_1_1_0 : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \beamY_RNI9DLCZ0Z_1\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal content_ram10_0 : std_logic;
signal content_awe10 : std_logic;
signal \content_N_35_cascade_\ : std_logic;
signal content_awe3_1 : std_logic;
signal \content_awe3_1_cascade_\ : std_logic;
signal content_ram2_0 : std_logic;
signal \content_N_40\ : std_logic;
signal \content_N_35\ : std_logic;
signal \content_awe1_0_a2_0_cascade_\ : std_logic;
signal content_ram1_0 : std_logic;
signal \un7_slaveselectlt5_cascade_\ : std_logic;
signal \N_190_i\ : std_logic;
signal un1_counter_0_1 : std_logic;
signal un7_slaveselectlt5 : std_logic;
signal \un1_counter_0_1_cascade_\ : std_logic;
signal \slaveselect_1lto5_0_cascade_\ : std_logic;
signal slaveselect_1lto5_1 : std_logic;
signal \SCLK1_0_i\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal un7_slaveselectlt2_0 : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal counter_cry_1 : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal counter_cry_2 : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal counter_cry_3 : std_logic;
signal \counter_RNI4HQB1Z0Z_5\ : std_logic;
signal counter_cry_4 : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal \SDATA1_c\ : std_logic;
signal \slaveselectZ0\ : std_logic;
signal un5_slaveselect : std_logic;
signal \SDATA2_c\ : std_logic;
signal \Clock12MHz_c_g\ : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_\ : std_logic;
signal \beamY_RNII78UPZ0Z_4\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axbxc5_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c4 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axb3 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc5_1 : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_c5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum : std_logic;
signal \beamY_RNIFC5HAZ0Z_4\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axbxc5_1 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_ac0_8 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axbxc5_2 : std_logic;
signal \chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axb4 : std_logic;
signal \beamY_RNI65RM4_0Z0Z_9\ : std_logic;
signal \beamY_RNIJNLCZ0Z_9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_c4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \beamY_RNIQ7DB_0Z0Z_9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal chary_if_generate_plus_mult1_un33_sum_axb3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \beamY_RNITSR8_0Z0Z_8\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \Clock12MHz_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \SDATA2_wire\ : std_logic;
signal \nCS1_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \SCLK1_wire\ : std_logic;
signal \SCLK2_wire\ : std_logic;
signal \nCS2_wire\ : std_logic;
signal \SDATA1_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \Clock12MHz_wire\ <= Clock12MHz;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    SDATA2 <= \SDATA2_wire\;
    nCS1 <= \nCS1_wire\;
    Pixel <= \Pixel_wire\;
    SCLK1 <= \SCLK1_wire\;
    SCLK2 <= \SCLK2_wire\;
    nCS2 <= \nCS2_wire\;
    \SDATA1_wire\ <= SDATA1;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__10363\,
            RESETB => \N__15601\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \Clock12MHz_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__15818\,
            GLOBALBUFFEROUTPUT => \Clock12MHz_c_g\
        );

    \Clock12MHz_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15820\,
            DIN => \N__15819\,
            DOUT => \N__15818\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15820\,
            PADOUT => \N__15819\,
            PADIN => \N__15818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15809\,
            DIN => \N__15808\,
            DOUT => \N__15807\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15809\,
            PADOUT => \N__15808\,
            PADIN => \N__15807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10753\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15800\,
            DIN => \N__15799\,
            DOUT => \N__15798\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15800\,
            PADOUT => \N__15799\,
            PADIN => \N__15798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8353\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDATA2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15791\,
            DIN => \N__15790\,
            DOUT => \N__15789\,
            PACKAGEPIN => \SDATA2_wire\
        );

    \SDATA2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15791\,
            PADOUT => \N__15790\,
            PADIN => \N__15789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14374\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15782\,
            DIN => \N__15781\,
            DOUT => \N__15780\,
            PACKAGEPIN => \nCS1_wire\
        );

    \nCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15782\,
            PADOUT => \N__15781\,
            PADIN => \N__15780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15773\,
            DIN => \N__15772\,
            DOUT => \N__15771\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15773\,
            PADOUT => \N__15772\,
            PADIN => \N__15771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8035\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15764\,
            DIN => \N__15763\,
            DOUT => \N__15762\,
            PACKAGEPIN => \SCLK1_wire\
        );

    \SCLK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15764\,
            PADOUT => \N__15763\,
            PADIN => \N__15762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15755\,
            DIN => \N__15754\,
            DOUT => \N__15753\,
            PACKAGEPIN => \SCLK2_wire\
        );

    \SCLK2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15755\,
            PADOUT => \N__15754\,
            PADIN => \N__15753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14133\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15746\,
            DIN => \N__15745\,
            DOUT => \N__15744\,
            PACKAGEPIN => \nCS2_wire\
        );

    \nCS2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15746\,
            PADOUT => \N__15745\,
            PADIN => \N__15744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDATA1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15737\,
            DIN => \N__15736\,
            DOUT => \N__15735\,
            PACKAGEPIN => \SDATA1_wire\
        );

    \SDATA1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15737\,
            PADOUT => \N__15736\,
            PADIN => \N__15735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SDATA1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3653\ : InMux
    port map (
            O => \N__15718\,
            I => \N__15713\
        );

    \I__3652\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15710\
        );

    \I__3651\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15701\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15696\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__15710\,
            I => \N__15696\
        );

    \I__3648\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15693\
        );

    \I__3647\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15690\
        );

    \I__3646\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15683\
        );

    \I__3645\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15683\
        );

    \I__3644\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15683\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15680\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__15701\,
            I => \N__15677\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__15696\,
            I => \N__15672\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__15693\,
            I => \N__15672\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__15690\,
            I => \N__15667\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__15683\,
            I => \N__15667\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__15680\,
            I => \N__15662\
        );

    \I__3636\ : Span4Mux_s3_h
    port map (
            O => \N__15677\,
            I => \N__15662\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__15672\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__3634\ : Odrv4
    port map (
            O => \N__15667\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__15662\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__3632\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15652\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__15652\,
            I => \beamY_RNITSR8_0Z0Z_8\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__3629\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__15643\,
            I => \N__15640\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__15640\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0\
        );

    \I__3626\ : InMux
    port map (
            O => \N__15637\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__15634\,
            I => \N__15631\
        );

    \I__3624\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15628\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15628\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0\
        );

    \I__3622\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15622\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15619\
        );

    \I__3620\ : Odrv12
    port map (
            O => \N__15619\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0\
        );

    \I__3619\ : InMux
    port map (
            O => \N__15616\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__3618\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15610\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__15610\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__15607\,
            I => \N__15603\
        );

    \I__3615\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15593\
        );

    \I__3614\ : InMux
    port map (
            O => \N__15603\,
            I => \N__15588\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15588\
        );

    \I__3612\ : IoInMux
    port map (
            O => \N__15601\,
            I => \N__15582\
        );

    \I__3611\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15579\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__15599\,
            I => \N__15576\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__15598\,
            I => \N__15572\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__15597\,
            I => \N__15569\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__15596\,
            I => \N__15566\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__15593\,
            I => \N__15561\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__15588\,
            I => \N__15561\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__15587\,
            I => \N__15558\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__15586\,
            I => \N__15555\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__15585\,
            I => \N__15552\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__15582\,
            I => \N__15547\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__15579\,
            I => \N__15544\
        );

    \I__3599\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15537\
        );

    \I__3598\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15537\
        );

    \I__3597\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15537\
        );

    \I__3596\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15534\
        );

    \I__3595\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15531\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__15561\,
            I => \N__15528\
        );

    \I__3593\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15525\
        );

    \I__3592\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15522\
        );

    \I__3591\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15519\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__15551\,
            I => \N__15516\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__15550\,
            I => \N__15513\
        );

    \I__3588\ : Span4Mux_s3_v
    port map (
            O => \N__15547\,
            I => \N__15510\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__15544\,
            I => \N__15507\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__15537\,
            I => \N__15504\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__15534\,
            I => \N__15493\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15493\
        );

    \I__3583\ : Sp12to4
    port map (
            O => \N__15528\,
            I => \N__15493\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__15525\,
            I => \N__15493\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15493\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__15519\,
            I => \N__15490\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15487\
        );

    \I__3578\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15484\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__15510\,
            I => \N__15480\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__15507\,
            I => \N__15477\
        );

    \I__3575\ : Span12Mux_s6_h
    port map (
            O => \N__15504\,
            I => \N__15474\
        );

    \I__3574\ : Span12Mux_s8_v
    port map (
            O => \N__15493\,
            I => \N__15465\
        );

    \I__3573\ : Span12Mux_s7_v
    port map (
            O => \N__15490\,
            I => \N__15465\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15465\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15465\
        );

    \I__3570\ : InMux
    port map (
            O => \N__15483\,
            I => \N__15462\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__15480\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__15477\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3567\ : Odrv12
    port map (
            O => \N__15474\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__15465\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__15462\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__3563\ : InMux
    port map (
            O => \N__15448\,
            I => \N__15445\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__15445\,
            I => \N__15442\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__15442\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15439\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__15436\,
            I => \N__15433\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15430\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__15430\,
            I => \N__15427\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__15427\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__3555\ : InMux
    port map (
            O => \N__15424\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__3554\ : InMux
    port map (
            O => \N__15421\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__15418\,
            I => \N__15413\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__15417\,
            I => \N__15409\
        );

    \I__3551\ : InMux
    port map (
            O => \N__15416\,
            I => \N__15397\
        );

    \I__3550\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15397\
        );

    \I__3549\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15397\
        );

    \I__3548\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15397\
        );

    \I__3547\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15397\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__15397\,
            I => \N__15394\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__15394\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\
        );

    \I__3544\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__3543\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15385\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__15385\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__3541\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15379\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__15379\,
            I => \N__15374\
        );

    \I__3539\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15369\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15369\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__15374\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__15369\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__3535\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15358\
        );

    \I__3534\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15358\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__15358\,
            I => chary_if_generate_plus_mult1_un47_sum_axbxc5_2
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__15355\,
            I => \chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_\
        );

    \I__3531\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__3530\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15346\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__15346\,
            I => chary_if_generate_plus_mult1_un47_sum_axb4
        );

    \I__3528\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15337\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15337\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__15337\,
            I => \N__15332\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15327\
        );

    \I__3524\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15327\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__15332\,
            I => \beamY_RNI65RM4_0Z0Z_9\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__15327\,
            I => \beamY_RNI65RM4_0Z0Z_9\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__15322\,
            I => \N__15316\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__15321\,
            I => \N__15313\
        );

    \I__3519\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15304\
        );

    \I__3518\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15304\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15304\
        );

    \I__3516\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15304\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__15304\,
            I => \N__15301\
        );

    \I__3514\ : Span4Mux_s3_h
    port map (
            O => \N__15301\,
            I => \N__15298\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__15298\,
            I => \beamY_RNIJNLCZ0Z_9\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__15295\,
            I => \N__15286\
        );

    \I__3511\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15281\
        );

    \I__3510\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15281\
        );

    \I__3509\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15275\
        );

    \I__3508\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15275\
        );

    \I__3507\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15268\
        );

    \I__3506\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15268\
        );

    \I__3505\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15265\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__15281\,
            I => \N__15262\
        );

    \I__3503\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15259\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__15275\,
            I => \N__15256\
        );

    \I__3501\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15253\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15250\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__15268\,
            I => \N__15245\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__15265\,
            I => \N__15245\
        );

    \I__3497\ : Span4Mux_s3_h
    port map (
            O => \N__15262\,
            I => \N__15242\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__15259\,
            I => \N__15239\
        );

    \I__3495\ : Span4Mux_s3_h
    port map (
            O => \N__15256\,
            I => \N__15232\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__15253\,
            I => \N__15232\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__15250\,
            I => \N__15232\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__15245\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__15242\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__15239\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__15232\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__3488\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15217\
        );

    \I__3487\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15217\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__15217\,
            I => chary_if_generate_plus_mult1_un47_sum_c4
        );

    \I__3485\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15211\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15208\
        );

    \I__3483\ : Span4Mux_s2_h
    port map (
            O => \N__15208\,
            I => \N__15205\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__15205\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\
        );

    \I__3481\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15199\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__15199\,
            I => \beamY_RNIQ7DB_0Z0Z_9\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15196\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__3478\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15185\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__15192\,
            I => \N__15182\
        );

    \I__3476\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15176\
        );

    \I__3475\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15173\
        );

    \I__3474\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15168\
        );

    \I__3473\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15168\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__15185\,
            I => \N__15165\
        );

    \I__3471\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15162\
        );

    \I__3470\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15155\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15155\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15179\,
            I => \N__15155\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__15176\,
            I => \N__15148\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15148\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15148\
        );

    \I__3464\ : Span4Mux_s3_h
    port map (
            O => \N__15165\,
            I => \N__15145\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__15162\,
            I => \N__15140\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__15155\,
            I => \N__15140\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__15148\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__15145\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3459\ : Odrv12
    port map (
            O => \N__15140\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__3458\ : InMux
    port map (
            O => \N__15133\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__3457\ : InMux
    port map (
            O => \N__15130\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__15127\,
            I => \N__15124\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15116\
        );

    \I__3454\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15116\
        );

    \I__3453\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15109\
        );

    \I__3452\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15106\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__15116\,
            I => \N__15103\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15096\
        );

    \I__3449\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15096\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15096\
        );

    \I__3447\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15093\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__15109\,
            I => \N__15088\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N__15088\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__15103\,
            I => \N__15083\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__15096\,
            I => \N__15083\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__15093\,
            I => \N__15080\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__15088\,
            I => \N__15075\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__15083\,
            I => \N__15075\
        );

    \I__3439\ : Span4Mux_s2_h
    port map (
            O => \N__15080\,
            I => \N__15072\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__15075\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__15072\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__3436\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15064\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__15064\,
            I => \N__15060\
        );

    \I__3434\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15053\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__15060\,
            I => \N__15049\
        );

    \I__3432\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15044\
        );

    \I__3431\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15044\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15039\
        );

    \I__3429\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15039\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__15036\
        );

    \I__3427\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15033\
        );

    \I__3426\ : Span4Mux_h
    port map (
            O => \N__15049\,
            I => \N__15030\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__15044\,
            I => \N__15025\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__15039\,
            I => \N__15025\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__15036\,
            I => \N__15020\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__15020\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__15030\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__15025\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__15020\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__3418\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15010\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__15010\,
            I => chary_if_generate_plus_mult1_un61_sum_c4
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__15007\,
            I => \N__15003\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__15006\,
            I => \N__15000\
        );

    \I__3414\ : InMux
    port map (
            O => \N__15003\,
            I => \N__14995\
        );

    \I__3413\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14995\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__14995\,
            I => \N__14992\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__14992\,
            I => chary_if_generate_plus_mult1_un47_sum_axb3
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__14986\,
            I => \N__14978\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__14985\,
            I => \N__14975\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__14984\,
            I => \N__14971\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__14983\,
            I => \N__14968\
        );

    \I__3405\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14959\
        );

    \I__3404\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14959\
        );

    \I__3403\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14959\
        );

    \I__3402\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14954\
        );

    \I__3401\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14954\
        );

    \I__3400\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14943\
        );

    \I__3399\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14943\
        );

    \I__3398\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14940\
        );

    \I__3397\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14937\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__14959\,
            I => \N__14932\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__14954\,
            I => \N__14932\
        );

    \I__3394\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14923\
        );

    \I__3393\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14923\
        );

    \I__3392\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14923\
        );

    \I__3391\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14923\
        );

    \I__3390\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14918\
        );

    \I__3389\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14918\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__14943\,
            I => \N__14914\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14911\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__14937\,
            I => \N__14904\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__14932\,
            I => \N__14904\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14904\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__14918\,
            I => \N__14901\
        );

    \I__3382\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14898\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__14914\,
            I => \N__14893\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__14911\,
            I => \N__14893\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__14904\,
            I => \N__14890\
        );

    \I__3378\ : Odrv12
    port map (
            O => \N__14901\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__14898\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__14893\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__14890\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__14881\,
            I => \N__14876\
        );

    \I__3373\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14868\
        );

    \I__3372\ : InMux
    port map (
            O => \N__14879\,
            I => \N__14868\
        );

    \I__3371\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14861\
        );

    \I__3370\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14861\
        );

    \I__3369\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14861\
        );

    \I__3368\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14858\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__14868\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__14861\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14858\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__3364\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14843\
        );

    \I__3363\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14836\
        );

    \I__3362\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14836\
        );

    \I__3361\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14836\
        );

    \I__3360\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14832\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__14846\,
            I => \N__14829\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__14843\,
            I => \N__14822\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__14836\,
            I => \N__14822\
        );

    \I__3356\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14819\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__14832\,
            I => \N__14816\
        );

    \I__3354\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14811\
        );

    \I__3353\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14811\
        );

    \I__3352\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14808\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__14822\,
            I => \N__14805\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__14819\,
            I => \N__14800\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__14816\,
            I => \N__14800\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__14811\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__14808\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__14805\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__14800\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__3344\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14777\
        );

    \I__3343\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14777\
        );

    \I__3342\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14770\
        );

    \I__3341\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14770\
        );

    \I__3340\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14770\
        );

    \I__3339\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14766\
        );

    \I__3338\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14757\
        );

    \I__3337\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14757\
        );

    \I__3336\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14757\
        );

    \I__3335\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14757\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__14777\,
            I => \N__14754\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__14770\,
            I => \N__14751\
        );

    \I__3332\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14748\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__14766\,
            I => \N__14742\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__14757\,
            I => \N__14742\
        );

    \I__3329\ : Span4Mux_h
    port map (
            O => \N__14754\,
            I => \N__14735\
        );

    \I__3328\ : Span4Mux_s3_h
    port map (
            O => \N__14751\,
            I => \N__14735\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__14748\,
            I => \N__14735\
        );

    \I__3326\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14732\
        );

    \I__3325\ : Span4Mux_s2_h
    port map (
            O => \N__14742\,
            I => \N__14729\
        );

    \I__3324\ : Sp12to4
    port map (
            O => \N__14735\,
            I => \N__14724\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__14732\,
            I => \N__14724\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__14729\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__3321\ : Odrv12
    port map (
            O => \N__14724\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__3320\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14712\
        );

    \I__3319\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14709\
        );

    \I__3318\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14706\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__14716\,
            I => \N__14699\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__14715\,
            I => \N__14696\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__14712\,
            I => \N__14693\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14690\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N__14687\
        );

    \I__3312\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14682\
        );

    \I__3311\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14682\
        );

    \I__3310\ : InMux
    port map (
            O => \N__14703\,
            I => \N__14677\
        );

    \I__3309\ : InMux
    port map (
            O => \N__14702\,
            I => \N__14677\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14672\
        );

    \I__3307\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14672\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__14693\,
            I => \N__14659\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__14690\,
            I => \N__14659\
        );

    \I__3304\ : Span4Mux_v
    port map (
            O => \N__14687\,
            I => \N__14659\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__14682\,
            I => \N__14659\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14659\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__14672\,
            I => \N__14659\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__14656\,
            I => \beamY_RNIFC5HAZ0Z_4\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__14653\,
            I => \N__14647\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__14652\,
            I => \N__14643\
        );

    \I__3296\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14633\
        );

    \I__3295\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14633\
        );

    \I__3294\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14633\
        );

    \I__3293\ : InMux
    port map (
            O => \N__14646\,
            I => \N__14633\
        );

    \I__3292\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14628\
        );

    \I__3291\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14628\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__14633\,
            I => \N__14625\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__14628\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__14625\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14614\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__14614\,
            I => chary_if_generate_plus_mult1_un47_sum_ac0_8
        );

    \I__3284\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14601\
        );

    \I__3283\ : InMux
    port map (
            O => \N__14610\,
            I => \N__14601\
        );

    \I__3282\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14596\
        );

    \I__3281\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14596\
        );

    \I__3280\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14591\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14591\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__14601\,
            I => \counter_RNI4HQB1Z0Z_5\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__14596\,
            I => \counter_RNI4HQB1Z0Z_5\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__14591\,
            I => \counter_RNI4HQB1Z0Z_5\
        );

    \I__3275\ : InMux
    port map (
            O => \N__14584\,
            I => counter_cry_4
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__14581\,
            I => \N__14578\
        );

    \I__3273\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14574\
        );

    \I__3272\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14566\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__14574\,
            I => \N__14563\
        );

    \I__3270\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14556\
        );

    \I__3269\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14556\
        );

    \I__3268\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14556\
        );

    \I__3267\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14551\
        );

    \I__3266\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14551\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__14566\,
            I => \counterZ0Z_5\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__14563\,
            I => \counterZ0Z_5\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__14556\,
            I => \counterZ0Z_5\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__14551\,
            I => \counterZ0Z_5\
        );

    \I__3261\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14527\
        );

    \I__3260\ : InMux
    port map (
            O => \N__14541\,
            I => \N__14522\
        );

    \I__3259\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14522\
        );

    \I__3258\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14518\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14515\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14508\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14508\
        );

    \I__3254\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14508\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14505\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14500\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14500\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14495\
        );

    \I__3249\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14495\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__14527\,
            I => \N__14490\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14490\
        );

    \I__3246\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14487\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14482\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14515\,
            I => \N__14482\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__14508\,
            I => \N__14479\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14474\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__14500\,
            I => \N__14474\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14495\,
            I => \N__14471\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__14490\,
            I => \N__14466\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__14487\,
            I => \N__14466\
        );

    \I__3237\ : Span12Mux_s9_h
    port map (
            O => \N__14482\,
            I => \N__14463\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__14479\,
            I => \N__14460\
        );

    \I__3235\ : Span4Mux_v
    port map (
            O => \N__14474\,
            I => \N__14455\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__14471\,
            I => \N__14455\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__14466\,
            I => \N__14452\
        );

    \I__3232\ : Odrv12
    port map (
            O => \N__14463\,
            I => \SDATA1_c\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__14460\,
            I => \SDATA1_c\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__14455\,
            I => \SDATA1_c\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__14452\,
            I => \SDATA1_c\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__3227\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14430\
        );

    \I__3226\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14427\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14424\
        );

    \I__3224\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14421\
        );

    \I__3223\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14418\
        );

    \I__3222\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14411\
        );

    \I__3221\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14411\
        );

    \I__3220\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14411\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__14430\,
            I => \N__14408\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__14427\,
            I => \slaveselectZ0\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__14424\,
            I => \slaveselectZ0\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__14421\,
            I => \slaveselectZ0\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__14418\,
            I => \slaveselectZ0\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__14411\,
            I => \slaveselectZ0\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__14408\,
            I => \slaveselectZ0\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__14395\,
            I => \N__14391\
        );

    \I__3211\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14387\
        );

    \I__3210\ : InMux
    port map (
            O => \N__14391\,
            I => \N__14384\
        );

    \I__3209\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14381\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__14387\,
            I => un5_slaveselect
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__14384\,
            I => un5_slaveselect
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14381\,
            I => un5_slaveselect
        );

    \I__3205\ : IoInMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14367\
        );

    \I__3203\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14364\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__14367\,
            I => \SDATA2_c\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__14364\,
            I => \SDATA2_c\
        );

    \I__3200\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14355\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14352\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14355\,
            I => \N__14348\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__14352\,
            I => \N__14336\
        );

    \I__3196\ : ClkMux
    port map (
            O => \N__14351\,
            I => \N__14311\
        );

    \I__3195\ : Glb2LocalMux
    port map (
            O => \N__14348\,
            I => \N__14311\
        );

    \I__3194\ : ClkMux
    port map (
            O => \N__14347\,
            I => \N__14311\
        );

    \I__3193\ : ClkMux
    port map (
            O => \N__14346\,
            I => \N__14311\
        );

    \I__3192\ : ClkMux
    port map (
            O => \N__14345\,
            I => \N__14311\
        );

    \I__3191\ : ClkMux
    port map (
            O => \N__14344\,
            I => \N__14311\
        );

    \I__3190\ : ClkMux
    port map (
            O => \N__14343\,
            I => \N__14311\
        );

    \I__3189\ : ClkMux
    port map (
            O => \N__14342\,
            I => \N__14311\
        );

    \I__3188\ : ClkMux
    port map (
            O => \N__14341\,
            I => \N__14311\
        );

    \I__3187\ : ClkMux
    port map (
            O => \N__14340\,
            I => \N__14311\
        );

    \I__3186\ : ClkMux
    port map (
            O => \N__14339\,
            I => \N__14311\
        );

    \I__3185\ : Glb2LocalMux
    port map (
            O => \N__14336\,
            I => \N__14311\
        );

    \I__3184\ : GlobalMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__3183\ : gio2CtrlBuf
    port map (
            O => \N__14308\,
            I => \Clock12MHz_c_g\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__14305\,
            I => \chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_\
        );

    \I__3181\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14299\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__14299\,
            I => \N__14296\
        );

    \I__3179\ : Span4Mux_v
    port map (
            O => \N__14296\,
            I => \N__14293\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__14293\,
            I => \beamY_RNII78UPZ0Z_4\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__14290\,
            I => \chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__14287\,
            I => \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_\
        );

    \I__3175\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14269\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14269\
        );

    \I__3173\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14260\
        );

    \I__3172\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14260\
        );

    \I__3171\ : InMux
    port map (
            O => \N__14280\,
            I => \N__14257\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14252\
        );

    \I__3169\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14252\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14245\
        );

    \I__3167\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14245\
        );

    \I__3166\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14245\
        );

    \I__3165\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14242\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__14269\,
            I => \N__14239\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14230\
        );

    \I__3162\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14230\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14230\
        );

    \I__3160\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14230\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__14260\,
            I => \N__14225\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__14257\,
            I => \N__14225\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__14252\,
            I => \N__14220\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__14245\,
            I => \N__14220\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14213\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__14239\,
            I => \N__14213\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__14230\,
            I => \N__14213\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__14225\,
            I => \N__14210\
        );

    \I__3151\ : Odrv12
    port map (
            O => \N__14220\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__14213\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__14210\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__3148\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14197\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__14197\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\
        );

    \I__3144\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14188\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__14188\,
            I => \N__14185\
        );

    \I__3142\ : Span4Mux_s3_v
    port map (
            O => \N__14185\,
            I => \N__14181\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14178\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__14181\,
            I => un1_counter_0_1
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__14178\,
            I => un1_counter_0_1
        );

    \I__3138\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14167\
        );

    \I__3137\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14164\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14161\
        );

    \I__3135\ : InMux
    port map (
            O => \N__14170\,
            I => \N__14158\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14167\,
            I => un7_slaveselectlt5
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__14164\,
            I => un7_slaveselectlt5
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__14161\,
            I => un7_slaveselectlt5
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14158\,
            I => un7_slaveselectlt5
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__14149\,
            I => \un1_counter_0_1_cascade_\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__14146\,
            I => \slaveselect_1lto5_0_cascade_\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14142\,
            I => \N__14137\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__14137\,
            I => slaveselect_1lto5_1
        );

    \I__3125\ : IoInMux
    port map (
            O => \N__14134\,
            I => \N__14130\
        );

    \I__3124\ : IoInMux
    port map (
            O => \N__14133\,
            I => \N__14127\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__14130\,
            I => \N__14122\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__14127\,
            I => \N__14122\
        );

    \I__3121\ : Span4Mux_s3_v
    port map (
            O => \N__14122\,
            I => \N__14119\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__14119\,
            I => \SCLK1_0_i\
        );

    \I__3119\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14102\
        );

    \I__3118\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14099\
        );

    \I__3117\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14094\
        );

    \I__3116\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14094\
        );

    \I__3115\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14089\
        );

    \I__3114\ : InMux
    port map (
            O => \N__14111\,
            I => \N__14089\
        );

    \I__3113\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14084\
        );

    \I__3112\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14084\
        );

    \I__3111\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14081\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14074\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14074\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14074\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__14102\,
            I => \counterZ0Z_1\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__14099\,
            I => \counterZ0Z_1\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__14094\,
            I => \counterZ0Z_1\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14089\,
            I => \counterZ0Z_1\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__14084\,
            I => \counterZ0Z_1\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__14081\,
            I => \counterZ0Z_1\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14074\,
            I => \counterZ0Z_1\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__14059\,
            I => \N__14050\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__14058\,
            I => \N__14039\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__14057\,
            I => \N__14036\
        );

    \I__3097\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14032\
        );

    \I__3096\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14025\
        );

    \I__3095\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14025\
        );

    \I__3094\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14025\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14022\
        );

    \I__3092\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14017\
        );

    \I__3091\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14017\
        );

    \I__3090\ : InMux
    port map (
            O => \N__14047\,
            I => \N__14010\
        );

    \I__3089\ : InMux
    port map (
            O => \N__14046\,
            I => \N__14010\
        );

    \I__3088\ : InMux
    port map (
            O => \N__14045\,
            I => \N__14010\
        );

    \I__3087\ : InMux
    port map (
            O => \N__14044\,
            I => \N__14003\
        );

    \I__3086\ : InMux
    port map (
            O => \N__14043\,
            I => \N__14003\
        );

    \I__3085\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14003\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14000\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14036\,
            I => \N__13995\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14035\,
            I => \N__13995\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__14032\,
            I => \counterZ0Z_0\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__14025\,
            I => \counterZ0Z_0\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14022\,
            I => \counterZ0Z_0\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__14017\,
            I => \counterZ0Z_0\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__14010\,
            I => \counterZ0Z_0\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__14003\,
            I => \counterZ0Z_0\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__14000\,
            I => \counterZ0Z_0\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__13995\,
            I => \counterZ0Z_0\
        );

    \I__3073\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13975\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__13975\,
            I => \N__13970\
        );

    \I__3071\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13965\
        );

    \I__3070\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13965\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__13970\,
            I => un7_slaveselectlt2_0
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__13965\,
            I => un7_slaveselectlt2_0
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \N__13957\
        );

    \I__3066\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13945\
        );

    \I__3064\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13940\
        );

    \I__3063\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13940\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13937\
        );

    \I__3061\ : InMux
    port map (
            O => \N__13950\,
            I => \N__13930\
        );

    \I__3060\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13930\
        );

    \I__3059\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13930\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__13945\,
            I => \counterZ0Z_2\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13940\,
            I => \counterZ0Z_2\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__13937\,
            I => \counterZ0Z_2\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__13930\,
            I => \counterZ0Z_2\
        );

    \I__3054\ : InMux
    port map (
            O => \N__13921\,
            I => counter_cry_1
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__13918\,
            I => \N__13912\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__13917\,
            I => \N__13909\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__13916\,
            I => \N__13905\
        );

    \I__3050\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13900\
        );

    \I__3049\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13897\
        );

    \I__3048\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13894\
        );

    \I__3047\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13889\
        );

    \I__3046\ : InMux
    port map (
            O => \N__13905\,
            I => \N__13889\
        );

    \I__3045\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13885\
        );

    \I__3044\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13882\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__13900\,
            I => \N__13877\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13877\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__13894\,
            I => \N__13874\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__13889\,
            I => \N__13871\
        );

    \I__3039\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13868\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__13885\,
            I => \counterZ0Z_3\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__13882\,
            I => \counterZ0Z_3\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__13877\,
            I => \counterZ0Z_3\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__13874\,
            I => \counterZ0Z_3\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__13871\,
            I => \counterZ0Z_3\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__13868\,
            I => \counterZ0Z_3\
        );

    \I__3032\ : InMux
    port map (
            O => \N__13855\,
            I => counter_cry_2
        );

    \I__3031\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13846\
        );

    \I__3030\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13843\
        );

    \I__3029\ : InMux
    port map (
            O => \N__13850\,
            I => \N__13838\
        );

    \I__3028\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13838\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__13846\,
            I => \counterZ0Z_4\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13843\,
            I => \counterZ0Z_4\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__13838\,
            I => \counterZ0Z_4\
        );

    \I__3024\ : InMux
    port map (
            O => \N__13831\,
            I => counter_cry_3
        );

    \I__3023\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__3022\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13822\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__13822\,
            I => content_ram10_0
        );

    \I__3020\ : CEMux
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__13816\,
            I => \N__13813\
        );

    \I__3018\ : Odrv12
    port map (
            O => \N__13813\,
            I => content_awe10
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \content_N_35_cascade_\
        );

    \I__3016\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13804\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__13804\,
            I => content_awe3_1
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__13801\,
            I => \content_awe3_1_cascade_\
        );

    \I__3013\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13793\
        );

    \I__3012\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13788\
        );

    \I__3011\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13788\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__13793\,
            I => content_ram2_0
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__13788\,
            I => content_ram2_0
        );

    \I__3008\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13778\
        );

    \I__3007\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13775\
        );

    \I__3006\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13772\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__13778\,
            I => \content_N_40\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__13775\,
            I => \content_N_40\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__13772\,
            I => \content_N_40\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__13764\,
            I => \N__13754\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__13763\,
            I => \N__13751\
        );

    \I__2999\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13748\
        );

    \I__2998\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13745\
        );

    \I__2997\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13736\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13736\
        );

    \I__2995\ : InMux
    port map (
            O => \N__13754\,
            I => \N__13736\
        );

    \I__2994\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13736\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__13748\,
            I => \content_N_35\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__13745\,
            I => \content_N_35\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__13736\,
            I => \content_N_35\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \content_awe1_0_a2_0_cascade_\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__13726\,
            I => \N__13722\
        );

    \I__2988\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13717\
        );

    \I__2987\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13717\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13713\
        );

    \I__2985\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13710\
        );

    \I__2984\ : Span4Mux_h
    port map (
            O => \N__13713\,
            I => \N__13707\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13710\,
            I => content_ram1_0
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__13707\,
            I => content_ram1_0
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__13702\,
            I => \un7_slaveselectlt5_cascade_\
        );

    \I__2980\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13692\
        );

    \I__2979\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13687\
        );

    \I__2978\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13687\
        );

    \I__2977\ : InMux
    port map (
            O => \N__13696\,
            I => \N__13682\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13682\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__13692\,
            I => \N_190_i\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N_190_i\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N_190_i\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__13675\,
            I => \N__13672\
        );

    \I__2971\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13669\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__13669\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\
        );

    \I__2969\ : InMux
    port map (
            O => \N__13666\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__13663\,
            I => \N__13660\
        );

    \I__2967\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13657\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__13657\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__13654\,
            I => \N__13651\
        );

    \I__2964\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13648\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__13648\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\
        );

    \I__2962\ : InMux
    port map (
            O => \N__13645\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2961\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13639\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__13639\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__13636\,
            I => \N__13632\
        );

    \I__2958\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13627\
        );

    \I__2957\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13627\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__13627\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02\
        );

    \I__2955\ : InMux
    port map (
            O => \N__13624\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__13621\,
            I => \N__13618\
        );

    \I__2953\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13615\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__13615\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81\
        );

    \I__2951\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13609\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__13609\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__2949\ : InMux
    port map (
            O => \N__13606\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__2948\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13600\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__13600\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__2946\ : InMux
    port map (
            O => \N__13597\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__2945\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13587\
        );

    \I__2944\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13584\
        );

    \I__2943\ : InMux
    port map (
            O => \N__13592\,
            I => \N__13577\
        );

    \I__2942\ : InMux
    port map (
            O => \N__13591\,
            I => \N__13577\
        );

    \I__2941\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13577\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__13587\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__13584\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__13577\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__13570\,
            I => \N__13565\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__13569\,
            I => \N__13561\
        );

    \I__2935\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13557\
        );

    \I__2934\ : InMux
    port map (
            O => \N__13565\,
            I => \N__13548\
        );

    \I__2933\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13548\
        );

    \I__2932\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13548\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13548\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__13557\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__13548\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\
        );

    \I__2928\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13540\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__13540\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__2926\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13534\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__13534\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__2924\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13526\
        );

    \I__2923\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13521\
        );

    \I__2922\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13521\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13515\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__13521\,
            I => \N__13512\
        );

    \I__2919\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13509\
        );

    \I__2918\ : InMux
    port map (
            O => \N__13519\,
            I => \N__13506\
        );

    \I__2917\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13503\
        );

    \I__2916\ : Span4Mux_h
    port map (
            O => \N__13515\,
            I => \N__13500\
        );

    \I__2915\ : Odrv4
    port map (
            O => \N__13512\,
            I => \beamY_RNI9DLCZ0Z_1\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__13509\,
            I => \beamY_RNI9DLCZ0Z_1\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13506\,
            I => \beamY_RNI9DLCZ0Z_1\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__13503\,
            I => \beamY_RNI9DLCZ0Z_1\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__13500\,
            I => \beamY_RNI9DLCZ0Z_1\
        );

    \I__2910\ : InMux
    port map (
            O => \N__13489\,
            I => \bfn_9_8_0_\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13482\
        );

    \I__2908\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13477\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13474\
        );

    \I__2906\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13469\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13480\,
            I => \N__13469\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13477\,
            I => \N__13459\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__13474\,
            I => \N__13459\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13459\
        );

    \I__2901\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13456\
        );

    \I__2900\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13453\
        );

    \I__2899\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13448\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__13459\,
            I => \N__13445\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__13456\,
            I => \N__13440\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__13453\,
            I => \N__13440\
        );

    \I__2895\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13435\
        );

    \I__2894\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13435\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__13448\,
            I => \beamYZ0Z_9\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__13445\,
            I => \beamYZ0Z_9\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__13440\,
            I => \beamYZ0Z_9\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__13435\,
            I => \beamYZ0Z_9\
        );

    \I__2889\ : ClkMux
    port map (
            O => \N__13426\,
            I => \N__13399\
        );

    \I__2888\ : ClkMux
    port map (
            O => \N__13425\,
            I => \N__13399\
        );

    \I__2887\ : ClkMux
    port map (
            O => \N__13424\,
            I => \N__13399\
        );

    \I__2886\ : ClkMux
    port map (
            O => \N__13423\,
            I => \N__13399\
        );

    \I__2885\ : ClkMux
    port map (
            O => \N__13422\,
            I => \N__13399\
        );

    \I__2884\ : ClkMux
    port map (
            O => \N__13421\,
            I => \N__13399\
        );

    \I__2883\ : ClkMux
    port map (
            O => \N__13420\,
            I => \N__13399\
        );

    \I__2882\ : ClkMux
    port map (
            O => \N__13419\,
            I => \N__13399\
        );

    \I__2881\ : ClkMux
    port map (
            O => \N__13418\,
            I => \N__13399\
        );

    \I__2880\ : GlobalMux
    port map (
            O => \N__13399\,
            I => \N__13396\
        );

    \I__2879\ : gio2CtrlBuf
    port map (
            O => \N__13396\,
            I => \PixelClock_g\
        );

    \I__2878\ : CEMux
    port map (
            O => \N__13393\,
            I => \N__13388\
        );

    \I__2877\ : CEMux
    port map (
            O => \N__13392\,
            I => \N__13385\
        );

    \I__2876\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13381\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__13388\,
            I => \N__13378\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__13385\,
            I => \N__13375\
        );

    \I__2873\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13370\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__13381\,
            I => \N__13367\
        );

    \I__2871\ : Span4Mux_v
    port map (
            O => \N__13378\,
            I => \N__13364\
        );

    \I__2870\ : Span4Mux_v
    port map (
            O => \N__13375\,
            I => \N__13361\
        );

    \I__2869\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13355\
        );

    \I__2868\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13355\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N__13352\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__13367\,
            I => \N__13345\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__13364\,
            I => \N__13345\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__13361\,
            I => \N__13345\
        );

    \I__2863\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13342\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13339\
        );

    \I__2861\ : Span12Mux_s8_v
    port map (
            O => \N__13352\,
            I => \N__13336\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__13345\,
            I => \N__13333\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__13342\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__13339\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__2857\ : Odrv12
    port map (
            O => \N__13336\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__13333\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__2855\ : InMux
    port map (
            O => \N__13324\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__2854\ : InMux
    port map (
            O => \N__13321\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__2853\ : InMux
    port map (
            O => \N__13318\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__2852\ : InMux
    port map (
            O => \N__13315\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__2851\ : InMux
    port map (
            O => \N__13312\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__2850\ : InMux
    port map (
            O => \N__13309\,
            I => \N__13306\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__13306\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__2848\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__13300\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__2846\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13291\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__13296\,
            I => \N__13284\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__13295\,
            I => \N__13280\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__13294\,
            I => \N__13277\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__13291\,
            I => \N__13273\
        );

    \I__2841\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13268\
        );

    \I__2840\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13268\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__13288\,
            I => \N__13259\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13253\
        );

    \I__2837\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13248\
        );

    \I__2836\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13243\
        );

    \I__2835\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13243\
        );

    \I__2834\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13240\
        );

    \I__2833\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13237\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__13273\,
            I => \N__13232\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__13268\,
            I => \N__13232\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13227\
        );

    \I__2829\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13227\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13223\
        );

    \I__2827\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13220\
        );

    \I__2826\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13213\
        );

    \I__2825\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13213\
        );

    \I__2824\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13213\
        );

    \I__2823\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13210\
        );

    \I__2822\ : InMux
    port map (
            O => \N__13257\,
            I => \N__13205\
        );

    \I__2821\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13205\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13202\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13198\
        );

    \I__2818\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13194\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__13248\,
            I => \N__13187\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13187\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__13240\,
            I => \N__13187\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__13237\,
            I => \N__13180\
        );

    \I__2813\ : Span4Mux_s2_v
    port map (
            O => \N__13232\,
            I => \N__13180\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__13227\,
            I => \N__13180\
        );

    \I__2811\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13175\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13175\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13166\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__13213\,
            I => \N__13166\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__13210\,
            I => \N__13166\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__13205\,
            I => \N__13166\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__13202\,
            I => \N__13163\
        );

    \I__2804\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13160\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__13198\,
            I => \N__13157\
        );

    \I__2802\ : InMux
    port map (
            O => \N__13197\,
            I => \N__13152\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__13194\,
            I => \N__13147\
        );

    \I__2800\ : Span12Mux_s6_h
    port map (
            O => \N__13187\,
            I => \N__13147\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__13180\,
            I => \N__13140\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13140\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__13166\,
            I => \N__13140\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__13163\,
            I => \N__13135\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__13160\,
            I => \N__13135\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__13157\,
            I => \N__13132\
        );

    \I__2793\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13127\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13127\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13152\,
            I => \beamYZ0Z_1\
        );

    \I__2790\ : Odrv12
    port map (
            O => \N__13147\,
            I => \beamYZ0Z_1\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__13140\,
            I => \beamYZ0Z_1\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__13135\,
            I => \beamYZ0Z_1\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__13132\,
            I => \beamYZ0Z_1\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__13127\,
            I => \beamYZ0Z_1\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \N__13110\
        );

    \I__2784\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13102\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13094\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13094\
        );

    \I__2781\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13086\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13083\
        );

    \I__2779\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13080\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__13105\,
            I => \N__13077\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__13102\,
            I => \N__13071\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13068\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13063\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13063\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13060\
        );

    \I__2772\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13057\
        );

    \I__2771\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13052\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13045\
        );

    \I__2769\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13045\
        );

    \I__2768\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13045\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__13086\,
            I => \N__13038\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__13083\,
            I => \N__13038\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13080\,
            I => \N__13038\
        );

    \I__2764\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13033\
        );

    \I__2763\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13033\
        );

    \I__2762\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13030\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \N__13027\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__13071\,
            I => \N__13023\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__13068\,
            I => \N__13020\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__13063\,
            I => \N__13017\
        );

    \I__2757\ : Span4Mux_h
    port map (
            O => \N__13060\,
            I => \N__13014\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__13057\,
            I => \N__13011\
        );

    \I__2755\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13006\
        );

    \I__2754\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13006\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13003\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__13045\,
            I => \N__12998\
        );

    \I__2751\ : Span4Mux_s3_v
    port map (
            O => \N__13038\,
            I => \N__12998\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__13033\,
            I => \N__12993\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__13030\,
            I => \N__12993\
        );

    \I__2748\ : InMux
    port map (
            O => \N__13027\,
            I => \N__12990\
        );

    \I__2747\ : InMux
    port map (
            O => \N__13026\,
            I => \N__12987\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__13023\,
            I => \N__12982\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__13020\,
            I => \N__12982\
        );

    \I__2744\ : Span4Mux_v
    port map (
            O => \N__13017\,
            I => \N__12975\
        );

    \I__2743\ : Span4Mux_v
    port map (
            O => \N__13014\,
            I => \N__12975\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__13011\,
            I => \N__12975\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__13006\,
            I => \N__12968\
        );

    \I__2740\ : Span4Mux_s3_v
    port map (
            O => \N__13003\,
            I => \N__12968\
        );

    \I__2739\ : Span4Mux_h
    port map (
            O => \N__12998\,
            I => \N__12968\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__12993\,
            I => \N__12965\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__12990\,
            I => \beamYZ0Z_0\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__12987\,
            I => \beamYZ0Z_0\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__12982\,
            I => \beamYZ0Z_0\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__12975\,
            I => \beamYZ0Z_0\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__12968\,
            I => \beamYZ0Z_0\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__12965\,
            I => \beamYZ0Z_0\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__12952\,
            I => \N__12949\
        );

    \I__2730\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12946\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12943\
        );

    \I__2728\ : Span4Mux_h
    port map (
            O => \N__12943\,
            I => \N__12940\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__12940\,
            I => \N__12937\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__12937\,
            I => g2_1_1_0
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__12934\,
            I => \N__12927\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__12933\,
            I => \N__12923\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__12932\,
            I => \N__12914\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__12931\,
            I => \N__12907\
        );

    \I__2721\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12904\
        );

    \I__2720\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12901\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12892\
        );

    \I__2718\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12892\
        );

    \I__2717\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12892\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12892\
        );

    \I__2715\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12889\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__12919\,
            I => \N__12883\
        );

    \I__2713\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12872\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12867\
        );

    \I__2711\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12867\
        );

    \I__2710\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12862\
        );

    \I__2709\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12862\
        );

    \I__2708\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12853\
        );

    \I__2707\ : InMux
    port map (
            O => \N__12910\,
            I => \N__12848\
        );

    \I__2706\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12848\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__12904\,
            I => \N__12839\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__12901\,
            I => \N__12839\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__12892\,
            I => \N__12839\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12839\
        );

    \I__2701\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12835\
        );

    \I__2700\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12830\
        );

    \I__2699\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12830\
        );

    \I__2698\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12825\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12825\
        );

    \I__2696\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12822\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12815\
        );

    \I__2694\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12815\
        );

    \I__2693\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12815\
        );

    \I__2692\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12808\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12808\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12808\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__12872\,
            I => \N__12799\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__12867\,
            I => \N__12799\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__12862\,
            I => \N__12796\
        );

    \I__2686\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12789\
        );

    \I__2685\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12789\
        );

    \I__2684\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12789\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12786\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12783\
        );

    \I__2681\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12780\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__12853\,
            I => \N__12775\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12775\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__12839\,
            I => \N__12772\
        );

    \I__2677\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12769\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__12835\,
            I => \N__12756\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__12830\,
            I => \N__12756\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12825\,
            I => \N__12756\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__12822\,
            I => \N__12756\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__12815\,
            I => \N__12756\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__12808\,
            I => \N__12756\
        );

    \I__2670\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12751\
        );

    \I__2669\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12751\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__12805\,
            I => \N__12747\
        );

    \I__2667\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12739\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__12799\,
            I => \N__12736\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__12796\,
            I => \N__12725\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__12789\,
            I => \N__12725\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__12786\,
            I => \N__12725\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__12783\,
            I => \N__12725\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__12780\,
            I => \N__12725\
        );

    \I__2660\ : Span12Mux_s6_v
    port map (
            O => \N__12775\,
            I => \N__12718\
        );

    \I__2659\ : Sp12to4
    port map (
            O => \N__12772\,
            I => \N__12718\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12718\
        );

    \I__2657\ : Span4Mux_v
    port map (
            O => \N__12756\,
            I => \N__12713\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__12751\,
            I => \N__12713\
        );

    \I__2655\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12710\
        );

    \I__2654\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12707\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12700\
        );

    \I__2652\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12700\
        );

    \I__2651\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12700\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12695\
        );

    \I__2649\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12695\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__12739\,
            I => \beamYZ0Z_2\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__12736\,
            I => \beamYZ0Z_2\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__12725\,
            I => \beamYZ0Z_2\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__12718\,
            I => \beamYZ0Z_2\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__12713\,
            I => \beamYZ0Z_2\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__12710\,
            I => \beamYZ0Z_2\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__12707\,
            I => \beamYZ0Z_2\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__12700\,
            I => \beamYZ0Z_2\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__12695\,
            I => \beamYZ0Z_2\
        );

    \I__2639\ : InMux
    port map (
            O => \N__12676\,
            I => un21_beamy_cry_1
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__12673\,
            I => \N__12666\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__12672\,
            I => \N__12661\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \N__12657\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__12670\,
            I => \N__12645\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__12669\,
            I => \N__12639\
        );

    \I__2633\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12631\
        );

    \I__2632\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12631\
        );

    \I__2631\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12628\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12625\
        );

    \I__2629\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12622\
        );

    \I__2628\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12617\
        );

    \I__2627\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12617\
        );

    \I__2626\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12608\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12608\
        );

    \I__2624\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12608\
        );

    \I__2623\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12608\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12601\
        );

    \I__2621\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12601\
        );

    \I__2620\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12601\
        );

    \I__2619\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12596\
        );

    \I__2618\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12589\
        );

    \I__2617\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12589\
        );

    \I__2616\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12589\
        );

    \I__2615\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12582\
        );

    \I__2614\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12575\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12575\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12575\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12572\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__12631\,
            I => \N__12563\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__12628\,
            I => \N__12563\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__12625\,
            I => \N__12563\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12622\,
            I => \N__12563\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__12617\,
            I => \N__12556\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__12608\,
            I => \N__12556\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12556\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12553\
        );

    \I__2602\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12550\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12596\,
            I => \N__12545\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__12589\,
            I => \N__12545\
        );

    \I__2599\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12542\
        );

    \I__2598\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12539\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__12586\,
            I => \N__12535\
        );

    \I__2596\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12526\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__12582\,
            I => \N__12523\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__12575\,
            I => \N__12516\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12516\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__12563\,
            I => \N__12516\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__12556\,
            I => \N__12513\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__12553\,
            I => \N__12508\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__12550\,
            I => \N__12508\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__12545\,
            I => \N__12501\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__12542\,
            I => \N__12501\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__12539\,
            I => \N__12501\
        );

    \I__2585\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12496\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12496\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12489\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12489\
        );

    \I__2581\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12489\
        );

    \I__2580\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12482\
        );

    \I__2579\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12482\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12482\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12526\,
            I => \beamYZ0Z_3\
        );

    \I__2576\ : Odrv12
    port map (
            O => \N__12523\,
            I => \beamYZ0Z_3\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__12516\,
            I => \beamYZ0Z_3\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__12513\,
            I => \beamYZ0Z_3\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__12508\,
            I => \beamYZ0Z_3\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__12501\,
            I => \beamYZ0Z_3\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__12496\,
            I => \beamYZ0Z_3\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__12489\,
            I => \beamYZ0Z_3\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12482\,
            I => \beamYZ0Z_3\
        );

    \I__2568\ : InMux
    port map (
            O => \N__12463\,
            I => un21_beamy_cry_2
        );

    \I__2567\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12452\
        );

    \I__2566\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12447\
        );

    \I__2565\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12447\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12442\
        );

    \I__2563\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12442\
        );

    \I__2562\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12429\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__12452\,
            I => \N__12424\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__12447\,
            I => \N__12424\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12421\
        );

    \I__2558\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12418\
        );

    \I__2557\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12413\
        );

    \I__2556\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12413\
        );

    \I__2555\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12410\
        );

    \I__2554\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12407\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__12436\,
            I => \N__12402\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__12435\,
            I => \N__12399\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__12434\,
            I => \N__12395\
        );

    \I__2550\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12391\
        );

    \I__2549\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12388\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__12429\,
            I => \N__12385\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__12424\,
            I => \N__12382\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__12421\,
            I => \N__12377\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__12418\,
            I => \N__12377\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12370\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12410\,
            I => \N__12370\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12370\
        );

    \I__2541\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12367\
        );

    \I__2540\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12364\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12357\
        );

    \I__2538\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12357\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12357\
        );

    \I__2536\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12352\
        );

    \I__2535\ : InMux
    port map (
            O => \N__12394\,
            I => \N__12352\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__12391\,
            I => \beamYZ0Z_4\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__12388\,
            I => \beamYZ0Z_4\
        );

    \I__2532\ : Odrv12
    port map (
            O => \N__12385\,
            I => \beamYZ0Z_4\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__12382\,
            I => \beamYZ0Z_4\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__12377\,
            I => \beamYZ0Z_4\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__12370\,
            I => \beamYZ0Z_4\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__12367\,
            I => \beamYZ0Z_4\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__12364\,
            I => \beamYZ0Z_4\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12357\,
            I => \beamYZ0Z_4\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__12352\,
            I => \beamYZ0Z_4\
        );

    \I__2524\ : InMux
    port map (
            O => \N__12331\,
            I => un21_beamy_cry_3
        );

    \I__2523\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12325\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__12325\,
            I => \N__12318\
        );

    \I__2521\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12315\
        );

    \I__2520\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12310\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12310\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12299\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__12318\,
            I => \N__12296\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12293\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__12310\,
            I => \N__12290\
        );

    \I__2514\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12285\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12285\
        );

    \I__2512\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12280\
        );

    \I__2511\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12280\
        );

    \I__2510\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12271\
        );

    \I__2509\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12271\
        );

    \I__2508\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12271\
        );

    \I__2507\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12271\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__12299\,
            I => \beamYZ0Z_5\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__12296\,
            I => \beamYZ0Z_5\
        );

    \I__2504\ : Odrv12
    port map (
            O => \N__12293\,
            I => \beamYZ0Z_5\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__12290\,
            I => \beamYZ0Z_5\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__12285\,
            I => \beamYZ0Z_5\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__12280\,
            I => \beamYZ0Z_5\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__12271\,
            I => \beamYZ0Z_5\
        );

    \I__2499\ : InMux
    port map (
            O => \N__12256\,
            I => un21_beamy_cry_4
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__2497\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12247\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__12247\,
            I => \N__12244\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__12244\,
            I => \N__12237\
        );

    \I__2494\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12234\
        );

    \I__2493\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12229\
        );

    \I__2492\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12229\
        );

    \I__2491\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12219\
        );

    \I__2490\ : Span4Mux_s3_h
    port map (
            O => \N__12237\,
            I => \N__12216\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12213\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__12229\,
            I => \N__12210\
        );

    \I__2487\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12205\
        );

    \I__2486\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12205\
        );

    \I__2485\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12202\
        );

    \I__2484\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12199\
        );

    \I__2483\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12192\
        );

    \I__2482\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12192\
        );

    \I__2481\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12192\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__12219\,
            I => \beamYZ0Z_6\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__12216\,
            I => \beamYZ0Z_6\
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__12213\,
            I => \beamYZ0Z_6\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__12210\,
            I => \beamYZ0Z_6\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__12205\,
            I => \beamYZ0Z_6\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__12202\,
            I => \beamYZ0Z_6\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__12199\,
            I => \beamYZ0Z_6\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__12192\,
            I => \beamYZ0Z_6\
        );

    \I__2472\ : InMux
    port map (
            O => \N__12175\,
            I => un21_beamy_cry_5
        );

    \I__2471\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12166\
        );

    \I__2470\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12166\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12157\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12154\
        );

    \I__2466\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12145\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__12160\,
            I => \N__12142\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__12157\,
            I => \N__12137\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__12154\,
            I => \N__12137\
        );

    \I__2462\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12132\
        );

    \I__2461\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12132\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12127\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12127\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12122\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12122\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__12145\,
            I => \beamYZ0Z_7\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__12142\,
            I => \beamYZ0Z_7\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__12137\,
            I => \beamYZ0Z_7\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__12132\,
            I => \beamYZ0Z_7\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__12127\,
            I => \beamYZ0Z_7\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__12122\,
            I => \beamYZ0Z_7\
        );

    \I__2450\ : InMux
    port map (
            O => \N__12109\,
            I => un21_beamy_cry_6
        );

    \I__2449\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12099\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__2447\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12094\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12089\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12086\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__12099\,
            I => \N__12081\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__12094\,
            I => \N__12081\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \N__12073\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12092\,
            I => \N__12070\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__12089\,
            I => \N__12067\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__12086\,
            I => \N__12064\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__12081\,
            I => \N__12061\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12058\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12051\
        );

    \I__2435\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12051\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12051\
        );

    \I__2433\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12046\
        );

    \I__2432\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12046\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__12070\,
            I => \beamYZ0Z_8\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__12067\,
            I => \beamYZ0Z_8\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__12064\,
            I => \beamYZ0Z_8\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__12061\,
            I => \beamYZ0Z_8\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__12058\,
            I => \beamYZ0Z_8\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12051\,
            I => \beamYZ0Z_8\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__12046\,
            I => \beamYZ0Z_8\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12031\,
            I => un21_beamy_cry_7
        );

    \I__2423\ : InMux
    port map (
            O => \N__12028\,
            I => \N__12025\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__12025\,
            I => un5_visibley_3_29
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__12022\,
            I => \g1_8_1_cascade_\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__12019\,
            I => \N__12015\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12011\
        );

    \I__2418\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12006\
        );

    \I__2417\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12006\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__12011\,
            I => \N__11999\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__12006\,
            I => \N__11996\
        );

    \I__2414\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11985\
        );

    \I__2413\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11985\
        );

    \I__2412\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11985\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11980\
        );

    \I__2410\ : Span4Mux_h
    port map (
            O => \N__11999\,
            I => \N__11977\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__11996\,
            I => \N__11974\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11967\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11967\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11967\
        );

    \I__2405\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11964\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11985\,
            I => \N__11961\
        );

    \I__2403\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11958\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11955\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__11980\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__11977\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__11974\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__11967\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__11964\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__11961\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__11958\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__11955\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2393\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11935\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__11935\,
            I => \N__11932\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__11932\,
            I => g1_3_0
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__11929\,
            I => \N__11926\
        );

    \I__2389\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11923\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__11923\,
            I => \N__11920\
        );

    \I__2387\ : Odrv12
    port map (
            O => \N__11920\,
            I => un5_visibley_1_0_28
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__11917\,
            I => \beamY_RNIJ0H2Z0Z_4_cascade_\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__11914\,
            I => \N__11911\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11908\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__11908\,
            I => un5_visibley_c5
        );

    \I__2382\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11902\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11902\,
            I => un5_visibley_c6_0_0_0
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__11899\,
            I => \un5_visibley_c6_0_0_0_cascade_\
        );

    \I__2379\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11892\
        );

    \I__2378\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11889\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__11892\,
            I => un5_visibley_c3
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__11889\,
            I => un5_visibley_c3
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__11884\,
            I => \un19_slaveselectlt5_0_cascade_\
        );

    \I__2374\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__2373\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11875\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__11875\,
            I => un19_slaveselectlt5_0
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__11872\,
            I => \counter_RNI4HQB1Z0Z_5_cascade_\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__11869\,
            I => \beamY_RNI4FVGVZ0Z_4_cascade_\
        );

    \I__2369\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11857\
        );

    \I__2368\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11857\
        );

    \I__2367\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11852\
        );

    \I__2366\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11852\
        );

    \I__2365\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11849\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__11857\,
            I => \N__11846\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__11852\,
            I => \N__11843\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11849\,
            I => \N__11840\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__11846\,
            I => \N__11837\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__11843\,
            I => \N__11834\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__11840\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__11837\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__11834\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2356\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__11824\,
            I => \N__11821\
        );

    \I__2354\ : Span4Mux_h
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__11818\,
            I => \N_596_2\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__11815\,
            I => \un5_visibley_4_28_cascade_\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__11812\,
            I => \N__11809\
        );

    \I__2350\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11805\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__11808\,
            I => \N__11802\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__2347\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__11799\,
            I => \N__11793\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__11796\,
            I => content_ram12_0
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__11793\,
            I => content_ram12_0
        );

    \I__2343\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__11785\,
            I => content_awe0_0_a2_0
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \content_awe0_0_a2_0_cascade_\
        );

    \I__2340\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11772\
        );

    \I__2338\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11769\
        );

    \I__2337\ : Span4Mux_h
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__11769\,
            I => content_ram4_0
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__11766\,
            I => content_ram4_0
        );

    \I__2334\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11752\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11752\
        );

    \I__2332\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11752\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__11752\,
            I => \content_N_36\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \content_N_36_cascade_\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__11746\,
            I => \content_awe7_1_cascade_\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11739\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11736\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__11739\,
            I => \N__11733\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__11736\,
            I => content_ram6_0
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__11733\,
            I => content_ram6_0
        );

    \I__2323\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11725\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__11725\,
            I => content_awe7_1
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__11722\,
            I => \N__11718\
        );

    \I__2320\ : InMux
    port map (
            O => \N__11721\,
            I => \N__11715\
        );

    \I__2319\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11712\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__11715\,
            I => \N__11709\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11704\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__11709\,
            I => \N__11704\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__11704\,
            I => content_ram7_0
        );

    \I__2314\ : SRMux
    port map (
            O => \N__11701\,
            I => \N__11698\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__11698\,
            I => \nCS1_0_sqmuxa\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__11692\,
            I => \N__11688\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11679\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11679\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__11684\,
            I => \N__11676\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__11679\,
            I => \N__11673\
        );

    \I__2305\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11670\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__11673\,
            I => \N__11665\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11665\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__11662\,
            I => \content_N_19\
        );

    \I__2300\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11654\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11647\
        );

    \I__2298\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11647\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__11654\,
            I => \N__11638\
        );

    \I__2296\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11633\
        );

    \I__2295\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11633\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__11647\,
            I => \N__11630\
        );

    \I__2293\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11623\
        );

    \I__2292\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11623\
        );

    \I__2291\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11623\
        );

    \I__2290\ : InMux
    port map (
            O => \N__11643\,
            I => \N__11620\
        );

    \I__2289\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11617\
        );

    \I__2288\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11614\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__11638\,
            I => content_column_1_i_2_2
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__11633\,
            I => content_column_1_i_2_2
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__11630\,
            I => content_column_1_i_2_2
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__11623\,
            I => content_column_1_i_2_2
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__11620\,
            I => content_column_1_i_2_2
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__11617\,
            I => content_column_1_i_2_2
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__11614\,
            I => content_column_1_i_2_2
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11594\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__11598\,
            I => \N__11591\
        );

    \I__2278\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11586\
        );

    \I__2277\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11581\
        );

    \I__2276\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11581\
        );

    \I__2275\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11576\
        );

    \I__2274\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11576\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__11586\,
            I => \N__11567\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__11581\,
            I => \N__11564\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__11576\,
            I => \N__11561\
        );

    \I__2270\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11552\
        );

    \I__2269\ : InMux
    port map (
            O => \N__11574\,
            I => \N__11552\
        );

    \I__2268\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11552\
        );

    \I__2267\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11552\
        );

    \I__2266\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11549\
        );

    \I__2265\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11546\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__11567\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__11564\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__11561\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__11552\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__11549\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__11546\,
            I => if_generate_plus_mult1_un61_sum_s_5
        );

    \I__2258\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__11530\,
            I => \content_content_ram10__e_0_RNIOLNMN1Z0Z_0\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__11527\,
            I => \N__11522\
        );

    \I__2255\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11517\
        );

    \I__2254\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11517\
        );

    \I__2253\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11514\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11511\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__11514\,
            I => content_ram3_0
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__11511\,
            I => content_ram3_0
        );

    \I__2249\ : CEMux
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__11503\,
            I => content_awe9
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__11500\,
            I => \N__11496\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11493\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11490\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__11493\,
            I => \N__11487\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__11490\,
            I => content_ram0_0
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__11487\,
            I => content_ram0_0
        );

    \I__2241\ : CEMux
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__2239\ : Span4Mux_h
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__11473\,
            I => content_awe8
        );

    \I__2237\ : CEMux
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__11464\,
            I => content_awe11
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__11461\,
            I => \N__11457\
        );

    \I__2233\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11454\
        );

    \I__2232\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11451\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__11454\,
            I => \N__11448\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11451\,
            I => content_ram5_0
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__11448\,
            I => content_ram5_0
        );

    \I__2228\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__11440\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__2226\ : InMux
    port map (
            O => \N__11437\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__2225\ : InMux
    port map (
            O => \N__11434\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11427\
        );

    \I__2223\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11418\
        );

    \I__2222\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11418\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11418\
        );

    \I__2220\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11415\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11418\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__11415\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__11410\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11404\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__11404\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__2214\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__11398\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__2211\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__11389\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__11386\,
            I => \N__11383\
        );

    \I__2208\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11380\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11377\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__11377\,
            I => \CO4_1\
        );

    \I__2205\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11371\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__11371\,
            I => \N__11368\
        );

    \I__2203\ : Odrv12
    port map (
            O => \N__11368\,
            I => \row_1_if_generate_plus_mult1_un47_sum_cZ0Z5\
        );

    \I__2202\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__11356\,
            I => content_ram8_0
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__11347\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28\
        );

    \I__2195\ : InMux
    port map (
            O => \N__11344\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2194\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11338\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__11338\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__2192\ : InMux
    port map (
            O => \N__11335\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__2191\ : InMux
    port map (
            O => \N__11332\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__11329\,
            I => \N__11324\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__11328\,
            I => \N__11320\
        );

    \I__2188\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11316\
        );

    \I__2187\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11307\
        );

    \I__2186\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11307\
        );

    \I__2185\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11307\
        );

    \I__2184\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11307\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__11316\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__11307\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__11302\,
            I => \N__11299\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11296\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__11296\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__2178\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__11290\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2\
        );

    \I__2176\ : InMux
    port map (
            O => \N__11287\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__2174\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__11278\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11275\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__11266\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3\
        );

    \I__2168\ : InMux
    port map (
            O => \N__11263\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__11260\,
            I => \un5_beamx_2_0_cascade_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__11254\,
            I => un5_beamx_3
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__11251\,
            I => \un5_visibley_ac0_11_0_1_cascade_\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \N__11245\
        );

    \I__2162\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11242\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__11242\,
            I => \beamY_RNI8325_0Z0Z_6\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__11239\,
            I => \N__11235\
        );

    \I__2159\ : InMux
    port map (
            O => \N__11238\,
            I => \N__11230\
        );

    \I__2158\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11230\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11225\
        );

    \I__2156\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11222\
        );

    \I__2155\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11219\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__11225\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__11222\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__11219\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__11212\,
            I => \N__11209\
        );

    \I__2150\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11206\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__11206\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4\
        );

    \I__2148\ : InMux
    port map (
            O => \N__11203\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__2147\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11197\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__11197\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7\
        );

    \I__2145\ : InMux
    port map (
            O => \N__11194\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__11191\,
            I => \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\
        );

    \I__2143\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__11185\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__2140\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11171\
        );

    \I__2139\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11171\
        );

    \I__2138\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11168\
        );

    \I__2137\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11164\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__11171\,
            I => \N__11159\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11159\
        );

    \I__2134\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11156\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11152\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__11159\,
            I => \N__11147\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__11156\,
            I => \N__11147\
        );

    \I__2130\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11144\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__11152\,
            I => \beamY_RNIVMI9D5Z0Z_3\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__11147\,
            I => \beamY_RNIVMI9D5Z0Z_3\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__11144\,
            I => \beamY_RNIVMI9D5Z0Z_3\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__11137\,
            I => \N__11134\
        );

    \I__2125\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11131\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__11131\,
            I => un5_visibley_1_29
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11124\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__11127\,
            I => \N__11120\
        );

    \I__2121\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11116\
        );

    \I__2120\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11111\
        );

    \I__2119\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11111\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__11119\,
            I => \N__11106\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__11116\,
            I => \N__11103\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__11111\,
            I => \N__11100\
        );

    \I__2115\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11095\
        );

    \I__2114\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11095\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11092\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__11103\,
            I => \N__11085\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__11100\,
            I => \N__11085\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__11095\,
            I => \N__11085\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__11092\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__11085\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \beamY_RNI8325Z0Z_6_cascade_\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__11077\,
            I => \un5_visibley_c5_cascade_\
        );

    \I__2105\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__11071\,
            I => un1_beamylto9_1
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \un5_visibley_c3_cascade_\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__11065\,
            I => \content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11059\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__11059\,
            I => \content_content_ram9__e_0_RNIFBHPN1Z0Z_0\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__11056\,
            I => \N__11053\
        );

    \I__2098\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11050\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__11050\,
            I => \content_content_ram5__RNIEM2QF3Z0Z_0\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__11047\,
            I => \N__11044\
        );

    \I__2095\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__2094\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11038\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__11038\,
            I => content_ram9_0
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__11035\,
            I => \N__11031\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__11034\,
            I => \N__11028\
        );

    \I__2090\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11023\
        );

    \I__2089\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11023\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__11023\,
            I => content_ram11_0
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__11020\,
            I => \N__11016\
        );

    \I__2086\ : IoInMux
    port map (
            O => \N__11019\,
            I => \N__11013\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__11008\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11008\
        );

    \I__2083\ : IoSpan4Mux
    port map (
            O => \N__11008\,
            I => \N__11005\
        );

    \I__2082\ : Span4Mux_s2_h
    port map (
            O => \N__11005\,
            I => \N__11001\
        );

    \I__2081\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10998\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__11001\,
            I => \nCS1_c\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10998\,
            I => \nCS1_c\
        );

    \I__2078\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10987\
        );

    \I__2077\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10987\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__10987\,
            I => un5_visibley_2_28
        );

    \I__2075\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10981\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__10981\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__2073\ : InMux
    port map (
            O => \N__10978\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__2072\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10969\
        );

    \I__2071\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10969\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10969\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0\
        );

    \I__2069\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10963\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__10963\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0\
        );

    \I__2067\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10957\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__10957\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__10954\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10947\
        );

    \I__2063\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10944\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__10947\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__10944\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0\
        );

    \I__2060\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10936\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N__10933\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__10930\,
            I => chessboardpixel_un178_pixel_26
        );

    \I__2056\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10924\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__10924\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__2054\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10918\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10915\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__10915\,
            I => \N__10912\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__10912\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z5\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__10909\,
            I => \N__10906\
        );

    \I__2049\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10903\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__10903\,
            I => \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3\
        );

    \I__2047\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10896\
        );

    \I__2046\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10893\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10890\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10887\
        );

    \I__2043\ : Span4Mux_h
    port map (
            O => \N__10890\,
            I => \N__10882\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__10887\,
            I => \N__10879\
        );

    \I__2041\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10874\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10874\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__10882\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__10879\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__10874\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__10867\,
            I => \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10861\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__10861\,
            I => \N__10858\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__10858\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__10855\,
            I => \chessboardpixel_un200_pixellto4_1_cascade_\
        );

    \I__2031\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10849\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__10846\,
            I => \N__10843\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__10843\,
            I => chessboardpixel_un200_pixellt10
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__10840\,
            I => \N__10835\
        );

    \I__2026\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10832\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10829\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10826\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__10832\,
            I => un8_beamy_3
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__10829\,
            I => un8_beamy_3
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__10826\,
            I => un8_beamy_3
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__10819\,
            I => \beamY_i_2_cascade_\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__10816\,
            I => \N__10811\
        );

    \I__2018\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10807\
        );

    \I__2017\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10802\
        );

    \I__2016\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10802\
        );

    \I__2015\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10799\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__10807\,
            I => \beamY_i_2\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__10802\,
            I => \beamY_i_2\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__10799\,
            I => \beamY_i_2\
        );

    \I__2011\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10786\
        );

    \I__2010\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10786\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__10786\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0\
        );

    \I__2008\ : InMux
    port map (
            O => \N__10783\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__2007\ : InMux
    port map (
            O => \N__10780\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__2006\ : InMux
    port map (
            O => \N__10777\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__2005\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10771\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10771\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__10768\,
            I => \g2_0_cascade_\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__10765\,
            I => \N__10762\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10759\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10756\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__10756\,
            I => chary_if_generate_plus_mult1_un68_sum_1_5
        );

    \I__1998\ : IoInMux
    port map (
            O => \N__10753\,
            I => \N__10750\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__10750\,
            I => \N__10747\
        );

    \I__1996\ : Span4Mux_s3_v
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__10744\,
            I => \VSync_c\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__10741\,
            I => \N__10738\
        );

    \I__1993\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10735\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__10735\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__10732\,
            I => \N__10729\
        );

    \I__1990\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10726\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__10726\,
            I => un5_visibley_3_28
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__10723\,
            I => \un5_visibley_3_28_cascade_\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__10720\,
            I => \g1_3_cascade_\
        );

    \I__1986\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10714\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__10714\,
            I => g2_0_1
        );

    \I__1984\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10708\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10705\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__10705\,
            I => un1_beamylto9_2
        );

    \I__1981\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10696\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10696\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__10696\,
            I => un5_visibley_1_28
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__10693\,
            I => \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10687\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__10687\,
            I => chary_if_generate_plus_mult1_un68_sum_2_5
        );

    \I__1975\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10681\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__10681\,
            I => un5_visibley_2_29
        );

    \I__1973\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10675\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__10675\,
            I => g2_0_0
        );

    \I__1971\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10669\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__10669\,
            I => \beamY_RNIMSO1N7Z0Z_2\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__10666\,
            I => \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_\
        );

    \I__1968\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10660\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__10660\,
            I => \N__10657\
        );

    \I__1966\ : Odrv12
    port map (
            O => \N__10657\,
            I => chary_if_generate_plus_mult1_un68_sum_1_0_5
        );

    \I__1965\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10651\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10648\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__10648\,
            I => g2_0
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__10645\,
            I => \N__10642\
        );

    \I__1961\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10639\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__10639\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__1959\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10633\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__10633\,
            I => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__1957\ : InMux
    port map (
            O => \N__10630\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__1956\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10624\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__10624\,
            I => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10621\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__10618\,
            I => \content_column_1_i_2_2_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10611\
        );

    \I__1951\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10608\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__10611\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10608\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__10603\,
            I => \N__10600\
        );

    \I__1947\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10597\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__10597\,
            I => if_generate_plus_mult1_un75_sum_axb_4_l_fx
        );

    \I__1945\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10586\
        );

    \I__1944\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10586\
        );

    \I__1943\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10582\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__10591\,
            I => \N__10579\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10576\
        );

    \I__1940\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10573\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10570\
        );

    \I__1938\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10567\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__10576\,
            I => \N__10564\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10561\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__10570\,
            I => \N__10556\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__10567\,
            I => \N__10556\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__10564\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__10561\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__10556\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__1930\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10546\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__10546\,
            I => \column_1_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__10543\,
            I => \content_m7_ns_1_cascade_\
        );

    \I__1927\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10533\
        );

    \I__1926\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10533\
        );

    \I__1925\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10530\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10533\,
            I => \N__10527\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__10530\,
            I => \N__10524\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__10524\,
            I => \N__10518\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__10521\,
            I => \content_N_8\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__10518\,
            I => \content_N_8\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__10513\,
            I => \content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10507\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10504\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__10504\,
            I => \content_content_ram7__RNI6B0NG3Z0Z_0\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__10498\,
            I => \content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__10495\,
            I => \N__10492\
        );

    \I__1911\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10489\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__10489\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__1909\ : InMux
    port map (
            O => \N__10486\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__1908\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10480\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__10480\,
            I => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__1906\ : InMux
    port map (
            O => \N__10477\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__1905\ : InMux
    port map (
            O => \N__10474\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__10471\,
            I => \N__10468\
        );

    \I__1903\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10465\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__10465\,
            I => content_column_1_i_2_i_2
        );

    \I__1901\ : InMux
    port map (
            O => \N__10462\,
            I => \N__10454\
        );

    \I__1900\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10454\
        );

    \I__1899\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10449\
        );

    \I__1898\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10449\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10440\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__10449\,
            I => \N__10440\
        );

    \I__1895\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10437\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10432\
        );

    \I__1893\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10432\
        );

    \I__1892\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10429\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__10440\,
            I => un6_rowlto1
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__10437\,
            I => un6_rowlto1
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__10432\,
            I => un6_rowlto1
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__10429\,
            I => un6_rowlto1
        );

    \I__1887\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10414\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10411\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__10411\,
            I => \N__10408\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__10408\,
            I => \content_N_25\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__10405\,
            I => \N__10402\
        );

    \I__1881\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10399\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__10399\,
            I => \column_1_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__10396\,
            I => \N__10393\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10390\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__10390\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__1876\ : InMux
    port map (
            O => \N__10387\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__10384\,
            I => \N__10381\
        );

    \I__1874\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10378\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10378\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__1872\ : InMux
    port map (
            O => \N__10375\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__1871\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__1870\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10366\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__10366\,
            I => column_1_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__1868\ : IoInMux
    port map (
            O => \N__10363\,
            I => \N__10360\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__10360\,
            I => \N__10357\
        );

    \I__1866\ : IoSpan4Mux
    port map (
            O => \N__10357\,
            I => \N__10354\
        );

    \I__1865\ : Sp12to4
    port map (
            O => \N__10354\,
            I => \N__10351\
        );

    \I__1864\ : Span12Mux_s7_v
    port map (
            O => \N__10351\,
            I => \N__10348\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__10348\,
            I => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__10345\,
            I => \N__10338\
        );

    \I__1861\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10334\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \N__10331\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__10342\,
            I => \N__10327\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10341\,
            I => \N__10323\
        );

    \I__1857\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10318\
        );

    \I__1856\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10318\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10315\
        );

    \I__1854\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10308\
        );

    \I__1853\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10308\
        );

    \I__1852\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10308\
        );

    \I__1851\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10305\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10300\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10300\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__10315\,
            I => \N__10297\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__10308\,
            I => \N__10292\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__10305\,
            I => \N__10292\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__10300\,
            I => \N__10289\
        );

    \I__1844\ : Span4Mux_h
    port map (
            O => \N__10297\,
            I => \N__10284\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__10292\,
            I => \N__10284\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__10289\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__10284\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__1840\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10273\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10273\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__10273\,
            I => \G_383\
        );

    \I__1837\ : InMux
    port map (
            O => \N__10270\,
            I => column_1_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__1836\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10257\
        );

    \I__1835\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10257\
        );

    \I__1834\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10257\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__10264\,
            I => \N__10254\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__10257\,
            I => \N__10250\
        );

    \I__1831\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10245\
        );

    \I__1830\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10245\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__10250\,
            I => un6_rowlto0
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__10245\,
            I => un6_rowlto0
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__10240\,
            I => \N__10237\
        );

    \I__1826\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__10234\,
            I => \column_1_if_generate_plus_mult1_un75_sum_iZ0\
        );

    \I__1824\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10227\
        );

    \I__1823\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10224\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__10227\,
            I => \N__10218\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10218\
        );

    \I__1820\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10215\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__10218\,
            I => \N__10209\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__10215\,
            I => \N__10209\
        );

    \I__1817\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10206\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__10209\,
            I => \N__10201\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__10206\,
            I => \N__10201\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__10201\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__10192\,
            I => if_generate_plus_mult1_un75_sum_cry_2_s
        );

    \I__1810\ : InMux
    port map (
            O => \N__10189\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \N__10182\
        );

    \I__1808\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10177\
        );

    \I__1807\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10177\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10177\,
            I => un5_visibley_0_28
        );

    \I__1805\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10171\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__10171\,
            I => g2
        );

    \I__1803\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10165\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10162\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__10162\,
            I => un5_visibley_0_29
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__10159\,
            I => \N__10156\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10153\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10153\,
            I => \N__10150\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__10150\,
            I => \Pixel_RNOZ0Z_67\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__10147\,
            I => \un4_beamylt6_cascade_\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__10144\,
            I => \N__10141\
        );

    \I__1794\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10138\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__10138\,
            I => \N__10135\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__10135\,
            I => un4_beamylt8_0
        );

    \I__1791\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10129\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__10129\,
            I => chary_0_24
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__10126\,
            I => \N__10121\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10112\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10112\
        );

    \I__1786\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10107\
        );

    \I__1785\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10107\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10100\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10100\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10100\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__10112\,
            I => chary_if_generate_plus_mult1_un75_sum_axbxc5_1
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__10107\,
            I => chary_if_generate_plus_mult1_un75_sum_axbxc5_1
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__10100\,
            I => chary_if_generate_plus_mult1_un75_sum_axbxc5_1
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__10093\,
            I => \chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_\
        );

    \I__1777\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10087\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10087\,
            I => g1_2_0
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__10084\,
            I => \beamY_RNIMSO1N7_0Z0Z_2_cascade_\
        );

    \I__1774\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10075\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10075\,
            I => g4_0
        );

    \I__1771\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10069\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10069\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \g2_1_0_cascade_\
        );

    \I__1768\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__10060\,
            I => chary_if_generate_plus_mult1_un68_sum_0_5
        );

    \I__1766\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10054\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__10054\,
            I => \Pixel_RNOZ0Z_66\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__1763\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10045\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10042\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__10042\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__1760\ : InMux
    port map (
            O => \N__10039\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__10036\,
            I => \N__10033\
        );

    \I__1758\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10030\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__10030\,
            I => \N__10027\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__10027\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__1755\ : InMux
    port map (
            O => \N__10024\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__1754\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10018\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__10015\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__10015\,
            I => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__1751\ : InMux
    port map (
            O => \N__10012\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__10009\,
            I => \if_generate_plus_mult1_un61_sum_s_5_cascade_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9998\
        );

    \I__1748\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9998\
        );

    \I__1747\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9992\
        );

    \I__1746\ : InMux
    port map (
            O => \N__10003\,
            I => \N__9989\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9986\
        );

    \I__1744\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9983\
        );

    \I__1743\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9978\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9978\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9992\,
            I => \N__9973\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9973\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__9986\,
            I => \N__9970\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__9983\,
            I => \N__9967\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__9978\,
            I => \N__9964\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__9973\,
            I => \N__9961\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__9970\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__9967\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__1733\ : Odrv12
    port map (
            O => \N__9964\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__9961\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__1731\ : InMux
    port map (
            O => \N__9952\,
            I => \N__9946\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9943\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9940\
        );

    \I__1728\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9937\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__9946\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__9943\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__9940\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__9937\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__1723\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9925\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__9925\,
            I => column_1_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__1721\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9919\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__9919\,
            I => \N__9916\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__9916\,
            I => \N__9913\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__9913\,
            I => chary_2_24
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__9910\,
            I => \N__9906\
        );

    \I__1716\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9903\
        );

    \I__1715\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9898\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__9903\,
            I => \N__9895\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9891\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__9901\,
            I => \N__9888\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9898\,
            I => \N__9884\
        );

    \I__1710\ : Span12Mux_s5_h
    port map (
            O => \N__9895\,
            I => \N__9881\
        );

    \I__1709\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9878\
        );

    \I__1708\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9875\
        );

    \I__1707\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9870\
        );

    \I__1706\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9870\
        );

    \I__1705\ : Span12Mux_s5_h
    port map (
            O => \N__9884\,
            I => \N__9867\
        );

    \I__1704\ : Odrv12
    port map (
            O => \N__9881\,
            I => \beamY_RNI539IG9Z0Z_3\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__9878\,
            I => \beamY_RNI539IG9Z0Z_3\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__9875\,
            I => \beamY_RNI539IG9Z0Z_3\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__9870\,
            I => \beamY_RNI539IG9Z0Z_3\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__9867\,
            I => \beamY_RNI539IG9Z0Z_3\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__9856\,
            I => \beamY_RNI539IG9Z0Z_3_cascade_\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9850\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__9850\,
            I => g4
        );

    \I__1696\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9843\
        );

    \I__1695\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9836\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__9843\,
            I => \N__9833\
        );

    \I__1693\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9830\
        );

    \I__1692\ : InMux
    port map (
            O => \N__9841\,
            I => \N__9827\
        );

    \I__1691\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9824\
        );

    \I__1690\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9821\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9818\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9813\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9813\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__9827\,
            I => \N__9808\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__9824\,
            I => \N__9808\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9805\
        );

    \I__1683\ : Span4Mux_h
    port map (
            O => \N__9818\,
            I => \N__9802\
        );

    \I__1682\ : Span4Mux_h
    port map (
            O => \N__9813\,
            I => \N__9799\
        );

    \I__1681\ : Odrv12
    port map (
            O => \N__9808\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__9805\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__9802\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__9799\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__9790\,
            I => \N__9787\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9784\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__1674\ : Odrv12
    port map (
            O => \N__9781\,
            I => charx_if_generate_plus_mult1_un40_sum_i
        );

    \I__1673\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__9775\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\
        );

    \I__1671\ : InMux
    port map (
            O => \N__9772\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__1670\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9765\
        );

    \I__1669\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9762\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__9765\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9762\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__1665\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__9751\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__9748\,
            I => \N__9744\
        );

    \I__1662\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9739\
        );

    \I__1661\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9739\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__9739\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\
        );

    \I__1659\ : InMux
    port map (
            O => \N__9736\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__1658\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__1657\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9727\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__9727\,
            I => charx_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__9724\,
            I => \N__9721\
        );

    \I__1654\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__9718\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\
        );

    \I__1652\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9712\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__9712\,
            I => charx_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__1650\ : InMux
    port map (
            O => \N__9709\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__1649\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9703\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__9703\,
            I => charx_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__1647\ : InMux
    port map (
            O => \N__9700\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__9697\,
            I => \N__9693\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9689\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9693\,
            I => \N__9684\
        );

    \I__1643\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9684\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__9689\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__9684\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__9679\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\
        );

    \I__1639\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__9673\,
            I => charx_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__1637\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__9667\,
            I => un5_visiblex_i_27
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__1634\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9658\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__9658\,
            I => \N__9654\
        );

    \I__1632\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9651\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__9654\,
            I => \column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__9651\,
            I => \column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO\
        );

    \I__1629\ : InMux
    port map (
            O => \N__9646\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__1628\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__9640\,
            I => \content_content_ram0__RNIR1C2R81_0Z0Z_0\
        );

    \I__1626\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9634\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__9634\,
            I => un6_rowlt7_0
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1623\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__9622\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\
        );

    \I__1620\ : InMux
    port map (
            O => \N__9619\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__1618\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__9607\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\
        );

    \I__1615\ : InMux
    port map (
            O => \N__9604\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__1614\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__9595\,
            I => charx_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__1611\ : InMux
    port map (
            O => \N__9592\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__1610\ : InMux
    port map (
            O => \N__9589\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1609\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9583\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9578\
        );

    \I__1607\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9575\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9572\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__9578\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__9575\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__9572\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__9565\,
            I => \N__9562\
        );

    \I__1601\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9559\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__9559\,
            I => charx_if_generate_plus_mult1_un47_sum_i
        );

    \I__1599\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9553\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__9553\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\
        );

    \I__1597\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9547\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__9547\,
            I => g4_1
        );

    \I__1595\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9541\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__9541\,
            I => \N__9538\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__9538\,
            I => \N__9535\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__9535\,
            I => g0_0_a3_5
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__9532\,
            I => \m4_rn_1_cascade_\
        );

    \I__1590\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__9523\,
            I => \N__9520\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__9520\,
            I => \Pixel_RNOZ0Z_40\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__9517\,
            I => \content_content_ram0__RNIR1C2R81Z0Z_0_cascade_\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9505\
        );

    \I__1584\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9499\
        );

    \I__1583\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9496\
        );

    \I__1582\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9493\
        );

    \I__1581\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9488\
        );

    \I__1580\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9483\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9483\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9480\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9473\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9473\
        );

    \I__1575\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9473\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9468\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__9496\,
            I => \N__9468\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__9493\,
            I => \N__9464\
        );

    \I__1571\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9459\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9459\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__9488\,
            I => \N__9455\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9446\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__9480\,
            I => \N__9446\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9446\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__9468\,
            I => \N__9446\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9443\
        );

    \I__1563\ : Span4Mux_s3_v
    port map (
            O => \N__9464\,
            I => \N__9438\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__9459\,
            I => \N__9438\
        );

    \I__1561\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9435\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__9455\,
            I => \N_331_i\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__9446\,
            I => \N_331_i\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N_331_i\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__9438\,
            I => \N_331_i\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__9435\,
            I => \N_331_i\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__9424\,
            I => \un4_row_m7_ns_1_cascade_\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__9421\,
            I => \N__9418\
        );

    \I__1553\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9415\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9415\,
            I => \beamY_RNIPAQ91Z0Z_6\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9409\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__9409\,
            I => un4_beamy_0
        );

    \I__1549\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9403\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__9403\,
            I => m4_sn
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__9400\,
            I => \chary_1_24_cascade_\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9394\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N_1737_0\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \chary_1_0_24_cascade_\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__9388\,
            I => \g2_3_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9382\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__9382\,
            I => g1_1_1
        );

    \I__1540\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__9376\,
            I => un116_pixel_0_0_0
        );

    \I__1538\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9370\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__9370\,
            I => \N_5_1\
        );

    \I__1536\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__9361\,
            I => \N__9358\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__9358\,
            I => g0_0_a3_4
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__9355\,
            I => \un8_beamylto9_1_cascade_\
        );

    \I__1531\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__9349\,
            I => un8_beamy
        );

    \I__1529\ : InMux
    port map (
            O => \N__9346\,
            I => \N__9343\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__9343\,
            I => \N_134_0\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__9340\,
            I => \font_un28_pixel_29_cascade_\
        );

    \I__1526\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__9331\,
            I => \beamY_RNIDA2GGA3Z0Z_0\
        );

    \I__1523\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9325\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__9325\,
            I => \N__9322\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__9322\,
            I => g0_1
        );

    \I__1520\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9312\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9309\
        );

    \I__1518\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9300\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9300\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__9315\,
            I => \N__9297\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9291\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9309\,
            I => \N__9288\
        );

    \I__1513\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9285\
        );

    \I__1512\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9278\
        );

    \I__1511\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9278\
        );

    \I__1510\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9278\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__9300\,
            I => \N__9275\
        );

    \I__1508\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9270\
        );

    \I__1507\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9270\
        );

    \I__1506\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9265\
        );

    \I__1505\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9265\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__9291\,
            I => \N__9262\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__9288\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__9285\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__9278\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__9275\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__9270\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__9265\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__9262\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__9247\,
            I => \beamY_RNIDA2GGA3Z0Z_0_cascade_\
        );

    \I__1495\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N_19_0_0\
        );

    \I__1493\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__9235\,
            I => font_un28_pixel_30
        );

    \I__1491\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9228\
        );

    \I__1490\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9225\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9222\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__9225\,
            I => font_un28_pixel_29
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__9222\,
            I => font_un28_pixel_29
        );

    \I__1486\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N_15_i\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \Pixel_RNOZ0Z_28_cascade_\
        );

    \I__1483\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__9205\,
            I => \N__9202\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__9202\,
            I => \Pixel_RNOZ0Z_9\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9193\
        );

    \I__1479\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9193\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9189\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9185\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__9189\,
            I => \N__9182\
        );

    \I__1475\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9179\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__9185\,
            I => chary_24
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__9182\,
            I => chary_24
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__9179\,
            I => chary_24
        );

    \I__1471\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9169\,
            I => \N__9165\
        );

    \I__1469\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9161\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__9165\,
            I => \N__9158\
        );

    \I__1467\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9155\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9152\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__9158\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__9155\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__9152\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__1461\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9139\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__9139\,
            I => charx_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__1459\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9127\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9127\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__9134\,
            I => \N__9123\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__9133\,
            I => \N__9120\
        );

    \I__1455\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9116\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9113\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9110\
        );

    \I__1452\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9105\
        );

    \I__1451\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9105\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9101\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__9116\,
            I => \N__9095\
        );

    \I__1448\ : Span4Mux_h
    port map (
            O => \N__9113\,
            I => \N__9092\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9087\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__9105\,
            I => \N__9087\
        );

    \I__1445\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9084\
        );

    \I__1444\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9081\
        );

    \I__1443\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9074\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9074\
        );

    \I__1441\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9074\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__9095\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__9092\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__9087\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__9084\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9081\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__9074\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__9061\,
            I => \N__9058\
        );

    \I__1433\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__9055\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__1431\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__9049\,
            I => \N__9046\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__9046\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\
        );

    \I__1428\ : InMux
    port map (
            O => \N__9043\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__1427\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9033\
        );

    \I__1426\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9033\
        );

    \I__1425\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9030\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__9033\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9030\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\
        );

    \I__1422\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9019\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9019\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__9019\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8
        );

    \I__1419\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__9010\
        );

    \I__1417\ : Odrv12
    port map (
            O => \N__9010\,
            I => \Pixel_RNOZ0Z_14\
        );

    \I__1416\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__9001\,
            I => font_un126_pixel_5_a0_1
        );

    \I__1413\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8992\
        );

    \I__1411\ : Span12Mux_s3_v
    port map (
            O => \N__8992\,
            I => \N__8989\
        );

    \I__1410\ : Odrv12
    port map (
            O => \N__8989\,
            I => \N_1740_0\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__8986\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_\
        );

    \I__1408\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8980\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__8980\,
            I => \N__8974\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8969\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8969\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8964\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__8974\,
            I => \N__8956\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8956\
        );

    \I__1401\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8953\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__8967\,
            I => \N__8950\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__8964\,
            I => \N__8947\
        );

    \I__1398\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8940\
        );

    \I__1397\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8940\
        );

    \I__1396\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8940\
        );

    \I__1395\ : Span4Mux_h
    port map (
            O => \N__8956\,
            I => \N__8937\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8934\
        );

    \I__1393\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8931\
        );

    \I__1392\ : Odrv12
    port map (
            O => \N__8947\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8940\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__8937\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__1389\ : Odrv12
    port map (
            O => \N__8934\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__8931\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__8920\,
            I => \N__8917\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8914\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__8914\,
            I => charx_if_generate_plus_mult1_un33_sum_i
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__8911\,
            I => \N__8908\
        );

    \I__1383\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8895\
        );

    \I__1382\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8895\
        );

    \I__1381\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8895\
        );

    \I__1380\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8888\
        );

    \I__1379\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8888\
        );

    \I__1378\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8888\
        );

    \I__1377\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8885\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8880\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__8888\,
            I => \N__8880\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8885\,
            I => \N__8875\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__8880\,
            I => \N__8872\
        );

    \I__1372\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8869\
        );

    \I__1371\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8866\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__8875\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__8872\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__8869\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__8866\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__8857\,
            I => \N__8854\
        );

    \I__1365\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__8851\,
            I => \N__8848\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__8848\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\
        );

    \I__1362\ : InMux
    port map (
            O => \N__8845\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__8842\,
            I => \N__8839\
        );

    \I__1360\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8836\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__8830\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__1355\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__8821\,
            I => \N__8818\
        );

    \I__1353\ : Odrv12
    port map (
            O => \N__8818\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\
        );

    \I__1352\ : InMux
    port map (
            O => \N__8815\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__8812\,
            I => \N__8809\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__8800\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\
        );

    \I__1346\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8794\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__8791\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__1343\ : InMux
    port map (
            O => \N__8788\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__1342\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8782\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8779\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__8779\,
            I => \N__8776\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__8776\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__1338\ : InMux
    port map (
            O => \N__8773\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__1337\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8767\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8762\
        );

    \I__1335\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8759\
        );

    \I__1334\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8756\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__8762\,
            I => \N__8751\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8751\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__8756\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__8751\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\
        );

    \I__1329\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8743\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__8743\,
            I => un4_row_9_0
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__8740\,
            I => \N__8737\
        );

    \I__1326\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8734\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__8731\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__1323\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8723\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8718\
        );

    \I__1321\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8718\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__8723\,
            I => \column_1_if_generate_plus_mult1_un47_sum_cZ0Z5\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__8718\,
            I => \column_1_if_generate_plus_mult1_un47_sum_cZ0Z5\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__8713\,
            I => \N__8710\
        );

    \I__1317\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8707\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__8707\,
            I => \N__8701\
        );

    \I__1315\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8698\
        );

    \I__1314\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8692\
        );

    \I__1313\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8692\
        );

    \I__1312\ : Span4Mux_v
    port map (
            O => \N__8701\,
            I => \N__8686\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__8698\,
            I => \N__8686\
        );

    \I__1310\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8680\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__8692\,
            I => \N__8677\
        );

    \I__1308\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8674\
        );

    \I__1307\ : Span4Mux_h
    port map (
            O => \N__8686\,
            I => \N__8671\
        );

    \I__1306\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8664\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8664\
        );

    \I__1304\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8664\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8661\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__8677\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__8674\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__8671\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__8664\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__8661\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__1297\ : InMux
    port map (
            O => \N__8650\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1295\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__8635\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8632\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__8629\,
            I => \N__8626\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8623\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8620\
        );

    \I__1287\ : Span4Mux_h
    port map (
            O => \N__8620\,
            I => \N__8617\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__8617\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8614\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__1284\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1282\ : Span4Mux_h
    port map (
            O => \N__8605\,
            I => \N__8602\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__8602\,
            I => charx_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__1280\ : InMux
    port map (
            O => \N__8599\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__1279\ : InMux
    port map (
            O => \N__8596\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__1278\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8590\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__8587\,
            I => \N__8584\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__8584\,
            I => if_generate_plus_mult1_un54_sum_axb_3_l_ofx
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1273\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8575\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__8575\,
            I => \N__8572\
        );

    \I__1271\ : Span4Mux_h
    port map (
            O => \N__8572\,
            I => \N__8569\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__8569\,
            I => \column_1_if_generate_plus_mult1_un47_sum_c5_iZ0\
        );

    \I__1269\ : InMux
    port map (
            O => \N__8566\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__8563\,
            I => \N__8560\
        );

    \I__1267\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1265\ : Span4Mux_h
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__8551\,
            I => if_generate_plus_mult1_un54_sum_axb_4_l_ofx
        );

    \I__1263\ : InMux
    port map (
            O => \N__8548\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__1262\ : InMux
    port map (
            O => \N__8545\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1261\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8536\
        );

    \I__1260\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8536\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8533\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__8533\,
            I => charx_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__1256\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8524\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__8524\,
            I => un5_visiblex_i_26
        );

    \I__1254\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8515\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__8515\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__8512\,
            I => \un4_row_9_2_cascade_\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8506\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8503\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__8503\,
            I => un4_row_9_5
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__8500\,
            I => \N__8496\
        );

    \I__1246\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8491\
        );

    \I__1245\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8491\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__8491\,
            I => \N__8488\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__8488\,
            I => \N__8483\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8478\
        );

    \I__1241\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8478\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__8483\,
            I => \N__8475\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__8478\,
            I => \beamXZ0Z_10\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__8475\,
            I => \beamXZ0Z_10\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8466\
        );

    \I__1236\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8462\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8459\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8456\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8451\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__8459\,
            I => \N__8451\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8448\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__8451\,
            I => \N__8445\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__8448\,
            I => un1_beamx_2
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__8445\,
            I => un1_beamx_2
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__8440\,
            I => \N__8436\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__8439\,
            I => \N__8431\
        );

    \I__1225\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8424\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8424\
        );

    \I__1223\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8421\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8417\
        );

    \I__1221\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8414\
        );

    \I__1220\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8411\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__8424\,
            I => \N__8406\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__8421\,
            I => \N__8406\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__8420\,
            I => \N__8402\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8397\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8397\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8394\
        );

    \I__1213\ : Span4Mux_s2_v
    port map (
            O => \N__8406\,
            I => \N__8391\
        );

    \I__1212\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8387\
        );

    \I__1211\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8384\
        );

    \I__1210\ : Span12Mux_s9_v
    port map (
            O => \N__8397\,
            I => \N__8381\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__8394\,
            I => \N__8376\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__8391\,
            I => \N__8376\
        );

    \I__1207\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8373\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__8387\,
            I => \beamXZ0Z_7\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__8384\,
            I => \beamXZ0Z_7\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__8381\,
            I => \beamXZ0Z_7\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__8376\,
            I => \beamXZ0Z_7\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__8373\,
            I => \beamXZ0Z_7\
        );

    \I__1201\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8359\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8356\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__8356\,
            I => un1_beamxlt10_0
        );

    \I__1198\ : IoInMux
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1196\ : Span4Mux_s3_v
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1195\ : Span4Mux_h
    port map (
            O => \N__8344\,
            I => \N__8341\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__8341\,
            I => \HSync_c\
        );

    \I__1193\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8331\
        );

    \I__1191\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8328\
        );

    \I__1190\ : Span4Mux_s2_v
    port map (
            O => \N__8331\,
            I => \N__8322\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8328\,
            I => \N__8319\
        );

    \I__1188\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8314\
        );

    \I__1187\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8314\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8311\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__8322\,
            I => \N__8308\
        );

    \I__1184\ : Span4Mux_s3_h
    port map (
            O => \N__8319\,
            I => \N__8303\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8303\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8300\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__8308\,
            I => un4_row
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__8303\,
            I => un4_row
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__8300\,
            I => un4_row
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1177\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__8284\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8281\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1172\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__8269\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\
        );

    \I__1169\ : InMux
    port map (
            O => \N__8266\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__1168\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__8257\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__1165\ : InMux
    port map (
            O => \N__8254\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__1164\ : InMux
    port map (
            O => \N__8251\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__1163\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8245\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8240\
        );

    \I__1161\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8237\
        );

    \I__1160\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8234\
        );

    \I__1159\ : Span4Mux_s1_h
    port map (
            O => \N__8240\,
            I => \N__8227\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__8237\,
            I => \N__8227\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8227\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__8227\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__8224\,
            I => \beamY_RNINKIU27Z0Z_0_cascade_\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__8221\,
            I => \Pixel_RNOZ0Z_29_cascade_\
        );

    \I__1153\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N_10\
        );

    \I__1151\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__8206\,
            I => chessboardpixel_un152_pixel_27
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__8203\,
            I => \N__8200\
        );

    \I__1147\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8194\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__8194\,
            I => chessboardpixel_un174_pixellt10
        );

    \I__1144\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__8188\,
            I => \N__8185\
        );

    \I__1142\ : Span4Mux_s3_h
    port map (
            O => \N__8185\,
            I => \N__8180\
        );

    \I__1141\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8175\
        );

    \I__1140\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8175\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__8180\,
            I => chessboardpixel_un175_pixel
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8175\,
            I => chessboardpixel_un175_pixel
        );

    \I__1137\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8167\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__8161\,
            I => g1_2_1
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \chessboardpixel_un175_pixel_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8152\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1130\ : Span4Mux_s3_h
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__8146\,
            I => g2_3_0_0
        );

    \I__1128\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8136\
        );

    \I__1127\ : InMux
    port map (
            O => \N__8142\,
            I => \N__8136\
        );

    \I__1126\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8133\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__8136\,
            I => \N__8130\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__8133\,
            I => \N__8127\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__8130\,
            I => un13_beamylt7
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__8127\,
            I => un13_beamylt7
        );

    \I__1121\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8118\
        );

    \I__1120\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8115\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8118\,
            I => un15_beamy
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__8115\,
            I => un15_beamy
        );

    \I__1117\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8107\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__8104\,
            I => un18_beamylt10_0
        );

    \I__1114\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8097\
        );

    \I__1113\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__8097\,
            I => \N__8089\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8089\
        );

    \I__1110\ : Span4Mux_s3_h
    port map (
            O => \N__8089\,
            I => \N__8084\
        );

    \I__1109\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8079\
        );

    \I__1108\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8079\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__8084\,
            I => un15_beamy_2
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__8079\,
            I => un15_beamy_2
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__8074\,
            I => \Pixel_RNOZ0Z_44_cascade_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1102\ : Span12Mux_s3_h
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__8062\,
            I => \N_10_0_0\
        );

    \I__1100\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__8050\,
            I => \N_20\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__8047\,
            I => \g0_4_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8041\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8038\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__8038\,
            I => \G_21_i_2\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__8032\,
            I => \N__8029\
        );

    \I__1090\ : Span4Mux_s1_v
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__8026\,
            I => \N__8023\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__8023\,
            I => \Pixel_c\
        );

    \I__1087\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__8017\,
            I => g1_1_0
        );

    \I__1085\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__8008\,
            I => g0_2_0
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__8005\,
            I => \g1_1_cascade_\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__7999\,
            I => g3_1
        );

    \I__1079\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__7993\,
            I => g0_5
        );

    \I__1077\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7986\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7983\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__7986\,
            I => g1_0_0
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__7983\,
            I => g1_0_0
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7972\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__7972\,
            I => \N__7969\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__7969\,
            I => g0_0_a3_0
        );

    \I__1069\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7957\
        );

    \I__1068\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7952\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7952\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__7963\,
            I => \N__7949\
        );

    \I__1065\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7945\
        );

    \I__1064\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7940\
        );

    \I__1063\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7940\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__7957\,
            I => \N__7934\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7934\
        );

    \I__1060\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7931\
        );

    \I__1059\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7927\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__7945\,
            I => \N__7922\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7922\
        );

    \I__1056\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7919\
        );

    \I__1055\ : Span4Mux_s2_v
    port map (
            O => \N__7934\,
            I => \N__7914\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7914\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__7930\,
            I => \N__7910\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7903\
        );

    \I__1051\ : Span4Mux_s2_v
    port map (
            O => \N__7922\,
            I => \N__7903\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__7919\,
            I => \N__7903\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__7914\,
            I => \N__7900\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \N__7896\
        );

    \I__1047\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7890\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__7903\,
            I => \N__7887\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__7900\,
            I => \N__7884\
        );

    \I__1044\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7875\
        );

    \I__1043\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7875\
        );

    \I__1042\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7875\
        );

    \I__1041\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7875\
        );

    \I__1040\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7872\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__7890\,
            I => \beamXZ0Z_0\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__7887\,
            I => \beamXZ0Z_0\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__7884\,
            I => \beamXZ0Z_0\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__7875\,
            I => \beamXZ0Z_0\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__7872\,
            I => \beamXZ0Z_0\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__7861\,
            I => \N__7858\
        );

    \I__1033\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__7852\,
            I => \N_35\
        );

    \I__1030\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__7843\,
            I => \N_58_mux\
        );

    \I__1027\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7834\
        );

    \I__1026\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7831\
        );

    \I__1025\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7826\
        );

    \I__1024\ : InMux
    port map (
            O => \N__7837\,
            I => \N__7826\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__7834\,
            I => \N__7816\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__7831\,
            I => \N__7816\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7809\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__7825\,
            I => \N__7805\
        );

    \I__1019\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7800\
        );

    \I__1018\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7800\
        );

    \I__1017\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7795\
        );

    \I__1016\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7795\
        );

    \I__1015\ : Span4Mux_s3_v
    port map (
            O => \N__7816\,
            I => \N__7792\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7783\
        );

    \I__1013\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7783\
        );

    \I__1012\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7783\
        );

    \I__1011\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7783\
        );

    \I__1010\ : Span4Mux_h
    port map (
            O => \N__7809\,
            I => \N__7780\
        );

    \I__1009\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7775\
        );

    \I__1008\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7775\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__7800\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__7795\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__7792\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__7783\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__7780\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__7775\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__7762\,
            I => \beamY_RNIDQG2Z0Z_0_cascade_\
        );

    \I__1000\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7753\
        );

    \I__999\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7748\
        );

    \I__998\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7748\
        );

    \I__997\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7742\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7734\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__7748\,
            I => \N__7731\
        );

    \I__994\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7724\
        );

    \I__993\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7724\
        );

    \I__992\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7724\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7721\
        );

    \I__990\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7714\
        );

    \I__989\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7714\
        );

    \I__988\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7714\
        );

    \I__987\ : InMux
    port map (
            O => \N__7738\,
            I => \N__7709\
        );

    \I__986\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7709\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__7734\,
            I => \N__7706\
        );

    \I__984\ : Span4Mux_h
    port map (
            O => \N__7731\,
            I => \N__7703\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__7724\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__7721\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__7714\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__7709\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__7706\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__7703\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__977\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7687\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__7684\,
            I => \beamY_RNINKIU27Z0Z_0\
        );

    \I__974\ : InMux
    port map (
            O => \N__7681\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__7678\,
            I => \g2_1_cascade_\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__7675\,
            I => \N_7_cascade_\
        );

    \I__971\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__7669\,
            I => g2_1
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__7666\,
            I => \g0_1_0_cascade_\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__7663\,
            I => \g0_1_3_cascade_\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__7660\,
            I => \g3_2_2_cascade_\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__965\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__7651\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\
        );

    \I__963\ : InMux
    port map (
            O => \N__7648\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__962\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__7642\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\
        );

    \I__960\ : InMux
    port map (
            O => \N__7639\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__7636\,
            I => \N__7633\
        );

    \I__958\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__7630\,
            I => un5_visiblex_i_24
        );

    \I__956\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7624\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__7624\,
            I => charx_if_generate_plus_mult1_un26_sum_i_5
        );

    \I__954\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7615\
        );

    \I__953\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7615\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__7615\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__951\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7603\
        );

    \I__950\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7603\
        );

    \I__949\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7603\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__7603\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__947\ : InMux
    port map (
            O => \N__7600\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__946\ : InMux
    port map (
            O => \N__7597\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__945\ : InMux
    port map (
            O => \N__7594\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__944\ : InMux
    port map (
            O => \N__7591\,
            I => un8_beamx_cry_9
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__942\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__941\ : InMux
    port map (
            O => \N__7584\,
            I => \N__7575\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__7583\,
            I => \N__7571\
        );

    \I__939\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7568\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7565\
        );

    \I__937\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7562\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7559\
        );

    \I__935\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7555\
        );

    \I__934\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7552\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7549\
        );

    \I__932\ : Span4Mux_h
    port map (
            O => \N__7565\,
            I => \N__7542\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__7562\,
            I => \N__7542\
        );

    \I__930\ : Span4Mux_s1_h
    port map (
            O => \N__7559\,
            I => \N__7542\
        );

    \I__929\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7539\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__7555\,
            I => \beamXZ0Z_4\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7552\,
            I => \beamXZ0Z_4\
        );

    \I__926\ : Odrv12
    port map (
            O => \N__7549\,
            I => \beamXZ0Z_4\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__7542\,
            I => \beamXZ0Z_4\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7539\,
            I => \beamXZ0Z_4\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__922\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7518\
        );

    \I__921\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7514\
        );

    \I__920\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7511\
        );

    \I__919\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7508\
        );

    \I__918\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7505\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__7518\,
            I => \N__7502\
        );

    \I__916\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7498\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7514\,
            I => \N__7491\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7491\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__7508\,
            I => \N__7491\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7486\
        );

    \I__911\ : Span12Mux_s9_v
    port map (
            O => \N__7502\,
            I => \N__7486\
        );

    \I__910\ : InMux
    port map (
            O => \N__7501\,
            I => \N__7483\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__7498\,
            I => \beamXZ0Z_6\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__7491\,
            I => \beamXZ0Z_6\
        );

    \I__907\ : Odrv12
    port map (
            O => \N__7486\,
            I => \beamXZ0Z_6\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__7483\,
            I => \beamXZ0Z_6\
        );

    \I__905\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__7471\,
            I => un3_beamx_5
        );

    \I__903\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__7462\,
            I => un3_beamx_7
        );

    \I__900\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7453\
        );

    \I__899\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7448\
        );

    \I__898\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7448\
        );

    \I__897\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7445\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__7453\,
            I => \beamXZ0Z_2\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7448\,
            I => \beamXZ0Z_2\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__7445\,
            I => \beamXZ0Z_2\
        );

    \I__893\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__7437\,
            I => \N__7429\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__7436\,
            I => \N__7426\
        );

    \I__890\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7422\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7419\
        );

    \I__888\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7416\
        );

    \I__887\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7413\
        );

    \I__886\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7410\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7422\,
            I => \beamXZ0Z_3\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__7419\,
            I => \beamXZ0Z_3\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__7416\,
            I => \beamXZ0Z_3\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__7413\,
            I => \beamXZ0Z_3\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7410\,
            I => \beamXZ0Z_3\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__7399\,
            I => \N__7395\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__7398\,
            I => \N__7392\
        );

    \I__878\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7388\
        );

    \I__877\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7385\
        );

    \I__876\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7382\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__7388\,
            I => \N__7375\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__7385\,
            I => \N__7375\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7375\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__7375\,
            I => \N__7372\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__7372\,
            I => un18_beamylt4
        );

    \I__870\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7362\
        );

    \I__869\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7355\
        );

    \I__868\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7355\
        );

    \I__867\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7355\
        );

    \I__866\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7352\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__7362\,
            I => \beamXZ0Z_1\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__7355\,
            I => \beamXZ0Z_1\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__7352\,
            I => \beamXZ0Z_1\
        );

    \I__862\ : InMux
    port map (
            O => \N__7345\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__860\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__7336\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\
        );

    \I__858\ : InMux
    port map (
            O => \N__7333\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__857\ : InMux
    port map (
            O => \N__7330\,
            I => un8_beamx_cry_1
        );

    \I__856\ : InMux
    port map (
            O => \N__7327\,
            I => un8_beamx_cry_2
        );

    \I__855\ : InMux
    port map (
            O => \N__7324\,
            I => un8_beamx_cry_3
        );

    \I__854\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7315\
        );

    \I__853\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7310\
        );

    \I__852\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7307\
        );

    \I__851\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7304\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__7315\,
            I => \N__7301\
        );

    \I__849\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7297\
        );

    \I__848\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7294\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7289\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__7307\,
            I => \N__7289\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__7304\,
            I => \N__7284\
        );

    \I__844\ : Span4Mux_s1_h
    port map (
            O => \N__7301\,
            I => \N__7284\
        );

    \I__843\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7281\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__7297\,
            I => \beamXZ0Z_5\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__7294\,
            I => \beamXZ0Z_5\
        );

    \I__840\ : Odrv12
    port map (
            O => \N__7289\,
            I => \beamXZ0Z_5\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__7284\,
            I => \beamXZ0Z_5\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__7281\,
            I => \beamXZ0Z_5\
        );

    \I__837\ : InMux
    port map (
            O => \N__7270\,
            I => un8_beamx_cry_4
        );

    \I__836\ : InMux
    port map (
            O => \N__7267\,
            I => un8_beamx_cry_5
        );

    \I__835\ : InMux
    port map (
            O => \N__7264\,
            I => un8_beamx_cry_6
        );

    \I__834\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7252\
        );

    \I__833\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7252\
        );

    \I__832\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7249\
        );

    \I__831\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7244\
        );

    \I__830\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7244\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__7252\,
            I => \N__7239\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__7249\,
            I => \N__7239\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__7244\,
            I => \N__7232\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__7239\,
            I => \N__7232\
        );

    \I__825\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7229\
        );

    \I__824\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7226\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__7232\,
            I => \N__7221\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7221\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__7226\,
            I => \beamXZ0Z_8\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__7221\,
            I => \beamXZ0Z_8\
        );

    \I__819\ : InMux
    port map (
            O => \N__7216\,
            I => un8_beamx_cry_7
        );

    \I__818\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7204\
        );

    \I__817\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7204\
        );

    \I__816\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7201\
        );

    \I__815\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7195\
        );

    \I__814\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7195\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7190\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__7201\,
            I => \N__7190\
        );

    \I__811\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7186\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7181\
        );

    \I__809\ : Sp12to4
    port map (
            O => \N__7190\,
            I => \N__7181\
        );

    \I__808\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7178\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__7186\,
            I => \beamXZ0Z_9\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__7181\,
            I => \beamXZ0Z_9\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__7178\,
            I => \beamXZ0Z_9\
        );

    \I__804\ : InMux
    port map (
            O => \N__7171\,
            I => \bfn_2_11_0_\
        );

    \I__803\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7162\
        );

    \I__802\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7162\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__7162\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__7159\,
            I => \N__7156\
        );

    \I__799\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__7153\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\
        );

    \I__797\ : InMux
    port map (
            O => \N__7150\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__795\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7141\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\
        );

    \I__793\ : InMux
    port map (
            O => \N__7138\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__792\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7132\,
            I => charx_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__790\ : InMux
    port map (
            O => \N__7129\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__789\ : InMux
    port map (
            O => \N__7126\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__788\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7119\
        );

    \I__787\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7116\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__7119\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__7116\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__7111\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7102\
        );

    \I__782\ : InMux
    port map (
            O => \N__7107\,
            I => \N__7102\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__7102\,
            I => charx_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__779\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__7093\,
            I => charx_if_generate_plus_mult1_un54_sum_i
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__7090\,
            I => \un13_beamylt7_0_cascade_\
        );

    \I__776\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7084\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__7081\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\
        );

    \I__773\ : InMux
    port map (
            O => \N__7078\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__771\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__7066\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\
        );

    \I__768\ : InMux
    port map (
            O => \N__7063\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__767\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__7054\,
            I => charx_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__764\ : InMux
    port map (
            O => \N__7051\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__763\ : InMux
    port map (
            O => \N__7048\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__761\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7035\
        );

    \I__760\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7035\
        );

    \I__759\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7032\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__7035\,
            I => \N__7029\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__7032\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__7029\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__754\ : InMux
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__7018\,
            I => charx_if_generate_plus_mult1_un61_sum_i
        );

    \I__752\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__7012\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \N__7004\
        );

    \I__749\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6999\
        );

    \I__748\ : InMux
    port map (
            O => \N__7007\,
            I => \N__6994\
        );

    \I__747\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6994\
        );

    \I__746\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6991\
        );

    \I__745\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6988\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__6999\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__6994\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__6991\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__6988\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__740\ : InMux
    port map (
            O => \N__6979\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__739\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6971\
        );

    \I__738\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6968\
        );

    \I__737\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6965\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__6971\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__6968\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__6965\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\
        );

    \I__733\ : InMux
    port map (
            O => \N__6958\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__732\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__731\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6949\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__6949\,
            I => charx_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__729\ : InMux
    port map (
            O => \N__6946\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__728\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6940\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__6940\,
            I => \N__6932\
        );

    \I__726\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6925\
        );

    \I__725\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6925\
        );

    \I__724\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6925\
        );

    \I__723\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6920\
        );

    \I__722\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6920\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__6932\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__6925\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__6920\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__717\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__6907\,
            I => charx_if_generate_plus_mult1_un68_sum_i
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__6904\,
            I => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\
        );

    \I__714\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__6898\,
            I => font_un126_pixel_5_a0_2
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__6895\,
            I => \G_19_i_a11_0_1_cascade_\
        );

    \I__711\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__6889\,
            I => \Pixel_RNOZ0Z_36\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \g1_1_0_0_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__6880\,
            I => g0_0
        );

    \I__706\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6873\
        );

    \I__705\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6870\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__6873\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__703\ : LocalMux
    port map (
            O => \N__6870\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__702\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6862\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__6862\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__6859\,
            I => \N__6855\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__6858\,
            I => \N__6852\
        );

    \I__698\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6847\
        );

    \I__697\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6847\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__6847\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\
        );

    \I__695\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6838\
        );

    \I__694\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6838\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__6838\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__6835\,
            I => \g3_3_cascade_\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__6832\,
            I => \g0_0_2_cascade_\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__6829\,
            I => \g0_3_cascade_\
        );

    \I__689\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6823\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N_21_0\
        );

    \I__687\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6817\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__6817\,
            I => \Pixel_RNOZ0Z_37\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__6814\,
            I => \font_un126_pixel_m_2_1_1_cascade_\
        );

    \I__684\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__6808\,
            I => \Pixel_RNOZ0Z_71\
        );

    \I__682\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6802\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__6802\,
            I => g0_0_1
        );

    \I__680\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6796\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__6796\,
            I => font_un3_pixel_29
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__6793\,
            I => \font_un126_pixel_m_2_1_cascade_\
        );

    \I__677\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__6787\,
            I => g2_2_0_1
        );

    \I__675\ : InMux
    port map (
            O => \N__6784\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__674\ : InMux
    port map (
            O => \N__6781\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__673\ : InMux
    port map (
            O => \N__6778\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__672\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__6772\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\
        );

    \I__670\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6766\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__6766\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3_i
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__6763\,
            I => \g1_2_cascade_\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__6760\,
            I => \g2_3_0_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6754\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__6754\,
            I => g2_2_0
        );

    \I__664\ : InMux
    port map (
            O => \N__6751\,
            I => un5_visiblex_cry_2
        );

    \I__663\ : InMux
    port map (
            O => \N__6748\,
            I => un5_visiblex_cry_3
        );

    \I__662\ : InMux
    port map (
            O => \N__6745\,
            I => un5_visiblex_cry_4
        );

    \I__661\ : InMux
    port map (
            O => \N__6742\,
            I => un5_visiblex_cry_5
        );

    \I__660\ : InMux
    port map (
            O => \N__6739\,
            I => un5_visiblex_cry_6
        );

    \I__659\ : InMux
    port map (
            O => \N__6736\,
            I => \bfn_1_12_0_\
        );

    \I__658\ : InMux
    port map (
            O => \N__6733\,
            I => un5_visiblex_cry_8
        );

    \I__657\ : InMux
    port map (
            O => \N__6730\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__6727\,
            I => \N__6724\
        );

    \I__655\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6721\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__6721\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__6718\,
            I => \N__6715\
        );

    \I__652\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__6712\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__650\ : InMux
    port map (
            O => \N__6709\,
            I => un5_visiblex_cry_0
        );

    \I__649\ : InMux
    port map (
            O => \N__6706\,
            I => un5_visiblex_cry_1
        );

    \I__648\ : InMux
    port map (
            O => \N__6703\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__647\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6695\
        );

    \I__646\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6692\
        );

    \I__645\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6689\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__6695\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6692\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__6689\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__6682\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_\
        );

    \I__640\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__6676\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__638\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6667\
        );

    \I__637\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6667\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__6667\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__634\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6658\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\
        );

    \I__632\ : InMux
    port map (
            O => \N__6655\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__630\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__6646\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\
        );

    \I__628\ : InMux
    port map (
            O => \N__6643\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__627\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__6637\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__625\ : InMux
    port map (
            O => \N__6634\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__624\ : InMux
    port map (
            O => \N__6631\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__623\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6623\
        );

    \I__622\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6618\
        );

    \I__621\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6618\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__6623\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__6618\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\
        );

    \I__618\ : InMux
    port map (
            O => \N__6613\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__617\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__6607\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\
        );

    \I__615\ : InMux
    port map (
            O => \N__6604\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__613\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6595\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__6592\,
            I => un18_beamylto9_2
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__609\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__6583\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__606\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6574\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\
        );

    \I__604\ : InMux
    port map (
            O => \N__6571\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__602\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__6562\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\
        );

    \I__600\ : InMux
    port map (
            O => \N__6559\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__599\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__6553\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__597\ : InMux
    port map (
            O => \N__6550\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__596\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__6544\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\
        );

    \I__594\ : InMux
    port map (
            O => \N__6541\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__592\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6532\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__6532\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3\
        );

    \I__590\ : InMux
    port map (
            O => \N__6529\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__588\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__6520\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\
        );

    \I__586\ : InMux
    port map (
            O => \N__6517\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3
        );

    \I__585\ : InMux
    port map (
            O => \N__6514\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__583\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__582\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6502\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__6502\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\
        );

    \I__580\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6496\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__6496\,
            I => charx_i_24
        );

    \I__578\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__6490\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3\
        );

    \I__576\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__6484\,
            I => charx_i_23
        );

    \I__574\ : InMux
    port map (
            O => \N__6481\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__573\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__6475\,
            I => g1
        );

    \I__571\ : InMux
    port map (
            O => \N__6472\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1
        );

    \I__570\ : InMux
    port map (
            O => \N__6469\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2
        );

    \I__569\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__6463\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5
        );

    \I__567\ : InMux
    port map (
            O => \N__6460\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__6457\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__6454\,
            I => \N__6450\
        );

    \I__564\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6442\
        );

    \I__563\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6442\
        );

    \I__562\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6442\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__6442\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__6439\,
            I => \font_un3_pixel_29_cascade_\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__6436\,
            I => \Pixel_RNOZ0Z_18_cascade_\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__6433\,
            I => \N_1214_0_cascade_\
        );

    \I__557\ : IoInMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__6427\,
            I => \N__6424\
        );

    \I__555\ : Span4Mux_s1_h
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__553\ : Sp12to4
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__6415\,
            I => \Clock50MHz.PixelClock\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_9_8_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6430\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \beamX_RNII5M_9_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7259\,
            in1 => \N__8434\,
            in2 => \N__7528\,
            in3 => \N__7211\,
            lcout => un18_beamylto9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_0_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__7821\,
            in1 => \N__9296\,
            in2 => \_gnd_net_\,
            in3 => \N__7737\,
            lcout => font_un3_pixel_29,
            ltout => \font_un3_pixel_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_18_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9513\,
            in2 => \N__6439\,
            in3 => \N__9529\,
            lcout => OPEN,
            ltout => \Pixel_RNOZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_5_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__13108\,
            in1 => \N__6478\,
            in2 => \N__6436\,
            in3 => \N__8998\,
            lcout => OPEN,
            ltout => \N_1214_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_0_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__6826\,
            in1 => \N__6757\,
            in2 => \N__6433\,
            in3 => \N__6883\,
            lcout => \G_21_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_20_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110100101"
        )
    port map (
            in0 => \N__7738\,
            in1 => \_gnd_net_\,
            in2 => \N__9315\,
            in3 => \N__7822\,
            lcout => g1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7825\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6487\,
            in2 => \N__6511\,
            in3 => \N__6472\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_71_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6547\,
            in2 => \N__6454\,
            in3 => \N__6469\,
            lcout => \Pixel_RNOZ0Z_71\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_inv_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6466\,
            in2 => \N__6538\,
            in3 => \N__6449\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_i_5,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6453\,
            in1 => \N__6877\,
            in2 => \N__6526\,
            in3 => \N__6460\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\,
            ltout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_30_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7808\,
            in2 => \N__6457\,
            in3 => \N__7939\,
            lcout => g0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6507\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7015\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6499\,
            in2 => \_gnd_net_\,
            in3 => \N__6541\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDB3_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6493\,
            in2 => \N__15585\,
            in3 => \N__6529\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2_c_RNI21CDBZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6876\,
            in2 => \_gnd_net_\,
            in3 => \N__6517\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6514\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011000110011"
        )
    port map (
            in0 => \N__7003\,
            in1 => \N__6974\,
            in2 => \N__10342\,
            in3 => \N__6937\,
            lcout => charx_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101001110101"
        )
    port map (
            in0 => \N__6938\,
            in1 => \N__10330\,
            in2 => \N__7009\,
            in3 => \N__6975\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDABZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7007\,
            in2 => \N__10343\,
            in3 => \N__6939\,
            lcout => charx_i_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9997\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6679\,
            in2 => \N__6589\,
            in3 => \N__6481\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6700\,
            in2 => \N__6580\,
            in3 => \N__6613\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6610\,
            in2 => \N__6568\,
            in3 => \N__6698\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6556\,
            in2 => \_gnd_net_\,
            in3 => \N__6604\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIVEM1_4_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__7391\,
            in1 => \N__7321\,
            in2 => \N__6601\,
            in3 => \N__7584\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_2_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9841\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9840\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6672\,
            in2 => \N__6718\,
            in3 => \N__6571\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6627\,
            in2 => \N__6664\,
            in3 => \N__6559\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6699\,
            in1 => \N__6673\,
            in2 => \N__6652\,
            in3 => \N__6550\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6640\,
            in2 => \_gnd_net_\,
            in3 => \N__6703\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\,
            ltout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6682\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6626\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8704\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7167\,
            in2 => \N__6727\,
            in3 => \N__6655\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8248\,
            in2 => \N__8293\,
            in3 => \N__6643\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6628\,
            in1 => \N__7168\,
            in2 => \N__8278\,
            in3 => \N__6634\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8263\,
            in2 => \_gnd_net_\,
            in3 => \N__6631\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8977\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8705\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8465\,
            in1 => \N__7468\,
            in2 => \N__8420\,
            in3 => \N__7314\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_3_l_ofx_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101010110101"
        )
    port map (
            in0 => \N__8961\,
            in1 => \N__8906\,
            in2 => \N__9133\,
            in3 => \N__8684\,
            lcout => if_generate_plus_mult1_un54_sum_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_l_ofx_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110111100"
        )
    port map (
            in0 => \N__9126\,
            in1 => \N__8691\,
            in2 => \N__8911\,
            in3 => \N__8963\,
            lcout => if_generate_plus_mult1_un54_sum_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_c5_i_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001111100111"
        )
    port map (
            in0 => \N__8962\,
            in1 => \N__8907\,
            in2 => \N__9134\,
            in3 => \N__8685\,
            lcout => \column_1_if_generate_plus_mult1_un47_sum_c5_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8683\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7893\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7365\,
            in2 => \_gnd_net_\,
            in3 => \N__6709\,
            lcout => charx_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7456\,
            in2 => \_gnd_net_\,
            in3 => \N__6706\,
            lcout => charx_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7425\,
            in2 => \N__15586\,
            in3 => \N__6751\,
            lcout => chessboardpixel_un152_pixel_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7558\,
            in2 => \_gnd_net_\,
            in3 => \N__6748\,
            lcout => charx_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7300\,
            in2 => \_gnd_net_\,
            in3 => \N__6745\,
            lcout => charx_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7501\,
            in2 => \N__15587\,
            in3 => \N__6742\,
            lcout => charx_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8390\,
            in2 => \_gnd_net_\,
            in3 => \N__6739\,
            lcout => charx_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7238\,
            in2 => \N__15596\,
            in3 => \N__6736\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7189\,
            in2 => \_gnd_net_\,
            in3 => \N__6733\,
            lcout => charx_if_generate_plus_mult1_un26_sum_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8878\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6769\,
            in2 => \_gnd_net_\,
            in3 => \N__6730\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6775\,
            in2 => \N__15597\,
            in3 => \N__6784\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9100\,
            in2 => \_gnd_net_\,
            in3 => \N__6781\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6778\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_2_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9098\,
            lcout => charx_if_generate_plus_mult1_un26_sum_axb_3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_48_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__7212\,
            in1 => \N__7260\,
            in2 => \N__8440\,
            in3 => \N__8143\,
            lcout => OPEN,
            ltout => \g1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_26_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__8101\,
            in1 => \N__8338\,
            in2 => \N__6763\,
            in3 => \N__8191\,
            lcout => OPEN,
            ltout => \g2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_7_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6790\,
            in2 => \N__6760\,
            in3 => \N__7962\,
            lcout => g2_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_73_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__8435\,
            in1 => \N__8142\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \g3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_56_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__7261\,
            in1 => \N__8100\,
            in2 => \N__6835\,
            in3 => \N__7213\,
            lcout => g0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_38_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__7813\,
            in1 => \N__7961\,
            in2 => \_gnd_net_\,
            in3 => \N__7739\,
            lcout => OPEN,
            ltout => \g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_17_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6892\,
            in1 => \N__8155\,
            in2 => \N__6832\,
            in3 => \N__6820\,
            lcout => OPEN,
            ltout => \g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_4_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__6901\,
            in1 => \N__9016\,
            in2 => \N__6829\,
            in3 => \N__9007\,
            lcout => \N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_37_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__9295\,
            in1 => \N__13106\,
            in2 => \N__13294\,
            in3 => \N__9512\,
            lcout => \Pixel_RNOZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_72_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__9294\,
            in2 => \_gnd_net_\,
            in3 => \N__7960\,
            lcout => OPEN,
            ltout => \font_un126_pixel_m_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_55_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000110"
        )
    port map (
            in0 => \N__7740\,
            in1 => \N__7814\,
            in2 => \N__6814\,
            in3 => \N__6811\,
            lcout => OPEN,
            ltout => \font_un126_pixel_m_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_33_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__6805\,
            in1 => \N__6799\,
            in2 => \N__6793\,
            in3 => \N__8334\,
            lcout => g0_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_25_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010001100010"
        )
    port map (
            in0 => \N__7741\,
            in1 => \N__7815\,
            in2 => \N__12952\,
            in3 => \N__9308\,
            lcout => g2_2_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10341\,
            in2 => \_gnd_net_\,
            in3 => \N__6943\,
            lcout => charx_if_generate_plus_mult1_un1_sum_axb1,
            ltout => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_16_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000110001"
        )
    port map (
            in0 => \N__7745\,
            in1 => \N__9199\,
            in2 => \N__6904\,
            in3 => \N__9305\,
            lcout => font_un126_pixel_5_a0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_8_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7948\,
            in1 => \N__7824\,
            in2 => \_gnd_net_\,
            in3 => \N__7747\,
            lcout => OPEN,
            ltout => \G_19_i_a11_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__9337\,
            in1 => \N__9307\,
            in2 => \N__6895\,
            in3 => \N__9208\,
            lcout => \N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_36_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9198\,
            in1 => \N__13107\,
            in2 => \_gnd_net_\,
            in3 => \N__13287\,
            lcout => \Pixel_RNOZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_24_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001000000"
        )
    port map (
            in0 => \N__9306\,
            in1 => \N__7823\,
            in2 => \N__7861\,
            in3 => \N__7746\,
            lcout => OPEN,
            ltout => \g1_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_6_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__9367\,
            in1 => \N__9544\,
            in2 => \N__6886\,
            in3 => \N__8071\,
            lcout => g0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__7008\,
            in1 => \N__6976\,
            in2 => \N__10345\,
            in3 => \N__6936\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIL5OEN1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001111001100"
        )
    port map (
            in0 => \N__10005\,
            in1 => \N__6865\,
            in2 => \N__6858\,
            in3 => \N__6843\,
            lcout => chessboardpixel_un152_pixel_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAKPE41_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010011010000"
        )
    port map (
            in0 => \N__10006\,
            in1 => \N__10592\,
            in2 => \N__6859\,
            in3 => \N__6844\,
            lcout => chessboardpixel_un174_pixellt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__10337\,
            in1 => \N__7002\,
            in2 => \_gnd_net_\,
            in3 => \N__6935\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI8P51_4_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__7522\,
            in1 => \N__7319\,
            in2 => \N__7398\,
            in3 => \N__7582\,
            lcout => un13_beamylt7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10326\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6954\,
            in2 => \N__6913\,
            in3 => \N__6979\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7087\,
            in2 => \N__7045\,
            in3 => \N__6958\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6955\,
            in2 => \N__7075\,
            in3 => \N__7041\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7060\,
            in2 => \_gnd_net_\,
            in3 => \N__6946\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_RNO_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7320\,
            in1 => \N__7438\,
            in2 => \N__7588\,
            in3 => \N__7524\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10223\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7209\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_77_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__7523\,
            in1 => \N__7318\,
            in2 => \N__7399\,
            in3 => \N__7578\,
            lcout => OPEN,
            ltout => \un13_beamylt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_61_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__7210\,
            in1 => \N__7258\,
            in2 => \N__7090\,
            in3 => \N__8429\,
            lcout => g1_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10214\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7107\,
            in2 => \N__7024\,
            in3 => \N__7078\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7123\,
            in2 => \N__7159\,
            in3 => \N__7063\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7040\,
            in1 => \N__7108\,
            in2 => \N__7147\,
            in3 => \N__7051\,
            lcout => charx_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7135\,
            in2 => \_gnd_net_\,
            in3 => \N__7048\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10585\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8243\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8541\,
            in2 => \N__7099\,
            in3 => \N__7150\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9586\,
            in2 => \N__9631\,
            in3 => \N__7138\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7122\,
            in1 => \N__8542\,
            in2 => \N__9616\,
            in3 => \N__7129\,
            lcout => charx_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9601\,
            in2 => \_gnd_net_\,
            in3 => \N__7126\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\,
            ltout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7111\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10004\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7369\,
            in2 => \N__7930\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7459\,
            in2 => \_gnd_net_\,
            in3 => \N__7330\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7435\,
            in2 => \_gnd_net_\,
            in3 => \N__7327\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13360\,
            in1 => \N__7574\,
            in2 => \_gnd_net_\,
            in3 => \N__7324\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7313\,
            in2 => \_gnd_net_\,
            in3 => \N__7270\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7521\,
            in2 => \_gnd_net_\,
            in3 => \N__7267\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8405\,
            in2 => \_gnd_net_\,
            in3 => \N__7264\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7237\,
            in2 => \_gnd_net_\,
            in3 => \N__7216\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__13418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7200\,
            in2 => \_gnd_net_\,
            in3 => \N__7171\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__13419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13373\,
            in1 => \N__8487\,
            in2 => \_gnd_net_\,
            in3 => \N__7591\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_10_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7367\,
            in1 => \N__7458\,
            in2 => \N__7583\,
            in3 => \N__8486\,
            lcout => un3_beamx_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13374\,
            in2 => \_gnd_net_\,
            in3 => \N__7899\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_3_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7895\,
            in1 => \N__7517\,
            in2 => \N__7437\,
            in3 => \N__7474\,
            lcout => un3_beamx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__7457\,
            in1 => \N__7366\,
            in2 => \N__7436\,
            in3 => \N__7894\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7368\,
            in1 => \_gnd_net_\,
            in2 => \N__7913\,
            in3 => \_gnd_net_\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_1_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8967\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7621\,
            in2 => \N__7636\,
            in3 => \N__7345\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7611\,
            in2 => \N__7342\,
            in3 => \N__7333\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9164\,
            in1 => \N__7627\,
            in2 => \N__7657\,
            in3 => \N__7648\,
            lcout => charx_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7645\,
            in1 => \N__7612\,
            in2 => \N__9119\,
            in3 => \N__7639\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8879\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7610\,
            lcout => charx_if_generate_plus_mult1_un26_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7620\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9104\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15602\,
            in2 => \_gnd_net_\,
            in3 => \N__7600\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15606\,
            in2 => \N__15607\,
            in3 => \N__7597\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7594\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7681\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__7837\,
            in1 => \N__9319\,
            in2 => \_gnd_net_\,
            in3 => \N__7757\,
            lcout => g2_1,
            ltout => \g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_74_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13109\,
            in2 => \N__7678\,
            in3 => \N__13289\,
            lcout => OPEN,
            ltout => \N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_58_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__7838\,
            in1 => \N__7965\,
            in2 => \N__7675\,
            in3 => \N__7758\,
            lcout => g1_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_76_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__13290\,
            in1 => \_gnd_net_\,
            in2 => \N__13114\,
            in3 => \N__7964\,
            lcout => OPEN,
            ltout => \g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_60_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7672\,
            in1 => \N__7989\,
            in2 => \N__7666\,
            in3 => \N__9511\,
            lcout => OPEN,
            ltout => \g0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_35_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__12911\,
            in1 => \N__9922\,
            in2 => \N__7663\,
            in3 => \N__9909\,
            lcout => g3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_13_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__7966\,
            in1 => \N__13113\,
            in2 => \N__13296\,
            in3 => \N__7990\,
            lcout => OPEN,
            ltout => \g3_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_3_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__9244\,
            in1 => \N__8218\,
            in2 => \N__7660\,
            in3 => \N__7996\,
            lcout => OPEN,
            ltout => \g0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__7849\,
            in1 => \N__8059\,
            in2 => \N__8047\,
            in3 => \N__8044\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_34_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010001000"
        )
    port map (
            in0 => \N__7690\,
            in1 => \N__8020\,
            in2 => \N__7978\,
            in3 => \N__9514\,
            lcout => OPEN,
            ltout => \g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_12_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9217\,
            in1 => \N__8014\,
            in2 => \N__8005\,
            in3 => \N__8002\,
            lcout => g0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI50PU65_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7839\,
            in2 => \_gnd_net_\,
            in3 => \N__7759\,
            lcout => g1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_57_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13090\,
            lcout => g0_0_a3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_46_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__8326\,
            in1 => \N__8183\,
            in2 => \N__7963\,
            in3 => \N__8121\,
            lcout => \N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_2_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8184\,
            in1 => \N__8122\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \N_58_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDQG2_0_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13089\,
            lcout => OPEN,
            ltout => \beamY_RNIDQG2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNINKIU27_0_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__7840\,
            in1 => \N__9316\,
            in2 => \N__7762\,
            in3 => \N__7756\,
            lcout => \beamY_RNINKIU27Z0Z_0\,
            ltout => \beamY_RNINKIU27Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_29_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110101101"
        )
    port map (
            in0 => \N__9508\,
            in1 => \N__13091\,
            in2 => \N__8224\,
            in3 => \N__13297\,
            lcout => OPEN,
            ltout => \Pixel_RNOZ0Z_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_10_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__9231\,
            in1 => \N__9317\,
            in2 => \N__8221\,
            in3 => \N__9509\,
            lcout => \N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGH4H57_1_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110110"
        )
    port map (
            in0 => \N__8212\,
            in1 => \N__10939\,
            in2 => \N__8203\,
            in3 => \N__10852\,
            lcout => chessboardpixel_un175_pixel,
            ltout => \chessboardpixel_un175_pixel_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_39_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__8170\,
            in1 => \N__8088\,
            in2 => \N__8158\,
            in3 => \N__8325\,
            lcout => g2_3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNISO4T_7_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__8141\,
            in1 => \N__8087\,
            in2 => \N__8470\,
            in3 => \N__8430\,
            lcout => un15_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIT9ER_10_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8110\,
            in1 => \N__9352\,
            in2 => \N__8500\,
            in3 => \N__9412\,
            lcout => un15_beamy_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_44_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__9188\,
            in1 => \N__12910\,
            in2 => \N__9910\,
            in3 => \N__9467\,
            lcout => OPEN,
            ltout => \Pixel_RNOZ0Z_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_21_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000110"
        )
    port map (
            in0 => \N__13257\,
            in1 => \N__13093\,
            in2 => \N__8074\,
            in3 => \N__9346\,
            lcout => \N_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_45_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__13256\,
            in1 => \_gnd_net_\,
            in2 => \N__12931\,
            in3 => \_gnd_net_\,
            lcout => g4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSyncZ0_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__8499\,
            in1 => \N__8469\,
            in2 => \N__8439\,
            in3 => \N__8362\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI627QC51_6_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10921\,
            in1 => \N__8509\,
            in2 => \N__9421\,
            in3 => \N__9637\,
            lcout => un4_row,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8983\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8520\,
            in2 => \N__8740\,
            in3 => \N__8281\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8770\,
            in2 => \N__8857\,
            in3 => \N__8266\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8244\,
            in1 => \N__8521\,
            in2 => \N__8827\,
            in3 => \N__8254\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8797\,
            in2 => \_gnd_net_\,
            in3 => \N__8251\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9846\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8726\,
            in2 => \N__8530\,
            in3 => \N__8596\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8593\,
            in2 => \N__8581\,
            in3 => \N__8566\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9950\,
            in1 => \N__8727\,
            in2 => \N__8563\,
            in3 => \N__8548\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_LUT4_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8545\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9581\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_2_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8706\,
            lcout => un5_visiblex_i_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8766\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIOHGI2_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8746\,
            in1 => \N__8728\,
            in2 => \_gnd_net_\,
            in3 => \N__9952\,
            lcout => OPEN,
            ltout => \un4_row_9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNI1GN17_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11374\,
            in1 => \N__10864\,
            in2 => \N__8512\,
            in3 => \N__10899\,
            lcout => un4_row_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_s_5_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9657\,
            lcout => if_generate_plus_mult1_un54_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIK2PQ_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__8979\,
            in1 => \N__8905\,
            in2 => \N__11386\,
            in3 => \N__9136\,
            lcout => un4_row_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_c5_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000111001000"
        )
    port map (
            in0 => \N__8978\,
            in1 => \N__8903\,
            in2 => \N__8713\,
            in3 => \N__9135\,
            lcout => \column_1_if_generate_plus_mult1_un47_sum_cZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8697\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9144\,
            in2 => \N__8920\,
            in3 => \N__8650\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9172\,
            in2 => \N__8647\,
            in3 => \N__8632\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9768\,
            in1 => \N__9145\,
            in2 => \N__8629\,
            in3 => \N__8614\,
            lcout => charx_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8611\,
            in2 => \_gnd_net_\,
            in3 => \N__8599\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\,
            ltout => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8986\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8968\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9839\,
            lcout => un5_visiblex_i_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8902\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9024\,
            in2 => \N__9061\,
            in3 => \N__8845\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9039\,
            in2 => \N__8842\,
            in3 => \N__8815\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8765\,
            in1 => \N__9025\,
            in2 => \N__8812\,
            in3 => \N__8788\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__8785\,
            in1 => \N__9040\,
            in2 => \_gnd_net_\,
            in3 => \N__8773\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9168\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9132\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15600\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9052\,
            in2 => \_gnd_net_\,
            in3 => \N__9043\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9038\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_14_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000010"
        )
    port map (
            in0 => \N__13092\,
            in1 => \N__9887\,
            in2 => \N__13295\,
            in3 => \N__12913\,
            lcout => \Pixel_RNOZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_15_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__12912\,
            in1 => \N__13283\,
            in2 => \N__9901\,
            in3 => \N__9510\,
            lcout => font_un126_pixel_5_a0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_19_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__9853\,
            in1 => \N__10132\,
            in2 => \N__13288\,
            in3 => \N__9504\,
            lcout => \N_1740_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_54_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100001000010"
        )
    port map (
            in0 => \N__11181\,
            in1 => \N__10125\,
            in2 => \N__12673\,
            in3 => \N__12917\,
            lcout => font_un28_pixel_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM1QKG9_0_3_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000100100"
        )
    port map (
            in0 => \N__10124\,
            in1 => \N__12665\,
            in2 => \N__12932\,
            in3 => \N__11180\,
            lcout => font_un28_pixel_29,
            ltout => \font_un28_pixel_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDA2GGA3_0_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101101100"
        )
    port map (
            in0 => \N__9503\,
            in1 => \N__13099\,
            in2 => \N__9340\,
            in3 => \N__13262\,
            lcout => \beamY_RNIDA2GGA3Z0Z_0\,
            ltout => \beamY_RNIDA2GGA3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_11_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__9328\,
            in1 => \N__9318\,
            in2 => \N__9247\,
            in3 => \N__9379\,
            lcout => \N_19_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_32_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__9238\,
            in1 => \N__13263\,
            in2 => \_gnd_net_\,
            in3 => \N__9232\,
            lcout => \N_15_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_28_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101100010100"
        )
    port map (
            in0 => \N__9192\,
            in1 => \N__12918\,
            in2 => \N__9902\,
            in3 => \N__9502\,
            lcout => OPEN,
            ltout => \Pixel_RNOZ0Z_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_9_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__13276\,
            in1 => \N__13100\,
            in2 => \N__9211\,
            in3 => \N__9397\,
            lcout => \Pixel_RNOZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_52_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__12644\,
            in1 => \N__9894\,
            in2 => \N__12933\,
            in3 => \N__10090\,
            lcout => g1_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM1QKG9_3_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010011001"
        )
    port map (
            in0 => \N__10117\,
            in1 => \N__12643\,
            in2 => \N__11182\,
            in3 => \N__12921\,
            lcout => chary_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_50_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110000111001"
        )
    port map (
            in0 => \N__12922\,
            in1 => \N__12648\,
            in2 => \N__10765\,
            in3 => \N__10119\,
            lcout => OPEN,
            ltout => \chary_1_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_27_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011101"
        )
    port map (
            in0 => \N__11827\,
            in1 => \N__10081\,
            in2 => \N__9400\,
            in3 => \N__9491\,
            lcout => \N_1737_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_70_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000101101"
        )
    port map (
            in0 => \N__12926\,
            in1 => \N__10663\,
            in2 => \N__12670\,
            in3 => \N__10118\,
            lcout => OPEN,
            ltout => \chary_1_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_53_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110011001"
        )
    port map (
            in0 => \N__13264\,
            in1 => \N__13056\,
            in2 => \N__9391\,
            in3 => \N__10080\,
            lcout => OPEN,
            ltout => \g2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_31_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101100010"
        )
    port map (
            in0 => \N__9492\,
            in1 => \N__9373\,
            in2 => \N__9388\,
            in3 => \N__9385\,
            lcout => un116_pixel_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_51_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13055\,
            in2 => \_gnd_net_\,
            in3 => \N__13258\,
            lcout => \N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_22_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13481\,
            in1 => \N__12105\,
            in2 => \N__12671\,
            in3 => \N__12172\,
            lcout => g0_0_a3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_4_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__12456\,
            in1 => \N__12656\,
            in2 => \N__10840\,
            in3 => \N__12920\,
            lcout => OPEN,
            ltout => \un8_beamylto9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_0_9_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13480\,
            in1 => \N__12104\,
            in2 => \N__9355\,
            in3 => \N__12171\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_43_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__10057\,
            in1 => \N__10174\,
            in2 => \N__10159\,
            in3 => \N__9458\,
            lcout => \N_134_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_23_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__12457\,
            in1 => \N__12328\,
            in2 => \N__12253\,
            in3 => \N__9550\,
            lcout => g0_0_a3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_62_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__10420\,
            in1 => \N__13226\,
            in2 => \N__11692\,
            in3 => \N__10267\,
            lcout => OPEN,
            ltout => \m4_rn_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_40_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__10540\,
            in1 => \_gnd_net_\,
            in2 => \N__9532\,
            in3 => \N__9406\,
            lcout => \Pixel_RNOZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram0__RNIR1C2R81_0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001111111011"
        )
    port map (
            in0 => \N__10461\,
            in1 => \N__10265\,
            in2 => \N__11691\,
            in3 => \N__10539\,
            lcout => OPEN,
            ltout => \content_content_ram0__RNIR1C2R81Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram0__RNIAENOV03_0_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9643\,
            in2 => \N__9517\,
            in3 => \N__10419\,
            lcout => \N_331_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0H2_0_4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12455\,
            lcout => OPEN,
            ltout => \un4_row_m7_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPAQ91_6_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110000010"
        )
    port map (
            in0 => \N__10900\,
            in1 => \N__12324\,
            in2 => \N__9424\,
            in3 => \N__12243\,
            lcout => \beamY_RNIPAQ91Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISI4A_9_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__12102\,
            in1 => \N__13486\,
            in2 => \N__10144\,
            in3 => \N__12164\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_63_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10266\,
            in1 => \_gnd_net_\,
            in2 => \N__13265\,
            in3 => \N__10462\,
            lcout => m4_sn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram0__RNIR1C2R81_0_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001000"
        )
    port map (
            in0 => \N__10459\,
            in1 => \N__10253\,
            in2 => \N__11684\,
            in3 => \N__10538\,
            lcout => \content_content_ram0__RNIR1C2R81_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un6_rowlto3_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__11659\,
            in1 => \N__10460\,
            in2 => \N__10264\,
            in3 => \N__11597\,
            lcout => un6_rowlt7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10003\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9676\,
            in2 => \N__9565\,
            in3 => \N__9619\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9778\,
            in2 => \N__9697\,
            in3 => \N__9604\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9582\,
            in1 => \N__9556\,
            in2 => \N__9748\,
            in3 => \N__9592\,
            lcout => charx_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9715\,
            in2 => \_gnd_net_\,
            in3 => \N__9589\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9847\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__9747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9692\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9842\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9732\,
            in2 => \N__9790\,
            in3 => \N__9772\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9769\,
            in2 => \N__9757\,
            in3 => \N__9736\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9696\,
            in1 => \N__9733\,
            in2 => \N__9724\,
            in3 => \N__9709\,
            lcout => charx_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9706\,
            in2 => \_gnd_net_\,
            in3 => \N__9700\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\,
            ltout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9679\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9995\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9670\,
            in2 => \N__9664\,
            in3 => \N__9646\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9951\,
            in2 => \N__10051\,
            in3 => \N__10039\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11570\,
            in1 => \N__9928\,
            in2 => \N__10036\,
            in3 => \N__10024\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_s_5_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10021\,
            in2 => \_gnd_net_\,
            in3 => \N__10012\,
            lcout => if_generate_plus_mult1_un61_sum_s_5,
            ltout => \if_generate_plus_mult1_un61_sum_s_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10009\,
            in3 => \_gnd_net_\,
            lcout => column_1_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_i_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9996\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9949\,
            lcout => column_1_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_59_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110101001"
        )
    port map (
            in0 => \N__12664\,
            in1 => \N__12930\,
            in2 => \N__10126\,
            in3 => \N__10690\,
            lcout => chary_2_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI539IG9_3_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12018\,
            in1 => \N__11862\,
            in2 => \N__11128\,
            in3 => \N__11179\,
            lcout => \beamY_RNI539IG9Z0Z_3\,
            ltout => \beamY_RNI539IG9Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_42_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9856\,
            in3 => \N__12886\,
            lcout => g4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_41_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100001001011"
        )
    port map (
            in0 => \N__10063\,
            in1 => \N__12887\,
            in2 => \N__12672\,
            in3 => \N__10120\,
            lcout => chary_0_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6CM834_3_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11109\,
            in1 => \N__12003\,
            in2 => \_gnd_net_\,
            in3 => \N__11863\,
            lcout => chary_if_generate_plus_mult1_un75_sum_axbxc5_1,
            ltout => \chary_if_generate_plus_mult1_un75_sum_axbxc5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_69_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000001111"
        )
    port map (
            in0 => \N__15059\,
            in1 => \N__11938\,
            in2 => \N__10093\,
            in3 => \N__12888\,
            lcout => g1_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_78_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000101010"
        )
    port map (
            in0 => \N__14718\,
            in1 => \N__14974\,
            in2 => \N__10186\,
            in3 => \N__14278\,
            lcout => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMSO1N7_0_2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12004\,
            in1 => \N__11167\,
            in2 => \N__12934\,
            in3 => \N__11110\,
            lcout => OPEN,
            ltout => \beamY_RNIMSO1N7_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJEAL7H_2_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10672\,
            in2 => \N__10084\,
            in3 => \N__11864\,
            lcout => g4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_79_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100000000"
        )
    port map (
            in0 => \N__14279\,
            in1 => \N__10185\,
            in2 => \N__14985\,
            in3 => \N__10168\,
            lcout => OPEN,
            ltout => \g2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_64_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000110110"
        )
    port map (
            in0 => \N__10072\,
            in1 => \N__15058\,
            in2 => \N__10066\,
            in3 => \N__12005\,
            lcout => chary_if_generate_plus_mult1_un68_sum_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_66_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000001"
        )
    port map (
            in0 => \N__12654\,
            in1 => \N__12014\,
            in2 => \N__11127\,
            in3 => \N__11865\,
            lcout => \Pixel_RNOZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_2_4_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12460\,
            in1 => \N__12652\,
            in2 => \_gnd_net_\,
            in3 => \N__12878\,
            lcout => un5_visibley_0_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_65_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101001"
        )
    port map (
            in0 => \N__12880\,
            in1 => \N__10717\,
            in2 => \N__10741\,
            in3 => \N__15067\,
            lcout => g2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_87_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12653\,
            in2 => \_gnd_net_\,
            in3 => \N__12879\,
            lcout => un5_visibley_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_67_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__11866\,
            in1 => \N__11123\,
            in2 => \N__12019\,
            in3 => \N__12655\,
            lcout => \Pixel_RNOZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4H2_6_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12241\,
            lcout => un8_beamy_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_1_3_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12588\,
            in2 => \_gnd_net_\,
            in3 => \N__12838\,
            lcout => OPEN,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2KA6_6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12242\,
            in1 => \N__12441\,
            in2 => \N__10147\,
            in3 => \N__12323\,
            lcout => un4_beamylt8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__13391\,
            in1 => \N__13531\,
            in2 => \_gnd_net_\,
            in3 => \N__13026\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13421\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10344\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10278\,
            in2 => \N__10240\,
            in3 => \N__10445\,
            lcout => \G_383\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10448\,
            in2 => \N__10198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_4_c_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10279\,
            in2 => \N__10495\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_s_5_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10483\,
            in2 => \_gnd_net_\,
            in3 => \N__10270\,
            lcout => un6_rowlto0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_i_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10231\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10230\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10549\,
            in2 => \N__10471\,
            in3 => \N__10189\,
            lcout => if_generate_plus_mult1_un75_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11643\,
            in2 => \N__10396\,
            in3 => \N__10486\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10446\,
            in1 => \N__10614\,
            in2 => \N__10603\,
            in3 => \N__10477\,
            lcout => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_s_5_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10636\,
            in2 => \_gnd_net_\,
            in3 => \N__10474\,
            lcout => un6_rowlto1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_column_1_i_2_sbtinv_2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11641\,
            lcout => content_column_1_i_2_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram5__RNIKAVJ9F_0_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10447\,
            in1 => \_gnd_net_\,
            in2 => \N__11056\,
            in3 => \N__10510\,
            lcout => \content_N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10593\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10371\,
            in2 => \N__10405\,
            in3 => \N__10387\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11571\,
            in2 => \N__10384\,
            in3 => \N__10375\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11642\,
            in1 => \N__10372\,
            in2 => \N__10645\,
            in3 => \N__10630\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_s_5_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10627\,
            in2 => \_gnd_net_\,
            in3 => \N__10621\,
            lcout => content_column_1_i_2_2,
            ltout => \content_column_1_i_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10618\,
            in3 => \N__10615\,
            lcout => if_generate_plus_mult1_un75_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_i_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram8__e_0_RNI0I9HN1_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__11646\,
            in1 => \N__11574\,
            in2 => \N__11812\,
            in3 => \N__11365\,
            lcout => OPEN,
            ltout => \content_m7_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram0__RNIEAKG02_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__11575\,
            in1 => \N__11779\,
            in2 => \N__10543\,
            in3 => \N__11499\,
            lcout => \content_N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram11__e_0_RNIQ1Q3O1_0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__11573\,
            in1 => \N__11526\,
            in2 => \N__11035\,
            in3 => \N__11645\,
            lcout => OPEN,
            ltout => \content_content_ram11__e_0_RNIQ1Q3O1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram7__RNI6B0NG3_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11721\,
            in2 => \N__10513\,
            in3 => \N__10501\,
            lcout => \content_content_ram7__RNI6B0NG3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram11__e_0_RNIQ1Q3O1_0_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__11572\,
            in1 => \N__11644\,
            in2 => \N__11034\,
            in3 => \N__11525\,
            lcout => \content_content_ram11__e_0_RNIQ1Q3O1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_92_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12660\,
            in2 => \_gnd_net_\,
            in3 => \N__12881\,
            lcout => un5_visibley_2_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_85_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000101010"
        )
    port map (
            in0 => \N__14719\,
            in1 => \N__10992\,
            in2 => \N__14984\,
            in3 => \N__14281\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_75_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000110110"
        )
    port map (
            in0 => \N__10678\,
            in1 => \N__15063\,
            in2 => \N__10693\,
            in3 => \N__12002\,
            lcout => chary_if_generate_plus_mult1_un68_sum_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_86_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__10684\,
            in1 => \N__10993\,
            in2 => \N__14983\,
            in3 => \N__14282\,
            lcout => g2_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMSO1N7_2_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11994\,
            in1 => \N__11155\,
            in2 => \N__11119\,
            in3 => \N__12882\,
            lcout => \beamY_RNIMSO1N7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_82_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010011001100"
        )
    port map (
            in0 => \N__14277\,
            in1 => \N__14703\,
            in2 => \N__14986\,
            in3 => \N__10702\,
            lcout => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_91_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000101010"
        )
    port map (
            in0 => \N__14702\,
            in1 => \N__14982\,
            in2 => \N__11929\,
            in3 => \N__14275\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_84_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101111110100"
        )
    port map (
            in0 => \N__11993\,
            in1 => \N__10654\,
            in2 => \N__10666\,
            in3 => \N__15056\,
            lcout => chary_if_generate_plus_mult1_un68_sum_1_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6C1MV_3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__10701\,
            in1 => \N__14981\,
            in2 => \N__11137\,
            in3 => \N__14276\,
            lcout => g2_0,
            ltout => \g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_68_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001111011100"
        )
    port map (
            in0 => \N__11995\,
            in1 => \N__10774\,
            in2 => \N__10768\,
            in3 => \N__15057\,
            lcout => chary_if_generate_plus_mult1_un68_sum_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSyncZ0_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101110111"
        )
    port map (
            in0 => \N__11074\,
            in1 => \N__10711\,
            in2 => \N__12919\,
            in3 => \N__13251\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_80_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000101010"
        )
    port map (
            in0 => \N__14717\,
            in1 => \N__14949\,
            in2 => \N__10732\,
            in3 => \N__14284\,
            lcout => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_4_4_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12458\,
            in1 => \N__12649\,
            in2 => \_gnd_net_\,
            in3 => \N__12875\,
            lcout => un5_visibley_3_28,
            ltout => \un5_visibley_3_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_88_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14948\,
            in2 => \N__10723\,
            in3 => \N__14283\,
            lcout => OPEN,
            ltout => \g1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_81_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__11984\,
            in1 => \N__12651\,
            in2 => \N__10720\,
            in3 => \N__12877\,
            lcout => g2_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_RNO_1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10839\,
            in1 => \N__13485\,
            in2 => \_gnd_net_\,
            in3 => \N__12106\,
            lcout => un1_beamylto9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_1_4_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12459\,
            in1 => \N__12650\,
            in2 => \_gnd_net_\,
            in3 => \N__12876\,
            lcout => un5_visibley_1_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001010101010"
        )
    port map (
            in0 => \N__13156\,
            in1 => \N__13520\,
            in2 => \N__13074\,
            in3 => \N__13384\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI70BUG1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010001000"
        )
    port map (
            in0 => \N__10792\,
            in1 => \N__10950\,
            in2 => \N__10816\,
            in3 => \N__10974\,
            lcout => OPEN,
            ltout => \chessboardpixel_un200_pixellto4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQF0E52_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__10975\,
            in1 => \N__13155\,
            in2 => \N__10855\,
            in3 => \N__10814\,
            lcout => chessboardpixel_un200_pixellt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIID25_0_7_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__12103\,
            in1 => \N__10838\,
            in2 => \_gnd_net_\,
            in3 => \N__12165\,
            lcout => un5_beamx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12587\,
            in2 => \_gnd_net_\,
            in3 => \N__12806\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12807\,
            in1 => \N__15483\,
            in2 => \_gnd_net_\,
            in3 => \N__10815\,
            lcout => \beamY_i_2\,
            ltout => \beamY_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10819\,
            in3 => \N__10791\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10810\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQB_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10927\,
            in2 => \N__11328\,
            in3 => \N__10783\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIA5IQBZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLG_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11323\,
            in2 => \N__11212\,
            in3 => \N__10780\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI1PBLGZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777J_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11200\,
            in2 => \N__11329\,
            in3 => \N__10777\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG777JZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10984\,
            in2 => \N__11353\,
            in3 => \N__11319\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEK_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11341\,
            in2 => \_gnd_net_\,
            in3 => \N__10978\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0\,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIS1DEKZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIN7I542_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__10966\,
            in1 => \N__10960\,
            in2 => \N__10954\,
            in3 => \N__10951\,
            lcout => chessboardpixel_un178_pixel_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11229\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111000010111"
        )
    port map (
            in0 => \N__15190\,
            in1 => \N__15709\,
            in2 => \N__15295\,
            in3 => \N__15121\,
            lcout => if_generate_plus_mult1_un54_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_c5_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111110100"
        )
    port map (
            in0 => \N__10886\,
            in1 => \N__14791\,
            in2 => \N__10909\,
            in3 => \N__15290\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_axb3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__15191\,
            in1 => \N__15717\,
            in2 => \_gnd_net_\,
            in3 => \N__15122\,
            lcout => \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3\,
            ltout => \row_1_if_generate_plus_mult1_un54_sum_axbZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__14790\,
            in2 => \N__10867\,
            in3 => \N__15289\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram9__e_0_RNIFBHPN1_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__11652\,
            in1 => \N__11589\,
            in2 => \N__13726\,
            in3 => \N__11043\,
            lcout => \content_content_ram9__e_0_RNIFBHPN1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram9__e_0_RNIFBHPN1_0_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__11590\,
            in1 => \N__13725\,
            in2 => \N__11047\,
            in3 => \N__11653\,
            lcout => OPEN,
            ltout => \content_content_ram9__e_0_RNIFBHPN1_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram5__RNIEM2QF3_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11460\,
            in2 => \N__11065\,
            in3 => \N__11062\,
            lcout => \content_content_ram5__RNIEM2QF3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram9__e_0_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14539\,
            lcout => content_ram9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14339\,
            ce => \N__11506\,
            sr => \_gnd_net_\
        );

    \content_content_ram11__e_0_0_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => content_ram11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14340\,
            ce => \N__11470\,
            sr => \_gnd_net_\
        );

    \nCS1_1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011111100010101"
        )
    port map (
            in0 => \N__14436\,
            in1 => \N__14191\,
            in2 => \N__14581\,
            in3 => \N__11004\,
            lcout => \nCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14344\,
            ce => 'H',
            sr => \N__11701\
        );

    \beamY_RNIBFP3_3_4_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12858\,
            in1 => \N__12438\,
            in2 => \_gnd_net_\,
            in3 => \N__12600\,
            lcout => un5_visibley_2_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4QL4A1_4_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000011110000"
        )
    port map (
            in0 => \N__14266\,
            in1 => \N__14951\,
            in2 => \N__14715\,
            in3 => \N__14827\,
            lcout => chary_if_generate_plus_mult1_un68_sum_ac0_7_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPAS0A1_4_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14267\,
            in1 => \_gnd_net_\,
            in2 => \N__14716\,
            in3 => \N__14950\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6C1MV_1_3_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__14952\,
            in1 => \N__14828\,
            in2 => \N__11239\,
            in3 => \N__14265\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVMI9D5_3_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011010"
        )
    port map (
            in0 => \N__15052\,
            in1 => \N__11983\,
            in2 => \N__11191\,
            in3 => \N__11188\,
            lcout => \beamY_RNIVMI9D5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12636\,
            in2 => \_gnd_net_\,
            in3 => \N__12857\,
            lcout => un5_visibley_1_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6C1MV_0_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100000110"
        )
    port map (
            in0 => \N__14268\,
            in1 => \N__14953\,
            in2 => \N__14846\,
            in3 => \N__11238\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8325_6_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__12308\,
            in2 => \N__12586\,
            in3 => \N__12750\,
            lcout => OPEN,
            ltout => \beamY_RNI8325Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPOR8_6_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__12309\,
            in1 => \N__12406\,
            in2 => \N__11080\,
            in3 => \N__12228\,
            lcout => un5_visibley_c5,
            ltout => \un5_visibley_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJNLC_9_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110111010101"
        )
    port map (
            in0 => \N__13467\,
            in1 => \N__12080\,
            in2 => \N__11077\,
            in3 => \N__12152\,
            lcout => \beamY_RNIJNLCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_RNO_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12538\,
            in1 => \N__12433\,
            in2 => \_gnd_net_\,
            in3 => \N__12153\,
            lcout => un1_beamylto9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_4_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12394\,
            in1 => \N__12529\,
            in2 => \_gnd_net_\,
            in3 => \N__12742\,
            lcout => un5_visibley_c3,
            ltout => \un5_visibley_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV7J7_7_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__12149\,
            in1 => \N__12223\,
            in2 => \N__11068\,
            in3 => \N__12303\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8325_9_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13452\,
            in1 => \N__12531\,
            in2 => \N__12434\,
            in3 => \N__13101\,
            lcout => OPEN,
            ltout => \un5_beamx_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__12743\,
            in1 => \N__13197\,
            in2 => \N__11260\,
            in3 => \N__11257\,
            lcout => \beamY_RNI9DLCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8325_0_6_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110011001"
        )
    port map (
            in0 => \N__12304\,
            in1 => \N__12226\,
            in2 => \N__12805\,
            in3 => \N__12530\,
            lcout => \beamY_RNI8325_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIID25_7_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12148\,
            in1 => \N__12222\,
            in2 => \N__12093\,
            in3 => \N__12302\,
            lcout => OPEN,
            ltout => \un5_visibley_ac0_11_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ7DB_9_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010100101"
        )
    port map (
            in0 => \N__13451\,
            in1 => \N__12076\,
            in2 => \N__11251\,
            in3 => \N__11895\,
            lcout => chary_if_generate_plus_mult1_un33_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPOR8_0_6_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010110001"
        )
    port map (
            in0 => \N__12405\,
            in1 => \N__12224\,
            in2 => \N__11248\,
            in3 => \N__12305\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11228\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOU4_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11426\,
            in2 => \N__11302\,
            in3 => \N__11203\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNITAOUZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIG7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11293\,
            in2 => \N__11431\,
            in3 => \N__11194\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNIBNIGZ0Z7\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5V28_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11430\,
            in2 => \N__11284\,
            in3 => \N__11344\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNII5VZ0Z28\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8PPUJ_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11327\,
            in1 => \N__11407\,
            in2 => \N__11272\,
            in3 => \N__11335\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37B_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11443\,
            in2 => \_gnd_net_\,
            in3 => \N__11332\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIJB37BZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14847\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLM2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13591\,
            in2 => \N__11395\,
            in3 => \N__11287\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNIDMLMZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJ2193_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13594\,
            in2 => \N__13675\,
            in3 => \N__11275\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIJZ0Z2193\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NT3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13592\,
            in2 => \N__13654\,
            in3 => \N__11263\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIL8NTZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNITBNTA_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11425\,
            in1 => \N__11401\,
            in2 => \N__13636\,
            in3 => \N__11437\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13612\,
            in2 => \_gnd_net_\,
            in3 => \N__11434\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4\,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KGZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIB7KG4_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11410\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJ54_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13635\,
            in2 => \_gnd_net_\,
            in3 => \N__13590\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIMJZ0Z54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14769\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN49K_8_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15123\,
            in2 => \_gnd_net_\,
            in3 => \N__15188\,
            lcout => \CO4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un47_sum_c5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000001010"
        )
    port map (
            in0 => \N__15189\,
            in1 => \_gnd_net_\,
            in2 => \N__15127\,
            in3 => \N__15718\,
            lcout => \row_1_if_generate_plus_mult1_un47_sum_cZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram8__e_0_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14538\,
            lcout => content_ram8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14341\,
            ce => \N__11482\,
            sr => \_gnd_net_\
        );

    \content_content_ram10__e_0_RNIOLNMN1_0_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__11658\,
            in1 => \N__13828\,
            in2 => \N__11599\,
            in3 => \N__13797\,
            lcout => OPEN,
            ltout => \content_content_ram10__e_0_RNIOLNMN1_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram6__RNI1FLOF3_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11743\,
            in2 => \N__11695\,
            in3 => \N__11533\,
            lcout => \content_N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram10__e_0_RNIOLNMN1_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__11657\,
            in1 => \N__13827\,
            in2 => \N__11598\,
            in3 => \N__13796\,
            lcout => \content_content_ram10__e_0_RNIOLNMN1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram3__0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__14541\,
            in1 => \N__13807\,
            in2 => \N__11527\,
            in3 => \N__14047\,
            lcout => content_ram3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram9__e_0_RNO_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__13782\,
            in1 => \N__13757\,
            in2 => \N__13918\,
            in3 => \N__14173\,
            lcout => content_awe9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram0__0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__11788\,
            in1 => \N__13758\,
            in2 => \N__11500\,
            in3 => \N__14540\,
            lcout => content_ram0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram8__e_0_RNO_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13698\,
            in1 => \N__14045\,
            in2 => \N__13763\,
            in3 => \N__14111\,
            lcout => content_awe8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram11__e_0_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13697\,
            in1 => \N__14046\,
            in2 => \N__13764\,
            in3 => \N__14112\,
            lcout => content_awe11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram5__0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__11760\,
            in1 => \N__13783\,
            in2 => \N__11461\,
            in3 => \N__14537\,
            lcout => content_ram5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_0_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14608\,
            in2 => \_gnd_net_\,
            in3 => \N__14044\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__14116\,
            in1 => \N__14043\,
            in2 => \_gnd_net_\,
            in3 => \N__14609\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram12__0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__11761\,
            in1 => \N__13699\,
            in2 => \N__11808\,
            in3 => \N__14535\,
            lcout => content_ram12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNINMOJ_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__14171\,
            in1 => \N__14110\,
            in2 => \N__14059\,
            in3 => \N__13903\,
            lcout => content_awe0_0_a2_0,
            ltout => \content_awe0_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram4__0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__11759\,
            in1 => \N__14536\,
            in2 => \N__11782\,
            in3 => \N__11775\,
            lcout => content_ram4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIHRI6_1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14042\,
            in2 => \_gnd_net_\,
            in3 => \N__14109\,
            lcout => \content_N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIVRML1_2_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__13973\,
            in1 => \N__14433\,
            in2 => \N__14395\,
            in3 => \N__13955\,
            lcout => \content_N_36\,
            ltout => \content_N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIGN9S1_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14115\,
            in2 => \N__11749\,
            in3 => \N__14053\,
            lcout => content_awe7_1,
            ltout => \content_awe7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram6__0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14054\,
            in1 => \N__14530\,
            in2 => \N__11746\,
            in3 => \N__11742\,
            lcout => content_ram6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram7__0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__11728\,
            in2 => \N__11722\,
            in3 => \N__14055\,
            lcout => content_ram7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nCS1_1_RNO_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__14571\,
            in1 => \N__11880\,
            in2 => \_gnd_net_\,
            in3 => \N__14434\,
            lcout => \nCS1_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIICFG_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__13954\,
            in1 => \N__13851\,
            in2 => \N__13917\,
            in3 => \N__13974\,
            lcout => un19_slaveselectlt5_0,
            ltout => \un19_slaveselectlt5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI4HQB1_5_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101110111"
        )
    port map (
            in0 => \N__14572\,
            in1 => \N__14184\,
            in2 => \N__11884\,
            in3 => \N__14435\,
            lcout => \counter_RNI4HQB1Z0Z_5\,
            ltout => \counter_RNI4HQB1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100001111"
        )
    port map (
            in0 => \N__11881\,
            in1 => \N__14573\,
            in2 => \N__11872\,
            in3 => \N__14440\,
            lcout => \slaveselectZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4FVGV_4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14967\,
            in1 => \N__14280\,
            in2 => \_gnd_net_\,
            in3 => \N__12437\,
            lcout => OPEN,
            ltout => \beamY_RNI4FVGVZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7LOHP1_3_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__12599\,
            in2 => \N__11869\,
            in3 => \N__12856\,
            lcout => chary_if_generate_plus_mult1_un75_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_90_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12637\,
            in2 => \_gnd_net_\,
            in3 => \N__12859\,
            lcout => un5_visibley_3_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_49_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13075\,
            in2 => \_gnd_net_\,
            in3 => \N__13252\,
            lcout => \N_596_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_93_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12861\,
            in1 => \_gnd_net_\,
            in2 => \N__12669\,
            in3 => \N__12440\,
            lcout => OPEN,
            ltout => \un5_visibley_4_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_89_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010011000001"
        )
    port map (
            in0 => \N__14704\,
            in1 => \N__14966\,
            in2 => \N__11815\,
            in3 => \N__14274\,
            lcout => OPEN,
            ltout => \g1_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_83_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__12028\,
            in1 => \N__14705\,
            in2 => \N__12022\,
            in3 => \N__11992\,
            lcout => g1_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_94_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12439\,
            in1 => \N__12638\,
            in2 => \_gnd_net_\,
            in3 => \N__12860\,
            lcout => un5_visibley_1_0_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_0_4_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__12534\,
            in1 => \N__12746\,
            in2 => \N__12436\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_5_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__12533\,
            in1 => \N__12745\,
            in2 => \N__12435\,
            in3 => \N__12307\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0H2_4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12398\,
            in2 => \_gnd_net_\,
            in3 => \N__12532\,
            lcout => OPEN,
            ltout => \beamY_RNIJ0H2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITSR8_8_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010010101"
        )
    port map (
            in0 => \N__12078\,
            in1 => \N__12744\,
            in2 => \N__11917\,
            in3 => \N__11905\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJNLC_0_9_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001000100101"
        )
    port map (
            in0 => \N__13468\,
            in1 => \N__12079\,
            in2 => \N__11914\,
            in3 => \N__12151\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKOP3_7_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__12150\,
            in1 => \N__12225\,
            in2 => \_gnd_net_\,
            in3 => \N__12306\,
            lcout => un5_visibley_c6_0_0_0,
            ltout => \un5_visibley_c6_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12077\,
            in2 => \N__11899\,
            in3 => \N__11896\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_47_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__13076\,
            in1 => \N__13201\,
            in2 => \N__13105\,
            in3 => \_gnd_net_\,
            lcout => g2_1_1_0,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12804\,
            in2 => \_gnd_net_\,
            in3 => \N__12676\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13529\,
            in1 => \N__12585\,
            in2 => \_gnd_net_\,
            in3 => \N__12463\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13518\,
            in1 => \N__12432\,
            in2 => \_gnd_net_\,
            in3 => \N__12331\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__12256\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12240\,
            in2 => \_gnd_net_\,
            in3 => \N__12175\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13530\,
            in1 => \N__12163\,
            in2 => \_gnd_net_\,
            in3 => \N__12109\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12092\,
            in2 => \_gnd_net_\,
            in3 => \N__12031\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \N__13426\,
            ce => \N__13392\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__13466\,
            in1 => \N__13519\,
            in2 => \_gnd_net_\,
            in3 => \N__13489\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13424\,
            ce => \N__13393\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15273\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13303\,
            in2 => \N__15417\,
            in3 => \N__13324\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBC41_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15412\,
            in2 => \N__15649\,
            in3 => \N__13321\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIDBCZ0Z41\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEG81_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15625\,
            in2 => \N__15418\,
            in3 => \N__13318\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIMEGZ0Z81\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIFFA42_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13568\,
            in1 => \N__13309\,
            in2 => \N__15451\,
            in3 => \N__13315\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15416\,
            in1 => \N__15382\,
            in2 => \N__15436\,
            in3 => \N__13312\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15408\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15704\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14747\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13537\,
            in2 => \N__13569\,
            in3 => \N__13666\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13564\,
            in2 => \N__13663\,
            in3 => \N__13645\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4L02_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13642\,
            in2 => \N__13570\,
            in3 => \N__13624\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNII4LZ0Z02\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNISRO94_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13593\,
            in1 => \N__13543\,
            in2 => \N__13621\,
            in3 => \N__13606\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IU42_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13603\,
            in2 => \_gnd_net_\,
            in3 => \N__13597\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI0IUZ0Z42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13560\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15274\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram10__e_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14534\,
            lcout => content_ram10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14343\,
            ce => \N__13819\,
            sr => \_gnd_net_\
        );

    \content_content_ram10__e_0_RNO_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14113\,
            in1 => \N__13696\,
            in2 => \N__13765\,
            in3 => \N__14048\,
            lcout => content_awe10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIVRML1_0_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__13978\,
            in1 => \N__14442\,
            in2 => \N__13960\,
            in3 => \N__14390\,
            lcout => \content_N_35\,
            ltout => \content_N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIMIF92_1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__13695\,
            in1 => \N__14056\,
            in2 => \N__13810\,
            in3 => \N__14114\,
            lcout => content_awe3_1,
            ltout => \content_awe3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram2__0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__14533\,
            in1 => \N__14049\,
            in2 => \N__13801\,
            in3 => \N__13798\,
            lcout => content_ram2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram1__RNO_0_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__13915\,
            in1 => \N__14172\,
            in2 => \_gnd_net_\,
            in3 => \N__13781\,
            lcout => OPEN,
            ltout => \content_awe1_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \content_content_ram1__0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__13762\,
            in2 => \N__13729\,
            in3 => \N__13716\,
            lcout => content_ram1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIRAS9_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__14105\,
            in1 => \N__13948\,
            in2 => \N__14058\,
            in3 => \_gnd_net_\,
            lcout => un7_slaveselectlt5,
            ltout => \un7_slaveselectlt5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_3_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13702\,
            in3 => \N__13908\,
            lcout => \N_190_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIN1J6_4_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13849\,
            in2 => \_gnd_net_\,
            in3 => \N__13888\,
            lcout => slaveselect_1lto5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIAV5D_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__14106\,
            in1 => \N__13949\,
            in2 => \N__13916\,
            in3 => \N__13850\,
            lcout => un1_counter_0_1,
            ltout => \un1_counter_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI9UU01_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__14569\,
            in1 => \N__14170\,
            in2 => \N__14149\,
            in3 => \N__14142\,
            lcout => un5_slaveselect,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI0GS9_5_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14107\,
            in1 => \N__13950\,
            in2 => \_gnd_net_\,
            in3 => \N__14570\,
            lcout => OPEN,
            ltout => \slaveselect_1lto5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_RNIK7MV_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__14441\,
            in1 => \N__14359\,
            in2 => \N__14146\,
            in3 => \N__14143\,
            lcout => \SCLK1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIHRI6_0_1_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__14035\,
            in1 => \N__14108\,
            in2 => \N__14057\,
            in3 => \_gnd_net_\,
            lcout => un7_slaveselectlt2_0,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14610\,
            in1 => \N__13956\,
            in2 => \_gnd_net_\,
            in3 => \N__13921\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => counter_cry_1,
            carryout => counter_cry_2,
            clk => \N__14351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14606\,
            in1 => \N__13904\,
            in2 => \_gnd_net_\,
            in3 => \N__13855\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => counter_cry_2,
            carryout => counter_cry_3,
            clk => \N__14351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14611\,
            in1 => \N__13852\,
            in2 => \_gnd_net_\,
            in3 => \N__13831\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => counter_cry_3,
            carryout => counter_cry_4,
            clk => \N__14351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_5_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14607\,
            in1 => \N__14577\,
            in2 => \_gnd_net_\,
            in3 => \N__14584\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SDATAZ0Z2_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__14521\,
            in2 => \N__14443\,
            in3 => \N__14394\,
            lcout => \SDATA2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUR98A_9_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__14650\,
            in1 => \N__14875\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un75_sum_c5_m3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII78UP_4_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001111000110"
        )
    port map (
            in0 => \N__14785\,
            in1 => \N__14202\,
            in2 => \N__14305\,
            in3 => \N__14850\,
            lcout => \beamY_RNII78UPZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5VO45_6_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__15342\,
            in1 => \N__14782\,
            in2 => \_gnd_net_\,
            in3 => \N__15293\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axbxc4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI3R2DF_6_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14873\,
            in2 => \N__14290\,
            in3 => \N__14646\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc4_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFC5HA_1_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001111101"
        )
    port map (
            in0 => \N__14848\,
            in1 => \N__14874\,
            in2 => \N__14653\,
            in3 => \N__14783\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKBULF_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100011011"
        )
    port map (
            in0 => \N__15294\,
            in1 => \N__14786\,
            in2 => \N__14287\,
            in3 => \N__15343\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c5,
            ltout => \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIS5VDP1_4_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14203\,
            in1 => \N__15013\,
            in2 => \N__14194\,
            in3 => \N__14917\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFC5HA_0_4_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111010100"
        )
    port map (
            in0 => \N__14784\,
            in1 => \N__14849\,
            in2 => \N__14881\,
            in3 => \N__14651\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIOMEH5_0_9_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111110100"
        )
    port map (
            in0 => \N__15335\,
            in1 => \N__14787\,
            in2 => \N__15006\,
            in3 => \N__15291\,
            lcout => chary_if_generate_plus_mult1_un54_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIOMEH5_9_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__15336\,
            in1 => \N__14788\,
            in2 => \N__15007\,
            in3 => \N__15292\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axbxc5_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIMIOPF_9_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14642\,
            in2 => \N__14989\,
            in3 => \N__14879\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFC5HA_4_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14880\,
            in1 => \N__14851\,
            in2 => \N__14652\,
            in3 => \N__14789\,
            lcout => \beamY_RNIFC5HAZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI94I81_9_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011000011"
        )
    port map (
            in0 => \N__15180\,
            in1 => \N__15706\,
            in2 => \N__15322\,
            in3 => \N__15114\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axb4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI94I81_0_9_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011101011000"
        )
    port map (
            in0 => \N__15115\,
            in1 => \N__15708\,
            in2 => \N__15192\,
            in3 => \N__15319\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axbxc5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI65RM4_9_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110001101001"
        )
    port map (
            in0 => \N__15223\,
            in1 => \N__15364\,
            in2 => \N__14620\,
            in3 => \N__15352\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI94I81_1_9_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__15181\,
            in1 => \N__15705\,
            in2 => \N__15321\,
            in3 => \N__15113\,
            lcout => chary_if_generate_plus_mult1_un47_sum_ac0_8,
            ltout => \chary_if_generate_plus_mult1_un47_sum_ac0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI65RM4_0_9_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000111100"
        )
    port map (
            in0 => \N__15222\,
            in1 => \N__15363\,
            in2 => \N__15355\,
            in3 => \N__15351\,
            lcout => \beamY_RNI65RM4_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBO4T_9_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__15320\,
            in1 => \N__15280\,
            in2 => \_gnd_net_\,
            in3 => \N__15707\,
            lcout => chary_if_generate_plus_mult1_un47_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ7DB_0_9_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15179\,
            lcout => \beamY_RNIQ7DB_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15214\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STC_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15202\,
            in2 => \N__15550\,
            in3 => \N__15196\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI4STCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUC_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15193\,
            in2 => \N__15551\,
            in3 => \N__15133\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI5UUCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15130\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITSR8_0_8_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15112\,
            lcout => \beamY_RNITSR8_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15716\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJG_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15655\,
            in2 => \N__15598\,
            in3 => \N__15637\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI5QJGZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMK_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15575\,
            in2 => \N__15634\,
            in3 => \N__15616\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIDRMKZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOK_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15613\,
            in2 => \N__15599\,
            in3 => \N__15439\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIFVOKZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15377\,
            in2 => \_gnd_net_\,
            in3 => \N__15424\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15391\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15421\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15390\,
            in2 => \_gnd_net_\,
            in3 => \N__15378\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
