// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 23 2015 22:12:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__16788;
    wire N__16787;
    wire N__16786;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16761;
    wire N__16760;
    wire N__16759;
    wire N__16752;
    wire N__16751;
    wire N__16750;
    wire N__16743;
    wire N__16742;
    wire N__16741;
    wire N__16734;
    wire N__16733;
    wire N__16732;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16708;
    wire N__16705;
    wire N__16704;
    wire N__16701;
    wire N__16696;
    wire N__16691;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16639;
    wire N__16636;
    wire N__16635;
    wire N__16632;
    wire N__16625;
    wire N__16622;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16582;
    wire N__16581;
    wire N__16580;
    wire N__16579;
    wire N__16578;
    wire N__16577;
    wire N__16574;
    wire N__16563;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16539;
    wire N__16536;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16520;
    wire N__16517;
    wire N__16516;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16492;
    wire N__16491;
    wire N__16490;
    wire N__16487;
    wire N__16486;
    wire N__16485;
    wire N__16482;
    wire N__16471;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16403;
    wire N__16400;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16327;
    wire N__16326;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16249;
    wire N__16244;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16145;
    wire N__16140;
    wire N__16137;
    wire N__16136;
    wire N__16135;
    wire N__16132;
    wire N__16131;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16109;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16087;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16082;
    wire N__16081;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16071;
    wire N__16070;
    wire N__16067;
    wire N__16066;
    wire N__16065;
    wire N__16062;
    wire N__16061;
    wire N__16060;
    wire N__16059;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16052;
    wire N__16051;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16038;
    wire N__16037;
    wire N__16036;
    wire N__16035;
    wire N__16026;
    wire N__16019;
    wire N__16018;
    wire N__16017;
    wire N__16016;
    wire N__16015;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16011;
    wire N__16010;
    wire N__16009;
    wire N__16004;
    wire N__16003;
    wire N__15994;
    wire N__15981;
    wire N__15978;
    wire N__15967;
    wire N__15956;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15923;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15907;
    wire N__15894;
    wire N__15875;
    wire N__15874;
    wire N__15873;
    wire N__15870;
    wire N__15869;
    wire N__15868;
    wire N__15865;
    wire N__15864;
    wire N__15863;
    wire N__15862;
    wire N__15859;
    wire N__15858;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15850;
    wire N__15849;
    wire N__15848;
    wire N__15843;
    wire N__15842;
    wire N__15841;
    wire N__15836;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15817;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15811;
    wire N__15808;
    wire N__15807;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15795;
    wire N__15794;
    wire N__15793;
    wire N__15790;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15770;
    wire N__15767;
    wire N__15758;
    wire N__15751;
    wire N__15740;
    wire N__15729;
    wire N__15718;
    wire N__15707;
    wire N__15686;
    wire N__15685;
    wire N__15684;
    wire N__15683;
    wire N__15682;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15676;
    wire N__15675;
    wire N__15674;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15666;
    wire N__15665;
    wire N__15664;
    wire N__15663;
    wire N__15662;
    wire N__15661;
    wire N__15660;
    wire N__15659;
    wire N__15658;
    wire N__15657;
    wire N__15656;
    wire N__15655;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15645;
    wire N__15640;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15624;
    wire N__15619;
    wire N__15614;
    wire N__15609;
    wire N__15598;
    wire N__15595;
    wire N__15594;
    wire N__15593;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15584;
    wire N__15583;
    wire N__15582;
    wire N__15571;
    wire N__15568;
    wire N__15563;
    wire N__15560;
    wire N__15551;
    wire N__15542;
    wire N__15533;
    wire N__15526;
    wire N__15519;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15497;
    wire N__15496;
    wire N__15495;
    wire N__15494;
    wire N__15493;
    wire N__15492;
    wire N__15491;
    wire N__15482;
    wire N__15481;
    wire N__15480;
    wire N__15479;
    wire N__15478;
    wire N__15477;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15471;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15462;
    wire N__15453;
    wire N__15450;
    wire N__15439;
    wire N__15434;
    wire N__15427;
    wire N__15420;
    wire N__15415;
    wire N__15414;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15406;
    wire N__15403;
    wire N__15396;
    wire N__15391;
    wire N__15386;
    wire N__15385;
    wire N__15384;
    wire N__15383;
    wire N__15378;
    wire N__15373;
    wire N__15366;
    wire N__15363;
    wire N__15358;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15286;
    wire N__15285;
    wire N__15284;
    wire N__15281;
    wire N__15280;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15166;
    wire N__15165;
    wire N__15164;
    wire N__15163;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15146;
    wire N__15145;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15138;
    wire N__15137;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15129;
    wire N__15128;
    wire N__15127;
    wire N__15124;
    wire N__15119;
    wire N__15110;
    wire N__15109;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15103;
    wire N__15102;
    wire N__15101;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15066;
    wire N__15063;
    wire N__15058;
    wire N__15053;
    wire N__15052;
    wire N__15049;
    wire N__15038;
    wire N__15037;
    wire N__15036;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15001;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14981;
    wire N__14974;
    wire N__14969;
    wire N__14964;
    wire N__14961;
    wire N__14942;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14934;
    wire N__14931;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14925;
    wire N__14924;
    wire N__14923;
    wire N__14922;
    wire N__14921;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14909;
    wire N__14908;
    wire N__14907;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14873;
    wire N__14870;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14855;
    wire N__14854;
    wire N__14851;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14825;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14787;
    wire N__14784;
    wire N__14779;
    wire N__14776;
    wire N__14769;
    wire N__14760;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14703;
    wire N__14700;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14617;
    wire N__14616;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14565;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14545;
    wire N__14540;
    wire N__14537;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14518;
    wire N__14513;
    wire N__14504;
    wire N__14503;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14499;
    wire N__14498;
    wire N__14497;
    wire N__14494;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14475;
    wire N__14474;
    wire N__14471;
    wire N__14466;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14383;
    wire N__14382;
    wire N__14381;
    wire N__14380;
    wire N__14377;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14351;
    wire N__14350;
    wire N__14347;
    wire N__14346;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14330;
    wire N__14329;
    wire N__14326;
    wire N__14321;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14278;
    wire N__14277;
    wire N__14276;
    wire N__14275;
    wire N__14274;
    wire N__14273;
    wire N__14272;
    wire N__14271;
    wire N__14270;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14250;
    wire N__14247;
    wire N__14242;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14226;
    wire N__14223;
    wire N__14222;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14196;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14176;
    wire N__14173;
    wire N__14168;
    wire N__14165;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14140;
    wire N__14137;
    wire N__14126;
    wire N__14119;
    wire N__14116;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14011;
    wire N__14010;
    wire N__14007;
    wire N__14002;
    wire N__13997;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13960;
    wire N__13959;
    wire N__13958;
    wire N__13957;
    wire N__13956;
    wire N__13955;
    wire N__13954;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13948;
    wire N__13947;
    wire N__13946;
    wire N__13945;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13922;
    wire N__13919;
    wire N__13918;
    wire N__13909;
    wire N__13906;
    wire N__13901;
    wire N__13894;
    wire N__13893;
    wire N__13892;
    wire N__13891;
    wire N__13890;
    wire N__13889;
    wire N__13888;
    wire N__13887;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13875;
    wire N__13872;
    wire N__13857;
    wire N__13852;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13805;
    wire N__13802;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13756;
    wire N__13753;
    wire N__13752;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13644;
    wire N__13639;
    wire N__13636;
    wire N__13631;
    wire N__13616;
    wire N__13615;
    wire N__13614;
    wire N__13613;
    wire N__13610;
    wire N__13609;
    wire N__13606;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13578;
    wire N__13575;
    wire N__13570;
    wire N__13565;
    wire N__13562;
    wire N__13553;
    wire N__13552;
    wire N__13551;
    wire N__13550;
    wire N__13547;
    wire N__13546;
    wire N__13543;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13535;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13517;
    wire N__13508;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13420;
    wire N__13417;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13387;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13372;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13360;
    wire N__13353;
    wire N__13350;
    wire N__13343;
    wire N__13340;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13249;
    wire N__13248;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13147;
    wire N__13146;
    wire N__13145;
    wire N__13144;
    wire N__13143;
    wire N__13142;
    wire N__13141;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13137;
    wire N__13136;
    wire N__13135;
    wire N__13134;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13040;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12965;
    wire N__12964;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12766;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12749;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12595;
    wire N__12592;
    wire N__12591;
    wire N__12588;
    wire N__12583;
    wire N__12578;
    wire N__12577;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12391;
    wire N__12388;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12361;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12332;
    wire N__12331;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12271;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12260;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12256;
    wire N__12255;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12244;
    wire N__12237;
    wire N__12236;
    wire N__12235;
    wire N__12234;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12198;
    wire N__12191;
    wire N__12176;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12158;
    wire N__12155;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12143;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12113;
    wire N__12112;
    wire N__12109;
    wire N__12108;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12091;
    wire N__12090;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12063;
    wire N__12062;
    wire N__12061;
    wire N__12060;
    wire N__12059;
    wire N__12058;
    wire N__12055;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12034;
    wire N__12027;
    wire N__12022;
    wire N__12019;
    wire N__12012;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11878;
    wire N__11877;
    wire N__11874;
    wire N__11869;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11854;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11830;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11824;
    wire N__11823;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11815;
    wire N__11812;
    wire N__11811;
    wire N__11810;
    wire N__11809;
    wire N__11808;
    wire N__11805;
    wire N__11800;
    wire N__11797;
    wire N__11796;
    wire N__11795;
    wire N__11794;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11782;
    wire N__11781;
    wire N__11780;
    wire N__11777;
    wire N__11776;
    wire N__11773;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11759;
    wire N__11756;
    wire N__11751;
    wire N__11748;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11729;
    wire N__11726;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11698;
    wire N__11693;
    wire N__11686;
    wire N__11683;
    wire N__11678;
    wire N__11677;
    wire N__11674;
    wire N__11673;
    wire N__11672;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11645;
    wire N__11642;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11622;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11602;
    wire N__11597;
    wire N__11594;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11570;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11554;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11539;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11510;
    wire N__11509;
    wire N__11508;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11496;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11466;
    wire N__11453;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11404;
    wire N__11401;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11376;
    wire N__11375;
    wire N__11374;
    wire N__11371;
    wire N__11370;
    wire N__11369;
    wire N__11368;
    wire N__11367;
    wire N__11366;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11337;
    wire N__11334;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11330;
    wire N__11329;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11307;
    wire N__11304;
    wire N__11295;
    wire N__11288;
    wire N__11285;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11255;
    wire N__11250;
    wire N__11245;
    wire N__11242;
    wire N__11237;
    wire N__11234;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11191;
    wire N__11190;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11170;
    wire N__11163;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11052;
    wire N__11051;
    wire N__11050;
    wire N__11049;
    wire N__11044;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10997;
    wire N__10994;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10943;
    wire N__10938;
    wire N__10935;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10915;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10856;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10846;
    wire N__10843;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10751;
    wire N__10748;
    wire N__10739;
    wire N__10738;
    wire N__10737;
    wire N__10736;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10715;
    wire N__10712;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10687;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10613;
    wire N__10610;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10568;
    wire N__10567;
    wire N__10566;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10560;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10541;
    wire N__10538;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10490;
    wire N__10489;
    wire N__10488;
    wire N__10487;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10444;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10310;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10302;
    wire N__10301;
    wire N__10296;
    wire N__10295;
    wire N__10292;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10262;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10254;
    wire N__10253;
    wire N__10250;
    wire N__10249;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10212;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10200;
    wire N__10199;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10155;
    wire N__10152;
    wire N__10147;
    wire N__10142;
    wire N__10137;
    wire N__10128;
    wire N__10119;
    wire N__10106;
    wire N__10105;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10044;
    wire N__10037;
    wire N__10034;
    wire N__10029;
    wire N__10022;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10017;
    wire N__10016;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9986;
    wire N__9985;
    wire N__9984;
    wire N__9981;
    wire N__9976;
    wire N__9973;
    wire N__9962;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9948;
    wire N__9943;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9891;
    wire N__9888;
    wire N__9883;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9868;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9853;
    wire N__9852;
    wire N__9851;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9844;
    wire N__9843;
    wire N__9840;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9822;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9799;
    wire N__9798;
    wire N__9793;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9722;
    wire N__9721;
    wire N__9718;
    wire N__9717;
    wire N__9714;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9702;
    wire N__9695;
    wire N__9692;
    wire N__9691;
    wire N__9690;
    wire N__9689;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9677;
    wire N__9674;
    wire N__9673;
    wire N__9672;
    wire N__9671;
    wire N__9670;
    wire N__9665;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9640;
    wire N__9637;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9616;
    wire N__9615;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9600;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9588;
    wire N__9585;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9530;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9516;
    wire N__9511;
    wire N__9510;
    wire N__9507;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9488;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9478;
    wire N__9473;
    wire N__9468;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9452;
    wire N__9447;
    wire N__9442;
    wire N__9431;
    wire N__9430;
    wire N__9427;
    wire N__9426;
    wire N__9425;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9382;
    wire N__9377;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9346;
    wire N__9345;
    wire N__9344;
    wire N__9341;
    wire N__9340;
    wire N__9337;
    wire N__9336;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9320;
    wire N__9315;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9290;
    wire N__9287;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9269;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9257;
    wire N__9248;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9179;
    wire N__9176;
    wire N__9175;
    wire N__9174;
    wire N__9171;
    wire N__9166;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9151;
    wire N__9150;
    wire N__9149;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9134;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9117;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9111;
    wire N__9110;
    wire N__9109;
    wire N__9106;
    wire N__9105;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9092;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9062;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9044;
    wire N__9041;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9012;
    wire N__9003;
    wire N__8998;
    wire N__8987;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8918;
    wire N__8915;
    wire N__8908;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8860;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8808;
    wire N__8807;
    wire N__8806;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8787;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8765;
    wire N__8764;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8741;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8652;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8640;
    wire N__8637;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8620;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8592;
    wire N__8589;
    wire N__8582;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8578;
    wire N__8577;
    wire N__8572;
    wire N__8571;
    wire N__8566;
    wire N__8561;
    wire N__8558;
    wire N__8557;
    wire N__8556;
    wire N__8553;
    wire N__8552;
    wire N__8547;
    wire N__8544;
    wire N__8535;
    wire N__8528;
    wire N__8525;
    wire N__8524;
    wire N__8523;
    wire N__8522;
    wire N__8521;
    wire N__8518;
    wire N__8509;
    wire N__8506;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8488;
    wire N__8487;
    wire N__8486;
    wire N__8483;
    wire N__8482;
    wire N__8481;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8475;
    wire N__8472;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8464;
    wire N__8463;
    wire N__8462;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8378;
    wire N__8375;
    wire N__8370;
    wire N__8357;
    wire N__8356;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8317;
    wire N__8316;
    wire N__8315;
    wire N__8312;
    wire N__8311;
    wire N__8308;
    wire N__8307;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8286;
    wire N__8279;
    wire N__8270;
    wire N__8269;
    wire N__8264;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8233;
    wire N__8230;
    wire N__8225;
    wire N__8220;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8164;
    wire N__8163;
    wire N__8160;
    wire N__8155;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8089;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8065;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8030;
    wire N__8027;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7966;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7937;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7919;
    wire N__7918;
    wire N__7917;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7899;
    wire N__7896;
    wire N__7891;
    wire N__7886;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7861;
    wire N__7860;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7838;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7821;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7771;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7756;
    wire N__7751;
    wire N__7748;
    wire N__7747;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7678;
    wire N__7677;
    wire N__7674;
    wire N__7669;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7651;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7643;
    wire N__7642;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7621;
    wire N__7618;
    wire N__7617;
    wire N__7616;
    wire N__7615;
    wire N__7608;
    wire N__7603;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7549;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7522;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7392;
    wire N__7391;
    wire N__7390;
    wire N__7385;
    wire N__7382;
    wire N__7377;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7357;
    wire N__7350;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7327;
    wire N__7326;
    wire N__7319;
    wire N__7312;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7279;
    wire N__7278;
    wire N__7275;
    wire N__7274;
    wire N__7271;
    wire N__7270;
    wire N__7269;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7257;
    wire N__7254;
    wire N__7249;
    wire N__7246;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7225;
    wire N__7224;
    wire N__7223;
    wire N__7216;
    wire N__7213;
    wire N__7208;
    wire N__7205;
    wire N__7204;
    wire N__7203;
    wire N__7200;
    wire N__7199;
    wire N__7190;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7178;
    wire N__7175;
    wire N__7174;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7111;
    wire N__7110;
    wire N__7107;
    wire N__7106;
    wire N__7103;
    wire N__7102;
    wire N__7099;
    wire N__7090;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7014;
    wire N__7013;
    wire N__7012;
    wire N__7009;
    wire N__7000;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6961;
    wire N__6958;
    wire N__6957;
    wire N__6956;
    wire N__6949;
    wire N__6946;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire Clock12MHz_c;
    wire \Clock50MHz.PixelClock ;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_4_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_;
    wire bfn_1_5_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0;
    wire bfn_1_6_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7;
    wire bfn_1_7_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0;
    wire chary_if_generate_plus_mult1_un47_sum_axb4_cascade_;
    wire beamY_RNIKM9GCZ0Z_9_cascade_;
    wire beamY_RNIM5433Z0Z_8;
    wire beamY_RNI93821Z0Z_9_cascade_;
    wire beamY_RNIM5433_0Z0Z_8;
    wire beamY_RNIIR4K3_0Z0Z_7;
    wire beamY_RNIIR4K3_0Z0Z_7_cascade_;
    wire beamY_RNIKM9GC_0Z0Z_9;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_;
    wire beamY_RNI9DSP2_0Z0Z_8;
    wire beamY_RNI41384Z0Z_7_cascade_;
    wire chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_;
    wire un8_beamylt9_0_cascade_;
    wire beamY_RNIP8FF1_1Z0Z_7;
    wire beamY_RNI93821Z0Z_9;
    wire beamY_RNIBV5E51Z0Z_8_cascade_;
    wire beamY_RNIBV5E51_0Z0Z_8;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_2;
    wire chary_if_generate_plus_mult1_un47_sum_c5;
    wire beamY_RNIVADQVZ0Z_8_cascade_;
    wire chary_if_generate_plus_mult1_un54_sum_ac0_5;
    wire beamY_RNIV5SUC3_0Z0Z_9_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_0_1;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_;
    wire beamY_RNIVADQVZ0Z_8;
    wire chary_if_generate_plus_mult1_un47_sum_c4;
    wire chary_if_generate_plus_mult1_un47_sum_axb4;
    wire beamY_RNIV5SUC3Z0Z_9;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_;
    wire g1_0_2;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_0;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_i_0;
    wire g1_1;
    wire g2_0_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_;
    wire un114_pixel_6_1_5__g0Z0Z_2;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_0;
    wire chary_if_generate_plus_mult1_un61_sum_c4_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb3_0;
    wire beamY_RNISDTA58Z0Z_5_cascade_;
    wire beamY_RNIJ0797KZ0Z_4;
    wire bfn_2_2_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5;
    wire beamY_RNI2B511_0Z0Z_9;
    wire bfn_2_3_0_;
    wire beamY_RNIUUEM_0Z0Z_8;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire bfn_2_4_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7;
    wire if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0;
    wire chary_if_generate_plus_mult1_un47_sum_axb3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0;
    wire beamY_i_2_cascade_;
    wire beamY_fast_RNIT5UFZ0Z_4_cascade_;
    wire un5_visibley_ac0_7;
    wire un5_visibley_ac0_7_cascade_;
    wire chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux;
    wire beamY_fastZ0Z_7;
    wire beamY_fastZ0Z_6;
    wire beamY_fastZ0Z_5;
    wire un5_visibley_ac0_11_0_1_cascade_;
    wire beamY_fastZ0Z_4;
    wire beamY_fastZ0Z_8;
    wire un5_visibley_c7;
    wire beamY_fastZ0Z_3;
    wire un5_visibley_c2_cascade_;
    wire beamY_fastZ0Z_2;
    wire bfn_2_12_0_;
    wire un21_beamy_cry_1_c_RNIALZ0Z73;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_2_c_RNICOZ0Z83;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3_c_RNIERZ0Z93;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4_c_RNIGUAZ0Z3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5_c_RNII1CZ0Z3;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6_c_RNIK4DZ0Z3;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7_c_RNIM7EZ0Z3;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire bfn_2_13_0_;
    wire if_generate_plus_mult1_un61_sum_axbxc5_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_c5_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_axb4_i;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1;
    wire row_1_if_i4_mux_i_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3;
    wire row_1_if_i4_mux_i;
    wire row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_;
    wire row_1_if_N_6;
    wire if_generate_plus_mult1_un75_sum_axbxc3_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_;
    wire row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0;
    wire if_generate_plus_mult1_un75_sum_axbxc3;
    wire row_1_if_generate_plus_mult1_un75_sum_c5;
    wire if_generate_plus_mult1_un82_sum_axb4_x1_cascade_;
    wire if_generate_plus_mult1_un82_sum_axb4_x0;
    wire beamY_RNIP8FF1_0Z0Z_7;
    wire un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_;
    wire un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_;
    wire beamY_RNIP8FF1Z0Z_7_cascade_;
    wire un5_visibley_c6;
    wire chary_if_generate_plus_mult1_un40_sum_c4;
    wire un5_visibley_c5;
    wire beamY_RNIP8FF1_2Z0Z_7;
    wire un4_beamylt6_cascade_;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1;
    wire chary_if_generate_plus_mult1_un54_sum_c5;
    wire beamY_RNIB6AOI5_0Z0Z_5_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_d;
    wire un5_visibley_c2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum;
    wire g2_1;
    wire chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_;
    wire chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_;
    wire chary_if_generate_plus_mult1_un54_sum_axb3;
    wire chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_0;
    wire chary_if_generate_plus_mult1_un68_sum_c5_0_0;
    wire un114_pixel_6_1_5__g0_17Z0Z_1_cascade_;
    wire chary_if_generate_plus_mult1_un75_sum_0_5;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_i;
    wire chary_if_generate_plus_mult1_un61_sum_c4;
    wire g1_0_3;
    wire bfn_5_4_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8;
    wire bfn_5_5_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i;
    wire bfn_5_6_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_5_7_0_;
    wire un8_beamx_cry_9;
    wire row_1_if_generate_plus_mult1_un82_sum_axb4_i;
    wire un114_pixel_6_1_5__un8_beamylto9Z0Z_0;
    wire un8_beamylt9_0;
    wire un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_;
    wire un114_pixel_6_1_5__un1_beamylto9_3_cascade_;
    wire VSync_c;
    wire un8_beamy_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_c5;
    wire row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum;
    wire un4_beamylt8_0;
    wire un114_pixel_6_1_5__g0_1Z0Z_4_cascade_;
    wire beamYZ0Z_5;
    wire beamYZ0Z_9;
    wire beamYZ0Z_7;
    wire beamYZ0Z_6;
    wire un114_pixel_6_1_5__g0_0Z0Z_4;
    wire un114_pixel_6_1_5__g0_0Z0Z_3_cascade_;
    wire un114_pixel_6_1_5__g2_0Z0Z_0_cascade_;
    wire beamYZ0Z_8;
    wire un114_pixel_6_1_5__g0_0_1Z0Z_1;
    wire g1;
    wire beamYZ0Z_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_;
    wire m511_0_x2_1_2;
    wire G_7_0_m2_1_1_1_cascade_;
    wire G_7_0_m2_1_1_cascade_;
    wire G_7_0_m2_1_0;
    wire chary_if_generate_plus_mult1_un75_sum_c5;
    wire chary_if_generate_plus_mult1_un68_sum_c4;
    wire chary_if_generate_plus_mult1_un61_sum_c5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_1;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_5;
    wire chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_;
    wire beamY_RNIL0E2QG2Z0Z_3;
    wire bfn_6_4_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i;
    wire bfn_6_5_0_;
    wire un5_visiblex_cry_0;
    wire un5_visiblex_cry_1;
    wire un5_visiblex_cry_2;
    wire un5_visiblex_cry_3;
    wire un5_visiblex_cry_4;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire bfn_6_6_0_;
    wire un5_visiblex_cry_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0;
    wire if_generate_plus_mult1_un54_sum_axbxc5;
    wire if_generate_plus_mult1_un61_sum_axbxc5;
    wire un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_;
    wire un114_pixel_6_1_5__un3_beamxZ0Z_7;
    wire un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0;
    wire un4_beamy_0;
    wire un13_beamylt10_0_cascade_;
    wire beamXZ0Z_4;
    wire beamXZ0Z_3;
    wire un18_beamylt5_0;
    wire beamXZ0Z_5;
    wire un18_beamylt5_0_cascade_;
    wire un114_pixel_6_1_5__un15_beamyZ0Z_0;
    wire beamXZ0Z_8;
    wire beamXZ0Z_9;
    wire beamXZ0Z_6;
    wire un114_pixel_6_1_5__un18_beamylto9Z0Z_2;
    wire beamXZ0Z_2;
    wire beamXZ0Z_1;
    wire un114_pixel_6_1_5__un13_beamylto2Z0Z_0;
    wire un114_pixel_6_1_5__un15_beamyZ0Z_1;
    wire un4_beamy_0_0;
    wire un114_pixel_6_1_5__g3_0_0_0;
    wire un13_beamylt10_0;
    wire un1_beamx_2;
    wire beamXZ0Z_7;
    wire beamXZ0Z_10;
    wire un1_beamxlt10_0;
    wire HSync_c;
    wire un114_pixel_6_1_5__un4_rowZ0Z_5;
    wire row_1_if_generate_plus_mult1_un68_sum_c5;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1;
    wire if_generate_plus_mult1_un75_sum_axbxc5;
    wire row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3;
    wire un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_;
    wire un114_pixel_6_1_5__un4_rowZ0Z_1;
    wire beamY_i_2;
    wire un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0;
    wire chessboardpixel_un200_pixellt10_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5;
    wire chary_if_generate_plus_mult1_un68_sum_c5_0;
    wire chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_;
    wire g1_0_1;
    wire beamYZ0Z_3;
    wire chary_if_generate_plus_mult1_un68_sum_axb4_i;
    wire g2;
    wire m511_0_o2_1;
    wire chary_if_generate_plus_mult1_un68_sum_axbxc5_0;
    wire N_80_i;
    wire un3_beamx_0;
    wire un5_beamx_0;
    wire beamYZ0Z_2;
    wire chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0;
    wire beamY_RNIJH2N2PZ0Z_3;
    wire bfn_7_3_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8;
    wire bfn_7_4_0_;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_1;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_2;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_3;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_4;
    wire column_1_if_generate_plus_mult1_un47_sum1_5_cascade_;
    wire un5_visiblex_i_0_25;
    wire charx_if_generate_plus_mult1_un26_sum_axb_3_i;
    wire column_1_if_generate_plus_mult1_un47_sum1_4;
    wire column_1_if_generate_plus_mult1_un47_sum1_3;
    wire if_generate_plus_mult1_un47_sum_m_5_cascade_;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_;
    wire N_11_0_i;
    wire if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3;
    wire chary_if_generate_plus_mult1_un33_sum_axb3;
    wire un114_pixel_6_1_5__un4_rowZ0Z_2;
    wire bfn_7_7_0_;
    wire if_generate_plus_mult1_un47_sum_m_1;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_1;
    wire if_generate_plus_mult1_un47_sum_m_5;
    wire if_generate_plus_mult1_un47_sum_m_2;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_2;
    wire if_generate_plus_mult1_un54_sum_axb_4_l_fx;
    wire N_571_i;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_4;
    wire if_generate_plus_mult1_un54_sum_s_5_cascade_;
    wire bfn_7_8_0_;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_s_5;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un54_sum_i_5;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_4;
    wire N_562_i;
    wire chessboardpixel_un174_pixel_0_1;
    wire chessboardpixel_un200_pixel_0_1;
    wire un114_pixel_6_1_5__un4_row_7Z0Z_1;
    wire N_357_0;
    wire N_18_0_cascade_;
    wire N_7_0_cascade_;
    wire font_un28_pixel_0_0_29;
    wire un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_;
    wire N_14_0;
    wire column_0111_0_cascade_;
    wire beamY_RNI05CI5A3_0Z0Z_0_cascade_;
    wire beamY_RNIBABJS01Z0Z_1_cascade_;
    wire N_21_0_cascade_;
    wire N_22_0;
    wire column_0111_0;
    wire un116_pixel_3_bmZ0Z_6_cascade_;
    wire beamY_RNISJITRQ2Z0Z_1_cascade_;
    wire N_12_0;
    wire N_248_0_cascade_;
    wire un116_pixel_3_ns_1_0_6;
    wire N_25_mux;
    wire un114_pixel_3_i_a3_7_cascade_;
    wire column_0001_0;
    wire un116_pixel_3_ns_1_2_cascade_;
    wire beamY_RNIDVSK5A3Z0Z_1;
    wire N_13_0;
    wire un114_pixel_0_1__N_6_mux_0;
    wire un116_pixel_1_amZ0Z_1_cascade_;
    wire un116_pixel_4_bmZ0Z_1;
    wire un116_pixel_4_amZ0Z_1_cascade_;
    wire un116_pixel_3_ns_1_1;
    wire beamY_RNIHIRVUS1Z0Z_1;
    wire un116_pixel_1_bmZ0Z_1;
    wire bfn_8_3_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i;
    wire bfn_8_4_0_;
    wire column_1_if_generate_plus_mult1_un47_sum0_2;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_1;
    wire column_1_if_generate_plus_mult1_un47_sum0_3;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_2;
    wire column_1_if_generate_plus_mult1_un47_sum0_4;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_3;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_4;
    wire if_generate_plus_mult1_un47_sum_0_cry_3_ma;
    wire if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx;
    wire N_200_0_i;
    wire bfn_8_5_0_;
    wire charx_if_generate_plus_mult1_un26_sum_s_2_sf;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4;
    wire if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx;
    wire un5_visiblex_i_25;
    wire column_1_if_generate_plus_mult1_un47_sum0_5;
    wire column_1_if_generate_plus_mult1_un47_sum1_5;
    wire un114_pixel_6_1_5__un4_rowZ0Z_0;
    wire un116_pixel_5_amZ0Z_6_cascade_;
    wire un116_pixel_5_bmZ0Z_6;
    wire un15_beamy;
    wire un114_pixel_6_1_5__g0Z0Z_0;
    wire un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_;
    wire un114_pixel_6_1_5__font_un126_pixel_m_4_1_0;
    wire un114_pixel_6_1_5__g0_2Z0Z_0_cascade_;
    wire un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0;
    wire un114_pixel_6_1_5__g0_1_0;
    wire un114_pixel_6_1_5__g1Z0Z_0_cascade_;
    wire un4_row;
    wire beamY_RNIPG1SS93Z0Z_2;
    wire N_23_0;
    wire N_15_0;
    wire N_342_0_0;
    wire N_1045_0_cascade_;
    wire bfn_8_10_0_;
    wire column_1_if_generate_plus_mult1_un61_sum_iZ0;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_1;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_2;
    wire un5_rowlto3_i;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_4;
    wire Pixel_3_sqmuxa;
    wire un114_pixel_6_1_5__font_un126_pixel_m_4;
    wire un1_beamy_0_0;
    wire Pixel_1_r_sn;
    wire Pixel_1_r_rn_0_cascade_;
    wire N_396;
    wire Pixel_c;
    wire PixelClock_g;
    wire m6Z0Z_1;
    wire G_7_0_m2_1;
    wire beamX_RNI1M3Q1V2Z0Z_0_cascade_;
    wire N_1039_0_0;
    wire font_un3_pixel_29_cascade_;
    wire G_7_0_m4_2_1_1_cascade_;
    wire G_7_0_m4_2_1;
    wire beamY_RNINIKJ5A3Z0Z_1;
    wire beamY_RNI7OTDJ61Z0Z_1_cascade_;
    wire beamY_RNIJDHE4C2Z0Z_1;
    wire font_un126_pixel_6_am_cascade_;
    wire font_un126_pixel_2_am;
    wire beamX_RNIQ6MATS2Z0Z_0;
    wire un114_pixel_7_1_7__N_11_i_1;
    wire N_37_cascade_;
    wire beamY_RNI05CI5A3_1Z0Z_0_cascade_;
    wire beamY_RNI05CI5A3Z0Z_0;
    wire beamY_RNII25UDD3_1Z0Z_0;
    wire un116_pixel_7_ns_1_4_cascade_;
    wire beamY_RNIFHEQCT1Z0Z_0;
    wire beamY_RNIA4V0NM1Z0Z_0_cascade_;
    wire beamY_RNII25UDD3_0Z0Z_0;
    wire un116_pixel_7_ns_1_6_cascade_;
    wire font_un3_pixel_29;
    wire beamY_RNIBHJ7AMZ0Z_0;
    wire bfn_8_13_0_;
    wire column_1_if_generate_plus_mult1_un75_sum_iZ0;
    wire G_340;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_1;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_2;
    wire G_341;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_4;
    wire un5_rowlto0_cascade_;
    wire beamY_RNIJ720T72Z0Z_0;
    wire un116_pixel_5_ns_1_2;
    wire bfn_8_14_0_;
    wire column_1_if_generate_plus_mult1_un68_sum_iZ0;
    wire if_generate_plus_mult1_un75_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_4;
    wire un116_pixel_2_ns_1_2;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire if_generate_plus_mult1_un75_sum_axb_4_l_fx;
    wire bfn_9_3_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0;
    wire if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx;
    wire bfn_9_4_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO;
    wire charx_if_generate_plus_mult1_un33_sum;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum;
    wire N_520;
    wire bfn_9_5_0_;
    wire un5_visiblex_i_24;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538;
    wire charx_if_generate_plus_mult1_un33_sum_cry_3;
    wire CO3_0;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5;
    wire bfn_9_6_0_;
    wire charx_if_generate_plus_mult1_un33_sum_i;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0;
    wire charx_if_generate_plus_mult1_un33_sum_i_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_3;
    wire charx_if_generate_plus_mult1_un40_sum_axb_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4;
    wire bfn_9_7_0_;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1;
    wire charx_if_generate_plus_mult1_un47_sum_cry_3;
    wire charx_if_generate_plus_mult1_un47_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1;
    wire charx_if_generate_plus_mult1_un40_sum_i_5;
    wire charx_if_generate_plus_mult1_un40_sum;
    wire charx_if_generate_plus_mult1_un40_sum_i;
    wire bfn_9_9_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1;
    wire CONSTANT_ONE_NET;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4;
    wire un114_pixel_6_1_5__g2_0_1;
    wire bfn_9_10_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_;
    wire un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1;
    wire charx_if_generate_plus_mult1_un1_sum_axb1;
    wire beamXZ0Z_0;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1;
    wire charx_if_generate_plus_mult1_un1_sum_axb1_cascade_;
    wire un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1;
    wire m15_cascade_;
    wire un114_pixel_0_1__N_6_mux;
    wire beamY_RNI4NRC8D1Z0Z_0_cascade_;
    wire beamY_RNII25UDD3Z0Z_0;
    wire N_14;
    wire un116_pixel_2_ns_1_6_cascade_;
    wire beamY_RNIH01F2SZ0Z_0;
    wire un116_pixel_2_ns_1Z0Z_5;
    wire N_276_0_cascade_;
    wire beamY_RNII25UDD3_3Z0Z_0;
    wire m7;
    wire m7_cascade_;
    wire N_302_i_0;
    wire beamY_RNITQPUS72Z0Z_0_cascade_;
    wire un116_pixel_3_1_0;
    wire beamY_RNI6B7UAL1Z0Z_1;
    wire m31;
    wire un116_pixel_4_1Z0Z_0;
    wire m38;
    wire beamYZ0Z_0;
    wire m38_cascade_;
    wire beamYZ0Z_1;
    wire un116_pixel_6_1_1_cascade_;
    wire N_17;
    wire N_321;
    wire un116_pixel_2_bmZ0Z_1;
    wire un5_rowlto2_i;
    wire un5_rowlto2;
    wire un5_rowlto0;
    wire un5_rowlto1;
    wire un5_rowlto3;
    wire un116_pixel_2_amZ0Z_1;
    wire bfn_11_5_0_;
    wire charx_if_generate_plus_mult1_un47_sum_i_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2;
    wire charx_if_generate_plus_mult1_un54_sum_cry_3;
    wire charx_if_generate_plus_mult1_un54_sum_axb_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_;
    wire charx_if_generate_plus_mult1_un47_sum;
    wire charx_if_generate_plus_mult1_un47_sum_i;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6;
    wire bfn_11_6_0_;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5;
    wire charx_if_generate_plus_mult1_un54_sum_i_5;
    wire charx_if_generate_plus_mult1_un61_sum_cry_3;
    wire charx_if_generate_plus_mult1_un61_sum_axb_5;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_;
    wire charx_if_generate_plus_mult1_un54_sum;
    wire charx_if_generate_plus_mult1_un54_sum_i;
    wire charx_if_generate_plus_mult1_un68_sum;
    wire bfn_11_7_0_;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0;
    wire charx_if_generate_plus_mult1_un61_sum_i_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_3;
    wire charx_if_generate_plus_mult1_un68_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un152_pixel_24;
    wire charx_if_generate_plus_mult1_un61_sum_i;
    wire bfn_11_8_0_;
    wire charx_if_generate_plus_mult1_un68_sum_i;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0;
    wire charx_if_generate_plus_mult1_un68_sum_i_5;
    wire charx_if_generate_plus_mult1_un75_sum_cry_3;
    wire charx_if_generate_plus_mult1_un75_sum_axb_5;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4;
    wire charx_i_24;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf;
    wire charx_i_23;
    wire charx_if_generate_plus_mult1_un75_sum;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__6839),
            .RESETB(N__14250),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__16788),
            .DIN(N__16787),
            .DOUT(N__16786),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__16788),
            .PADOUT(N__16787),
            .PADIN(N__16786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9202),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__16779),
            .DIN(N__16778),
            .DOUT(N__16777),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__16779),
            .PADOUT(N__16778),
            .PADIN(N__16777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__16770),
            .DIN(N__16769),
            .DOUT(N__16768),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__16770),
            .PADOUT(N__16769),
            .PADIN(N__16768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13178),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__16761),
            .DIN(N__16760),
            .DOUT(N__16759),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__16761),
            .PADOUT(N__16760),
            .PADIN(N__16759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9209),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__16752),
            .DIN(N__16751),
            .DOUT(N__16750),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__16752),
            .PADOUT(N__16751),
            .PADIN(N__16750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__16743),
            .DIN(N__16742),
            .DOUT(N__16741),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__16743),
            .PADOUT(N__16742),
            .PADIN(N__16741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11102),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__16734),
            .DIN(N__16733),
            .DOUT(N__16732),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__16734),
            .PADOUT(N__16733),
            .PADIN(N__16732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3889 (
            .O(N__16715),
            .I(N__16712));
    LocalMux I__3888 (
            .O(N__16712),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0));
    CascadeMux I__3887 (
            .O(N__16709),
            .I(N__16705));
    InMux I__3886 (
            .O(N__16708),
            .I(N__16701));
    InMux I__3885 (
            .O(N__16705),
            .I(N__16696));
    InMux I__3884 (
            .O(N__16704),
            .I(N__16696));
    LocalMux I__3883 (
            .O(N__16701),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0));
    LocalMux I__3882 (
            .O(N__16696),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0));
    CascadeMux I__3881 (
            .O(N__16691),
            .I(N__16687));
    CascadeMux I__3880 (
            .O(N__16690),
            .I(N__16684));
    InMux I__3879 (
            .O(N__16687),
            .I(N__16679));
    InMux I__3878 (
            .O(N__16684),
            .I(N__16679));
    LocalMux I__3877 (
            .O(N__16679),
            .I(charx_if_generate_plus_mult1_un68_sum_i_5));
    CascadeMux I__3876 (
            .O(N__16676),
            .I(N__16673));
    InMux I__3875 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__3874 (
            .O(N__16670),
            .I(charx_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__3873 (
            .O(N__16667),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__3872 (
            .O(N__16664),
            .I(N__16661));
    InMux I__3871 (
            .O(N__16661),
            .I(N__16658));
    LocalMux I__3870 (
            .O(N__16658),
            .I(N__16655));
    Odrv4 I__3869 (
            .O(N__16655),
            .I(charx_i_24));
    CascadeMux I__3868 (
            .O(N__16652),
            .I(N__16649));
    InMux I__3867 (
            .O(N__16649),
            .I(N__16646));
    LocalMux I__3866 (
            .O(N__16646),
            .I(N__16643));
    Odrv4 I__3865 (
            .O(N__16643),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0));
    CascadeMux I__3864 (
            .O(N__16640),
            .I(N__16636));
    CascadeMux I__3863 (
            .O(N__16639),
            .I(N__16632));
    InMux I__3862 (
            .O(N__16636),
            .I(N__16625));
    InMux I__3861 (
            .O(N__16635),
            .I(N__16625));
    InMux I__3860 (
            .O(N__16632),
            .I(N__16625));
    LocalMux I__3859 (
            .O(N__16625),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1));
    InMux I__3858 (
            .O(N__16622),
            .I(N__16618));
    CascadeMux I__3857 (
            .O(N__16621),
            .I(N__16615));
    LocalMux I__3856 (
            .O(N__16618),
            .I(N__16612));
    InMux I__3855 (
            .O(N__16615),
            .I(N__16609));
    Span4Mux_h I__3854 (
            .O(N__16612),
            .I(N__16606));
    LocalMux I__3853 (
            .O(N__16609),
            .I(N__16603));
    Odrv4 I__3852 (
            .O(N__16606),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    Odrv4 I__3851 (
            .O(N__16603),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    CascadeMux I__3850 (
            .O(N__16598),
            .I(N__16595));
    InMux I__3849 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__3848 (
            .O(N__16592),
            .I(N__16589));
    Span4Mux_h I__3847 (
            .O(N__16589),
            .I(N__16586));
    Odrv4 I__3846 (
            .O(N__16586),
            .I(charx_i_23));
    InMux I__3845 (
            .O(N__16583),
            .I(N__16574));
    InMux I__3844 (
            .O(N__16582),
            .I(N__16563));
    InMux I__3843 (
            .O(N__16581),
            .I(N__16563));
    InMux I__3842 (
            .O(N__16580),
            .I(N__16563));
    InMux I__3841 (
            .O(N__16579),
            .I(N__16563));
    InMux I__3840 (
            .O(N__16578),
            .I(N__16563));
    InMux I__3839 (
            .O(N__16577),
            .I(N__16559));
    LocalMux I__3838 (
            .O(N__16574),
            .I(N__16556));
    LocalMux I__3837 (
            .O(N__16563),
            .I(N__16553));
    InMux I__3836 (
            .O(N__16562),
            .I(N__16550));
    LocalMux I__3835 (
            .O(N__16559),
            .I(N__16547));
    Span4Mux_v I__3834 (
            .O(N__16556),
            .I(N__16544));
    Span4Mux_h I__3833 (
            .O(N__16553),
            .I(N__16539));
    LocalMux I__3832 (
            .O(N__16550),
            .I(N__16539));
    Span4Mux_h I__3831 (
            .O(N__16547),
            .I(N__16536));
    Span4Mux_v I__3830 (
            .O(N__16544),
            .I(N__16531));
    Span4Mux_v I__3829 (
            .O(N__16539),
            .I(N__16531));
    Span4Mux_v I__3828 (
            .O(N__16536),
            .I(N__16528));
    Span4Mux_h I__3827 (
            .O(N__16531),
            .I(N__16525));
    Odrv4 I__3826 (
            .O(N__16528),
            .I(charx_if_generate_plus_mult1_un75_sum));
    Odrv4 I__3825 (
            .O(N__16525),
            .I(charx_if_generate_plus_mult1_un75_sum));
    CascadeMux I__3824 (
            .O(N__16520),
            .I(N__16517));
    InMux I__3823 (
            .O(N__16517),
            .I(N__16502));
    InMux I__3822 (
            .O(N__16516),
            .I(N__16502));
    InMux I__3821 (
            .O(N__16515),
            .I(N__16502));
    InMux I__3820 (
            .O(N__16514),
            .I(N__16502));
    InMux I__3819 (
            .O(N__16513),
            .I(N__16502));
    LocalMux I__3818 (
            .O(N__16502),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0));
    InMux I__3817 (
            .O(N__16499),
            .I(N__16496));
    LocalMux I__3816 (
            .O(N__16496),
            .I(N__16492));
    CascadeMux I__3815 (
            .O(N__16495),
            .I(N__16487));
    Span4Mux_h I__3814 (
            .O(N__16492),
            .I(N__16482));
    InMux I__3813 (
            .O(N__16491),
            .I(N__16471));
    InMux I__3812 (
            .O(N__16490),
            .I(N__16471));
    InMux I__3811 (
            .O(N__16487),
            .I(N__16471));
    InMux I__3810 (
            .O(N__16486),
            .I(N__16471));
    InMux I__3809 (
            .O(N__16485),
            .I(N__16471));
    Odrv4 I__3808 (
            .O(N__16482),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1));
    LocalMux I__3807 (
            .O(N__16471),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1));
    CascadeMux I__3806 (
            .O(N__16466),
            .I(N__16463));
    InMux I__3805 (
            .O(N__16463),
            .I(N__16460));
    LocalMux I__3804 (
            .O(N__16460),
            .I(N__16457));
    Odrv4 I__3803 (
            .O(N__16457),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0));
    InMux I__3802 (
            .O(N__16454),
            .I(N__16451));
    LocalMux I__3801 (
            .O(N__16451),
            .I(N__16448));
    Span4Mux_v I__3800 (
            .O(N__16448),
            .I(N__16443));
    CascadeMux I__3799 (
            .O(N__16447),
            .I(N__16440));
    InMux I__3798 (
            .O(N__16446),
            .I(N__16436));
    Span4Mux_v I__3797 (
            .O(N__16443),
            .I(N__16433));
    InMux I__3796 (
            .O(N__16440),
            .I(N__16430));
    InMux I__3795 (
            .O(N__16439),
            .I(N__16427));
    LocalMux I__3794 (
            .O(N__16436),
            .I(N__16424));
    Sp12to4 I__3793 (
            .O(N__16433),
            .I(N__16419));
    LocalMux I__3792 (
            .O(N__16430),
            .I(N__16419));
    LocalMux I__3791 (
            .O(N__16427),
            .I(N__16416));
    Span4Mux_h I__3790 (
            .O(N__16424),
            .I(N__16413));
    Span12Mux_s6_h I__3789 (
            .O(N__16419),
            .I(N__16410));
    Odrv12 I__3788 (
            .O(N__16416),
            .I(charx_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3787 (
            .O(N__16413),
            .I(charx_if_generate_plus_mult1_un68_sum));
    Odrv12 I__3786 (
            .O(N__16410),
            .I(charx_if_generate_plus_mult1_un68_sum));
    InMux I__3785 (
            .O(N__16403),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__3784 (
            .O(N__16400),
            .I(N__16396));
    InMux I__3783 (
            .O(N__16399),
            .I(N__16393));
    LocalMux I__3782 (
            .O(N__16396),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0));
    LocalMux I__3781 (
            .O(N__16393),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0));
    CascadeMux I__3780 (
            .O(N__16388),
            .I(N__16385));
    InMux I__3779 (
            .O(N__16385),
            .I(N__16382));
    LocalMux I__3778 (
            .O(N__16382),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7));
    InMux I__3777 (
            .O(N__16379),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__3776 (
            .O(N__16376),
            .I(N__16373));
    LocalMux I__3775 (
            .O(N__16373),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0));
    CascadeMux I__3774 (
            .O(N__16370),
            .I(N__16366));
    CascadeMux I__3773 (
            .O(N__16369),
            .I(N__16363));
    InMux I__3772 (
            .O(N__16366),
            .I(N__16358));
    InMux I__3771 (
            .O(N__16363),
            .I(N__16358));
    LocalMux I__3770 (
            .O(N__16358),
            .I(charx_if_generate_plus_mult1_un61_sum_i_5));
    InMux I__3769 (
            .O(N__16355),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__3768 (
            .O(N__16352),
            .I(N__16349));
    LocalMux I__3767 (
            .O(N__16349),
            .I(charx_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__3766 (
            .O(N__16346),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__3765 (
            .O(N__16343),
            .I(N__16340));
    LocalMux I__3764 (
            .O(N__16340),
            .I(N__16336));
    InMux I__3763 (
            .O(N__16339),
            .I(N__16333));
    Span4Mux_v I__3762 (
            .O(N__16336),
            .I(N__16328));
    LocalMux I__3761 (
            .O(N__16333),
            .I(N__16328));
    Span4Mux_h I__3760 (
            .O(N__16328),
            .I(N__16322));
    InMux I__3759 (
            .O(N__16327),
            .I(N__16319));
    InMux I__3758 (
            .O(N__16326),
            .I(N__16316));
    CascadeMux I__3757 (
            .O(N__16325),
            .I(N__16313));
    Sp12to4 I__3756 (
            .O(N__16322),
            .I(N__16306));
    LocalMux I__3755 (
            .O(N__16319),
            .I(N__16306));
    LocalMux I__3754 (
            .O(N__16316),
            .I(N__16306));
    InMux I__3753 (
            .O(N__16313),
            .I(N__16303));
    Span12Mux_s11_v I__3752 (
            .O(N__16306),
            .I(N__16300));
    LocalMux I__3751 (
            .O(N__16303),
            .I(chessboardpixel_un152_pixel_24));
    Odrv12 I__3750 (
            .O(N__16300),
            .I(chessboardpixel_un152_pixel_24));
    InMux I__3749 (
            .O(N__16295),
            .I(N__16292));
    LocalMux I__3748 (
            .O(N__16292),
            .I(charx_if_generate_plus_mult1_un61_sum_i));
    InMux I__3747 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__3746 (
            .O(N__16286),
            .I(N__16283));
    Odrv4 I__3745 (
            .O(N__16283),
            .I(charx_if_generate_plus_mult1_un68_sum_i));
    InMux I__3744 (
            .O(N__16280),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__3743 (
            .O(N__16277),
            .I(N__16274));
    LocalMux I__3742 (
            .O(N__16274),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0));
    InMux I__3741 (
            .O(N__16271),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__3740 (
            .O(N__16268),
            .I(N__16262));
    InMux I__3739 (
            .O(N__16267),
            .I(N__16262));
    LocalMux I__3738 (
            .O(N__16262),
            .I(N__16259));
    Span4Mux_v I__3737 (
            .O(N__16259),
            .I(N__16256));
    Odrv4 I__3736 (
            .O(N__16256),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2));
    CascadeMux I__3735 (
            .O(N__16253),
            .I(N__16250));
    InMux I__3734 (
            .O(N__16250),
            .I(N__16244));
    InMux I__3733 (
            .O(N__16249),
            .I(N__16244));
    LocalMux I__3732 (
            .O(N__16244),
            .I(N__16240));
    InMux I__3731 (
            .O(N__16243),
            .I(N__16237));
    Span4Mux_s2_h I__3730 (
            .O(N__16240),
            .I(N__16234));
    LocalMux I__3729 (
            .O(N__16237),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    Odrv4 I__3728 (
            .O(N__16234),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3));
    CascadeMux I__3727 (
            .O(N__16229),
            .I(N__16226));
    InMux I__3726 (
            .O(N__16226),
            .I(N__16223));
    LocalMux I__3725 (
            .O(N__16223),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6));
    InMux I__3724 (
            .O(N__16220),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__3723 (
            .O(N__16217),
            .I(N__16213));
    InMux I__3722 (
            .O(N__16216),
            .I(N__16210));
    LocalMux I__3721 (
            .O(N__16213),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7));
    LocalMux I__3720 (
            .O(N__16210),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7));
    CascadeMux I__3719 (
            .O(N__16205),
            .I(N__16202));
    InMux I__3718 (
            .O(N__16202),
            .I(N__16199));
    LocalMux I__3717 (
            .O(N__16199),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3));
    InMux I__3716 (
            .O(N__16196),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__3715 (
            .O(N__16193),
            .I(N__16190));
    LocalMux I__3714 (
            .O(N__16190),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5));
    CascadeMux I__3713 (
            .O(N__16187),
            .I(N__16183));
    CascadeMux I__3712 (
            .O(N__16186),
            .I(N__16180));
    InMux I__3711 (
            .O(N__16183),
            .I(N__16175));
    InMux I__3710 (
            .O(N__16180),
            .I(N__16175));
    LocalMux I__3709 (
            .O(N__16175),
            .I(charx_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__3708 (
            .O(N__16172),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__3707 (
            .O(N__16169),
            .I(N__16166));
    LocalMux I__3706 (
            .O(N__16166),
            .I(charx_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__3705 (
            .O(N__16163),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__3704 (
            .O(N__16160),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_));
    InMux I__3703 (
            .O(N__16157),
            .I(N__16152));
    InMux I__3702 (
            .O(N__16156),
            .I(N__16149));
    InMux I__3701 (
            .O(N__16155),
            .I(N__16146));
    LocalMux I__3700 (
            .O(N__16152),
            .I(N__16140));
    LocalMux I__3699 (
            .O(N__16149),
            .I(N__16140));
    LocalMux I__3698 (
            .O(N__16146),
            .I(N__16137));
    InMux I__3697 (
            .O(N__16145),
            .I(N__16132));
    Span4Mux_v I__3696 (
            .O(N__16140),
            .I(N__16126));
    Span4Mux_v I__3695 (
            .O(N__16137),
            .I(N__16126));
    InMux I__3694 (
            .O(N__16136),
            .I(N__16123));
    InMux I__3693 (
            .O(N__16135),
            .I(N__16120));
    LocalMux I__3692 (
            .O(N__16132),
            .I(N__16117));
    InMux I__3691 (
            .O(N__16131),
            .I(N__16114));
    Sp12to4 I__3690 (
            .O(N__16126),
            .I(N__16109));
    LocalMux I__3689 (
            .O(N__16123),
            .I(N__16109));
    LocalMux I__3688 (
            .O(N__16120),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__3687 (
            .O(N__16117),
            .I(charx_if_generate_plus_mult1_un54_sum));
    LocalMux I__3686 (
            .O(N__16114),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv12 I__3685 (
            .O(N__16109),
            .I(charx_if_generate_plus_mult1_un54_sum));
    InMux I__3684 (
            .O(N__16100),
            .I(N__16097));
    LocalMux I__3683 (
            .O(N__16097),
            .I(charx_if_generate_plus_mult1_un54_sum_i));
    InMux I__3682 (
            .O(N__16094),
            .I(N__16091));
    LocalMux I__3681 (
            .O(N__16091),
            .I(un5_rowlto2_i));
    CascadeMux I__3680 (
            .O(N__16088),
            .I(N__16075));
    CascadeMux I__3679 (
            .O(N__16087),
            .I(N__16072));
    CascadeMux I__3678 (
            .O(N__16086),
            .I(N__16067));
    CascadeMux I__3677 (
            .O(N__16085),
            .I(N__16062));
    CascadeMux I__3676 (
            .O(N__16084),
            .I(N__16045));
    CascadeMux I__3675 (
            .O(N__16083),
            .I(N__16042));
    CascadeMux I__3674 (
            .O(N__16082),
            .I(N__16039));
    InMux I__3673 (
            .O(N__16081),
            .I(N__16026));
    InMux I__3672 (
            .O(N__16080),
            .I(N__16026));
    InMux I__3671 (
            .O(N__16079),
            .I(N__16026));
    InMux I__3670 (
            .O(N__16078),
            .I(N__16026));
    InMux I__3669 (
            .O(N__16075),
            .I(N__16019));
    InMux I__3668 (
            .O(N__16072),
            .I(N__16019));
    InMux I__3667 (
            .O(N__16071),
            .I(N__16019));
    InMux I__3666 (
            .O(N__16070),
            .I(N__16004));
    InMux I__3665 (
            .O(N__16067),
            .I(N__16004));
    InMux I__3664 (
            .O(N__16066),
            .I(N__15994));
    InMux I__3663 (
            .O(N__16065),
            .I(N__15994));
    InMux I__3662 (
            .O(N__16062),
            .I(N__15994));
    InMux I__3661 (
            .O(N__16061),
            .I(N__15994));
    InMux I__3660 (
            .O(N__16060),
            .I(N__15981));
    InMux I__3659 (
            .O(N__16059),
            .I(N__15981));
    InMux I__3658 (
            .O(N__16058),
            .I(N__15981));
    InMux I__3657 (
            .O(N__16057),
            .I(N__15981));
    InMux I__3656 (
            .O(N__16056),
            .I(N__15981));
    InMux I__3655 (
            .O(N__16055),
            .I(N__15981));
    InMux I__3654 (
            .O(N__16054),
            .I(N__15978));
    InMux I__3653 (
            .O(N__16053),
            .I(N__15967));
    InMux I__3652 (
            .O(N__16052),
            .I(N__15967));
    InMux I__3651 (
            .O(N__16051),
            .I(N__15967));
    InMux I__3650 (
            .O(N__16050),
            .I(N__15967));
    InMux I__3649 (
            .O(N__16049),
            .I(N__15967));
    InMux I__3648 (
            .O(N__16048),
            .I(N__15956));
    InMux I__3647 (
            .O(N__16045),
            .I(N__15956));
    InMux I__3646 (
            .O(N__16042),
            .I(N__15956));
    InMux I__3645 (
            .O(N__16039),
            .I(N__15956));
    InMux I__3644 (
            .O(N__16038),
            .I(N__15956));
    InMux I__3643 (
            .O(N__16037),
            .I(N__15949));
    InMux I__3642 (
            .O(N__16036),
            .I(N__15949));
    InMux I__3641 (
            .O(N__16035),
            .I(N__15949));
    LocalMux I__3640 (
            .O(N__16026),
            .I(N__15946));
    LocalMux I__3639 (
            .O(N__16019),
            .I(N__15943));
    InMux I__3638 (
            .O(N__16018),
            .I(N__15936));
    InMux I__3637 (
            .O(N__16017),
            .I(N__15936));
    InMux I__3636 (
            .O(N__16016),
            .I(N__15936));
    InMux I__3635 (
            .O(N__16015),
            .I(N__15933));
    InMux I__3634 (
            .O(N__16014),
            .I(N__15930));
    InMux I__3633 (
            .O(N__16013),
            .I(N__15923));
    InMux I__3632 (
            .O(N__16012),
            .I(N__15923));
    InMux I__3631 (
            .O(N__16011),
            .I(N__15923));
    InMux I__3630 (
            .O(N__16010),
            .I(N__15918));
    InMux I__3629 (
            .O(N__16009),
            .I(N__15918));
    LocalMux I__3628 (
            .O(N__16004),
            .I(N__15915));
    InMux I__3627 (
            .O(N__16003),
            .I(N__15912));
    LocalMux I__3626 (
            .O(N__15994),
            .I(N__15907));
    LocalMux I__3625 (
            .O(N__15981),
            .I(N__15907));
    LocalMux I__3624 (
            .O(N__15978),
            .I(N__15894));
    LocalMux I__3623 (
            .O(N__15967),
            .I(N__15894));
    LocalMux I__3622 (
            .O(N__15956),
            .I(N__15894));
    LocalMux I__3621 (
            .O(N__15949),
            .I(N__15894));
    Span4Mux_s3_v I__3620 (
            .O(N__15946),
            .I(N__15894));
    Span4Mux_s3_v I__3619 (
            .O(N__15943),
            .I(N__15894));
    LocalMux I__3618 (
            .O(N__15936),
            .I(un5_rowlto2));
    LocalMux I__3617 (
            .O(N__15933),
            .I(un5_rowlto2));
    LocalMux I__3616 (
            .O(N__15930),
            .I(un5_rowlto2));
    LocalMux I__3615 (
            .O(N__15923),
            .I(un5_rowlto2));
    LocalMux I__3614 (
            .O(N__15918),
            .I(un5_rowlto2));
    Odrv4 I__3613 (
            .O(N__15915),
            .I(un5_rowlto2));
    LocalMux I__3612 (
            .O(N__15912),
            .I(un5_rowlto2));
    Odrv4 I__3611 (
            .O(N__15907),
            .I(un5_rowlto2));
    Odrv4 I__3610 (
            .O(N__15894),
            .I(un5_rowlto2));
    CascadeMux I__3609 (
            .O(N__15875),
            .I(N__15870));
    CascadeMux I__3608 (
            .O(N__15874),
            .I(N__15865));
    CascadeMux I__3607 (
            .O(N__15873),
            .I(N__15859));
    InMux I__3606 (
            .O(N__15870),
            .I(N__15843));
    InMux I__3605 (
            .O(N__15869),
            .I(N__15843));
    InMux I__3604 (
            .O(N__15868),
            .I(N__15836));
    InMux I__3603 (
            .O(N__15865),
            .I(N__15836));
    CascadeMux I__3602 (
            .O(N__15864),
            .I(N__15832));
    CascadeMux I__3601 (
            .O(N__15863),
            .I(N__15829));
    InMux I__3600 (
            .O(N__15862),
            .I(N__15825));
    InMux I__3599 (
            .O(N__15859),
            .I(N__15822));
    InMux I__3598 (
            .O(N__15858),
            .I(N__15817));
    InMux I__3597 (
            .O(N__15857),
            .I(N__15817));
    CascadeMux I__3596 (
            .O(N__15856),
            .I(N__15814));
    CascadeMux I__3595 (
            .O(N__15855),
            .I(N__15808));
    CascadeMux I__3594 (
            .O(N__15854),
            .I(N__15803));
    CascadeMux I__3593 (
            .O(N__15853),
            .I(N__15800));
    CascadeMux I__3592 (
            .O(N__15852),
            .I(N__15795));
    CascadeMux I__3591 (
            .O(N__15851),
            .I(N__15790));
    CascadeMux I__3590 (
            .O(N__15850),
            .I(N__15784));
    CascadeMux I__3589 (
            .O(N__15849),
            .I(N__15781));
    InMux I__3588 (
            .O(N__15848),
            .I(N__15778));
    LocalMux I__3587 (
            .O(N__15843),
            .I(N__15775));
    InMux I__3586 (
            .O(N__15842),
            .I(N__15770));
    InMux I__3585 (
            .O(N__15841),
            .I(N__15770));
    LocalMux I__3584 (
            .O(N__15836),
            .I(N__15767));
    InMux I__3583 (
            .O(N__15835),
            .I(N__15758));
    InMux I__3582 (
            .O(N__15832),
            .I(N__15758));
    InMux I__3581 (
            .O(N__15829),
            .I(N__15758));
    InMux I__3580 (
            .O(N__15828),
            .I(N__15758));
    LocalMux I__3579 (
            .O(N__15825),
            .I(N__15751));
    LocalMux I__3578 (
            .O(N__15822),
            .I(N__15751));
    LocalMux I__3577 (
            .O(N__15817),
            .I(N__15751));
    InMux I__3576 (
            .O(N__15814),
            .I(N__15740));
    InMux I__3575 (
            .O(N__15813),
            .I(N__15740));
    InMux I__3574 (
            .O(N__15812),
            .I(N__15740));
    InMux I__3573 (
            .O(N__15811),
            .I(N__15740));
    InMux I__3572 (
            .O(N__15808),
            .I(N__15740));
    InMux I__3571 (
            .O(N__15807),
            .I(N__15729));
    InMux I__3570 (
            .O(N__15806),
            .I(N__15729));
    InMux I__3569 (
            .O(N__15803),
            .I(N__15729));
    InMux I__3568 (
            .O(N__15800),
            .I(N__15729));
    InMux I__3567 (
            .O(N__15799),
            .I(N__15729));
    InMux I__3566 (
            .O(N__15798),
            .I(N__15718));
    InMux I__3565 (
            .O(N__15795),
            .I(N__15718));
    InMux I__3564 (
            .O(N__15794),
            .I(N__15718));
    InMux I__3563 (
            .O(N__15793),
            .I(N__15718));
    InMux I__3562 (
            .O(N__15790),
            .I(N__15718));
    InMux I__3561 (
            .O(N__15789),
            .I(N__15707));
    InMux I__3560 (
            .O(N__15788),
            .I(N__15707));
    InMux I__3559 (
            .O(N__15787),
            .I(N__15707));
    InMux I__3558 (
            .O(N__15784),
            .I(N__15707));
    InMux I__3557 (
            .O(N__15781),
            .I(N__15707));
    LocalMux I__3556 (
            .O(N__15778),
            .I(un5_rowlto0));
    Odrv12 I__3555 (
            .O(N__15775),
            .I(un5_rowlto0));
    LocalMux I__3554 (
            .O(N__15770),
            .I(un5_rowlto0));
    Odrv4 I__3553 (
            .O(N__15767),
            .I(un5_rowlto0));
    LocalMux I__3552 (
            .O(N__15758),
            .I(un5_rowlto0));
    Odrv4 I__3551 (
            .O(N__15751),
            .I(un5_rowlto0));
    LocalMux I__3550 (
            .O(N__15740),
            .I(un5_rowlto0));
    LocalMux I__3549 (
            .O(N__15729),
            .I(un5_rowlto0));
    LocalMux I__3548 (
            .O(N__15718),
            .I(un5_rowlto0));
    LocalMux I__3547 (
            .O(N__15707),
            .I(un5_rowlto0));
    InMux I__3546 (
            .O(N__15686),
            .I(N__15670));
    InMux I__3545 (
            .O(N__15685),
            .I(N__15667));
    CascadeMux I__3544 (
            .O(N__15684),
            .I(N__15650));
    InMux I__3543 (
            .O(N__15683),
            .I(N__15645));
    InMux I__3542 (
            .O(N__15682),
            .I(N__15645));
    InMux I__3541 (
            .O(N__15681),
            .I(N__15640));
    InMux I__3540 (
            .O(N__15680),
            .I(N__15640));
    InMux I__3539 (
            .O(N__15679),
            .I(N__15633));
    InMux I__3538 (
            .O(N__15678),
            .I(N__15633));
    InMux I__3537 (
            .O(N__15677),
            .I(N__15633));
    CascadeMux I__3536 (
            .O(N__15676),
            .I(N__15628));
    CascadeMux I__3535 (
            .O(N__15675),
            .I(N__15625));
    InMux I__3534 (
            .O(N__15674),
            .I(N__15619));
    InMux I__3533 (
            .O(N__15673),
            .I(N__15619));
    LocalMux I__3532 (
            .O(N__15670),
            .I(N__15614));
    LocalMux I__3531 (
            .O(N__15667),
            .I(N__15614));
    InMux I__3530 (
            .O(N__15666),
            .I(N__15609));
    InMux I__3529 (
            .O(N__15665),
            .I(N__15609));
    InMux I__3528 (
            .O(N__15664),
            .I(N__15598));
    InMux I__3527 (
            .O(N__15663),
            .I(N__15598));
    InMux I__3526 (
            .O(N__15662),
            .I(N__15598));
    InMux I__3525 (
            .O(N__15661),
            .I(N__15598));
    InMux I__3524 (
            .O(N__15660),
            .I(N__15598));
    CascadeMux I__3523 (
            .O(N__15659),
            .I(N__15595));
    CascadeMux I__3522 (
            .O(N__15658),
            .I(N__15590));
    CascadeMux I__3521 (
            .O(N__15657),
            .I(N__15584));
    InMux I__3520 (
            .O(N__15656),
            .I(N__15571));
    InMux I__3519 (
            .O(N__15655),
            .I(N__15571));
    InMux I__3518 (
            .O(N__15654),
            .I(N__15571));
    InMux I__3517 (
            .O(N__15653),
            .I(N__15571));
    InMux I__3516 (
            .O(N__15650),
            .I(N__15571));
    LocalMux I__3515 (
            .O(N__15645),
            .I(N__15568));
    LocalMux I__3514 (
            .O(N__15640),
            .I(N__15563));
    LocalMux I__3513 (
            .O(N__15633),
            .I(N__15563));
    InMux I__3512 (
            .O(N__15632),
            .I(N__15560));
    InMux I__3511 (
            .O(N__15631),
            .I(N__15551));
    InMux I__3510 (
            .O(N__15628),
            .I(N__15551));
    InMux I__3509 (
            .O(N__15625),
            .I(N__15551));
    InMux I__3508 (
            .O(N__15624),
            .I(N__15551));
    LocalMux I__3507 (
            .O(N__15619),
            .I(N__15542));
    Span4Mux_v I__3506 (
            .O(N__15614),
            .I(N__15542));
    LocalMux I__3505 (
            .O(N__15609),
            .I(N__15542));
    LocalMux I__3504 (
            .O(N__15598),
            .I(N__15542));
    InMux I__3503 (
            .O(N__15595),
            .I(N__15533));
    InMux I__3502 (
            .O(N__15594),
            .I(N__15533));
    InMux I__3501 (
            .O(N__15593),
            .I(N__15533));
    InMux I__3500 (
            .O(N__15590),
            .I(N__15533));
    InMux I__3499 (
            .O(N__15589),
            .I(N__15526));
    InMux I__3498 (
            .O(N__15588),
            .I(N__15526));
    InMux I__3497 (
            .O(N__15587),
            .I(N__15526));
    InMux I__3496 (
            .O(N__15584),
            .I(N__15519));
    InMux I__3495 (
            .O(N__15583),
            .I(N__15519));
    InMux I__3494 (
            .O(N__15582),
            .I(N__15519));
    LocalMux I__3493 (
            .O(N__15571),
            .I(un5_rowlto1));
    Odrv12 I__3492 (
            .O(N__15568),
            .I(un5_rowlto1));
    Odrv4 I__3491 (
            .O(N__15563),
            .I(un5_rowlto1));
    LocalMux I__3490 (
            .O(N__15560),
            .I(un5_rowlto1));
    LocalMux I__3489 (
            .O(N__15551),
            .I(un5_rowlto1));
    Odrv4 I__3488 (
            .O(N__15542),
            .I(un5_rowlto1));
    LocalMux I__3487 (
            .O(N__15533),
            .I(un5_rowlto1));
    LocalMux I__3486 (
            .O(N__15526),
            .I(un5_rowlto1));
    LocalMux I__3485 (
            .O(N__15519),
            .I(un5_rowlto1));
    InMux I__3484 (
            .O(N__15500),
            .I(N__15482));
    InMux I__3483 (
            .O(N__15499),
            .I(N__15482));
    InMux I__3482 (
            .O(N__15498),
            .I(N__15482));
    InMux I__3481 (
            .O(N__15497),
            .I(N__15482));
    InMux I__3480 (
            .O(N__15496),
            .I(N__15462));
    InMux I__3479 (
            .O(N__15495),
            .I(N__15462));
    InMux I__3478 (
            .O(N__15494),
            .I(N__15453));
    InMux I__3477 (
            .O(N__15493),
            .I(N__15453));
    InMux I__3476 (
            .O(N__15492),
            .I(N__15453));
    InMux I__3475 (
            .O(N__15491),
            .I(N__15453));
    LocalMux I__3474 (
            .O(N__15482),
            .I(N__15450));
    InMux I__3473 (
            .O(N__15481),
            .I(N__15439));
    InMux I__3472 (
            .O(N__15480),
            .I(N__15439));
    InMux I__3471 (
            .O(N__15479),
            .I(N__15439));
    InMux I__3470 (
            .O(N__15478),
            .I(N__15439));
    InMux I__3469 (
            .O(N__15477),
            .I(N__15439));
    InMux I__3468 (
            .O(N__15476),
            .I(N__15434));
    InMux I__3467 (
            .O(N__15475),
            .I(N__15434));
    InMux I__3466 (
            .O(N__15474),
            .I(N__15427));
    InMux I__3465 (
            .O(N__15473),
            .I(N__15427));
    InMux I__3464 (
            .O(N__15472),
            .I(N__15427));
    InMux I__3463 (
            .O(N__15471),
            .I(N__15420));
    InMux I__3462 (
            .O(N__15470),
            .I(N__15420));
    InMux I__3461 (
            .O(N__15469),
            .I(N__15420));
    InMux I__3460 (
            .O(N__15468),
            .I(N__15415));
    InMux I__3459 (
            .O(N__15467),
            .I(N__15415));
    LocalMux I__3458 (
            .O(N__15462),
            .I(N__15406));
    LocalMux I__3457 (
            .O(N__15453),
            .I(N__15406));
    Span4Mux_v I__3456 (
            .O(N__15450),
            .I(N__15403));
    LocalMux I__3455 (
            .O(N__15439),
            .I(N__15396));
    LocalMux I__3454 (
            .O(N__15434),
            .I(N__15396));
    LocalMux I__3453 (
            .O(N__15427),
            .I(N__15396));
    LocalMux I__3452 (
            .O(N__15420),
            .I(N__15391));
    LocalMux I__3451 (
            .O(N__15415),
            .I(N__15391));
    InMux I__3450 (
            .O(N__15414),
            .I(N__15386));
    InMux I__3449 (
            .O(N__15413),
            .I(N__15386));
    InMux I__3448 (
            .O(N__15412),
            .I(N__15378));
    InMux I__3447 (
            .O(N__15411),
            .I(N__15378));
    Span4Mux_v I__3446 (
            .O(N__15406),
            .I(N__15373));
    Span4Mux_v I__3445 (
            .O(N__15403),
            .I(N__15373));
    Span4Mux_v I__3444 (
            .O(N__15396),
            .I(N__15366));
    Span4Mux_v I__3443 (
            .O(N__15391),
            .I(N__15366));
    LocalMux I__3442 (
            .O(N__15386),
            .I(N__15366));
    InMux I__3441 (
            .O(N__15385),
            .I(N__15363));
    InMux I__3440 (
            .O(N__15384),
            .I(N__15358));
    InMux I__3439 (
            .O(N__15383),
            .I(N__15358));
    LocalMux I__3438 (
            .O(N__15378),
            .I(un5_rowlto3));
    Odrv4 I__3437 (
            .O(N__15373),
            .I(un5_rowlto3));
    Odrv4 I__3436 (
            .O(N__15366),
            .I(un5_rowlto3));
    LocalMux I__3435 (
            .O(N__15363),
            .I(un5_rowlto3));
    LocalMux I__3434 (
            .O(N__15358),
            .I(un5_rowlto3));
    InMux I__3433 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__3432 (
            .O(N__15344),
            .I(un116_pixel_2_amZ0Z_1));
    CascadeMux I__3431 (
            .O(N__15341),
            .I(N__15338));
    InMux I__3430 (
            .O(N__15338),
            .I(N__15335));
    LocalMux I__3429 (
            .O(N__15335),
            .I(N__15332));
    Span4Mux_s2_h I__3428 (
            .O(N__15332),
            .I(N__15329));
    Odrv4 I__3427 (
            .O(N__15329),
            .I(charx_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__3426 (
            .O(N__15326),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__3425 (
            .O(N__15323),
            .I(N__15320));
    LocalMux I__3424 (
            .O(N__15320),
            .I(N__15317));
    Span4Mux_s2_h I__3423 (
            .O(N__15317),
            .I(N__15314));
    Odrv4 I__3422 (
            .O(N__15314),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1));
    InMux I__3421 (
            .O(N__15311),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__3420 (
            .O(N__15308),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__3419 (
            .O(N__15305),
            .I(N__15302));
    LocalMux I__3418 (
            .O(N__15302),
            .I(N__15299));
    Span4Mux_v I__3417 (
            .O(N__15299),
            .I(N__15296));
    Odrv4 I__3416 (
            .O(N__15296),
            .I(charx_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__3415 (
            .O(N__15293),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__3414 (
            .O(N__15290),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_));
    InMux I__3413 (
            .O(N__15287),
            .I(N__15281));
    InMux I__3412 (
            .O(N__15286),
            .I(N__15276));
    InMux I__3411 (
            .O(N__15285),
            .I(N__15273));
    InMux I__3410 (
            .O(N__15284),
            .I(N__15270));
    LocalMux I__3409 (
            .O(N__15281),
            .I(N__15267));
    InMux I__3408 (
            .O(N__15280),
            .I(N__15264));
    InMux I__3407 (
            .O(N__15279),
            .I(N__15261));
    LocalMux I__3406 (
            .O(N__15276),
            .I(N__15256));
    LocalMux I__3405 (
            .O(N__15273),
            .I(N__15256));
    LocalMux I__3404 (
            .O(N__15270),
            .I(N__15253));
    Span4Mux_h I__3403 (
            .O(N__15267),
            .I(N__15250));
    LocalMux I__3402 (
            .O(N__15264),
            .I(charx_if_generate_plus_mult1_un47_sum));
    LocalMux I__3401 (
            .O(N__15261),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3400 (
            .O(N__15256),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv12 I__3399 (
            .O(N__15253),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__3398 (
            .O(N__15250),
            .I(charx_if_generate_plus_mult1_un47_sum));
    InMux I__3397 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__3396 (
            .O(N__15236),
            .I(charx_if_generate_plus_mult1_un47_sum_i));
    CascadeMux I__3395 (
            .O(N__15233),
            .I(N__15230));
    InMux I__3394 (
            .O(N__15230),
            .I(N__15227));
    LocalMux I__3393 (
            .O(N__15227),
            .I(N__15224));
    Span4Mux_h I__3392 (
            .O(N__15224),
            .I(N__15221));
    Odrv4 I__3391 (
            .O(N__15221),
            .I(N_302_i_0));
    CascadeMux I__3390 (
            .O(N__15218),
            .I(beamY_RNITQPUS72Z0Z_0_cascade_));
    InMux I__3389 (
            .O(N__15215),
            .I(N__15212));
    LocalMux I__3388 (
            .O(N__15212),
            .I(un116_pixel_3_1_0));
    CascadeMux I__3387 (
            .O(N__15209),
            .I(N__15206));
    InMux I__3386 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__3385 (
            .O(N__15203),
            .I(beamY_RNI6B7UAL1Z0Z_1));
    InMux I__3384 (
            .O(N__15200),
            .I(N__15197));
    LocalMux I__3383 (
            .O(N__15197),
            .I(N__15194));
    Span4Mux_h I__3382 (
            .O(N__15194),
            .I(N__15190));
    InMux I__3381 (
            .O(N__15193),
            .I(N__15187));
    Odrv4 I__3380 (
            .O(N__15190),
            .I(m31));
    LocalMux I__3379 (
            .O(N__15187),
            .I(m31));
    InMux I__3378 (
            .O(N__15182),
            .I(N__15179));
    LocalMux I__3377 (
            .O(N__15179),
            .I(un116_pixel_4_1Z0Z_0));
    InMux I__3376 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__3375 (
            .O(N__15173),
            .I(m38));
    InMux I__3374 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__3373 (
            .O(N__15167),
            .I(N__15157));
    InMux I__3372 (
            .O(N__15166),
            .I(N__15154));
    CascadeMux I__3371 (
            .O(N__15165),
            .I(N__15150));
    CascadeMux I__3370 (
            .O(N__15164),
            .I(N__15147));
    CascadeMux I__3369 (
            .O(N__15163),
            .I(N__15139));
    CascadeMux I__3368 (
            .O(N__15162),
            .I(N__15134));
    CascadeMux I__3367 (
            .O(N__15161),
            .I(N__15129));
    CascadeMux I__3366 (
            .O(N__15160),
            .I(N__15124));
    Span4Mux_h I__3365 (
            .O(N__15157),
            .I(N__15119));
    LocalMux I__3364 (
            .O(N__15154),
            .I(N__15119));
    InMux I__3363 (
            .O(N__15153),
            .I(N__15110));
    InMux I__3362 (
            .O(N__15150),
            .I(N__15110));
    InMux I__3361 (
            .O(N__15147),
            .I(N__15110));
    InMux I__3360 (
            .O(N__15146),
            .I(N__15110));
    CascadeMux I__3359 (
            .O(N__15145),
            .I(N__15103));
    CascadeMux I__3358 (
            .O(N__15144),
            .I(N__15098));
    CascadeMux I__3357 (
            .O(N__15143),
            .I(N__15094));
    InMux I__3356 (
            .O(N__15142),
            .I(N__15091));
    InMux I__3355 (
            .O(N__15139),
            .I(N__15088));
    InMux I__3354 (
            .O(N__15138),
            .I(N__15085));
    InMux I__3353 (
            .O(N__15137),
            .I(N__15082));
    InMux I__3352 (
            .O(N__15134),
            .I(N__15079));
    InMux I__3351 (
            .O(N__15133),
            .I(N__15076));
    InMux I__3350 (
            .O(N__15132),
            .I(N__15073));
    InMux I__3349 (
            .O(N__15129),
            .I(N__15066));
    InMux I__3348 (
            .O(N__15128),
            .I(N__15066));
    InMux I__3347 (
            .O(N__15127),
            .I(N__15066));
    InMux I__3346 (
            .O(N__15124),
            .I(N__15063));
    Span4Mux_h I__3345 (
            .O(N__15119),
            .I(N__15058));
    LocalMux I__3344 (
            .O(N__15110),
            .I(N__15058));
    InMux I__3343 (
            .O(N__15109),
            .I(N__15053));
    InMux I__3342 (
            .O(N__15108),
            .I(N__15053));
    InMux I__3341 (
            .O(N__15107),
            .I(N__15049));
    InMux I__3340 (
            .O(N__15106),
            .I(N__15038));
    InMux I__3339 (
            .O(N__15103),
            .I(N__15038));
    InMux I__3338 (
            .O(N__15102),
            .I(N__15038));
    InMux I__3337 (
            .O(N__15101),
            .I(N__15038));
    InMux I__3336 (
            .O(N__15098),
            .I(N__15038));
    CascadeMux I__3335 (
            .O(N__15097),
            .I(N__15032));
    InMux I__3334 (
            .O(N__15094),
            .I(N__15029));
    LocalMux I__3333 (
            .O(N__15091),
            .I(N__15026));
    LocalMux I__3332 (
            .O(N__15088),
            .I(N__15019));
    LocalMux I__3331 (
            .O(N__15085),
            .I(N__15019));
    LocalMux I__3330 (
            .O(N__15082),
            .I(N__15019));
    LocalMux I__3329 (
            .O(N__15079),
            .I(N__15016));
    LocalMux I__3328 (
            .O(N__15076),
            .I(N__15013));
    LocalMux I__3327 (
            .O(N__15073),
            .I(N__15010));
    LocalMux I__3326 (
            .O(N__15066),
            .I(N__15001));
    LocalMux I__3325 (
            .O(N__15063),
            .I(N__15001));
    Span4Mux_v I__3324 (
            .O(N__15058),
            .I(N__15001));
    LocalMux I__3323 (
            .O(N__15053),
            .I(N__15001));
    InMux I__3322 (
            .O(N__15052),
            .I(N__14997));
    LocalMux I__3321 (
            .O(N__15049),
            .I(N__14994));
    LocalMux I__3320 (
            .O(N__15038),
            .I(N__14991));
    InMux I__3319 (
            .O(N__15037),
            .I(N__14988));
    InMux I__3318 (
            .O(N__15036),
            .I(N__14981));
    InMux I__3317 (
            .O(N__15035),
            .I(N__14981));
    InMux I__3316 (
            .O(N__15032),
            .I(N__14981));
    LocalMux I__3315 (
            .O(N__15029),
            .I(N__14974));
    Span4Mux_h I__3314 (
            .O(N__15026),
            .I(N__14974));
    Span4Mux_h I__3313 (
            .O(N__15019),
            .I(N__14974));
    Span4Mux_h I__3312 (
            .O(N__15016),
            .I(N__14969));
    Span4Mux_h I__3311 (
            .O(N__15013),
            .I(N__14969));
    Span4Mux_h I__3310 (
            .O(N__15010),
            .I(N__14964));
    Span4Mux_h I__3309 (
            .O(N__15001),
            .I(N__14964));
    InMux I__3308 (
            .O(N__15000),
            .I(N__14961));
    LocalMux I__3307 (
            .O(N__14997),
            .I(beamYZ0Z_0));
    Odrv4 I__3306 (
            .O(N__14994),
            .I(beamYZ0Z_0));
    Odrv4 I__3305 (
            .O(N__14991),
            .I(beamYZ0Z_0));
    LocalMux I__3304 (
            .O(N__14988),
            .I(beamYZ0Z_0));
    LocalMux I__3303 (
            .O(N__14981),
            .I(beamYZ0Z_0));
    Odrv4 I__3302 (
            .O(N__14974),
            .I(beamYZ0Z_0));
    Odrv4 I__3301 (
            .O(N__14969),
            .I(beamYZ0Z_0));
    Odrv4 I__3300 (
            .O(N__14964),
            .I(beamYZ0Z_0));
    LocalMux I__3299 (
            .O(N__14961),
            .I(beamYZ0Z_0));
    CascadeMux I__3298 (
            .O(N__14942),
            .I(m38_cascade_));
    CascadeMux I__3297 (
            .O(N__14939),
            .I(N__14931));
    InMux I__3296 (
            .O(N__14938),
            .I(N__14926));
    InMux I__3295 (
            .O(N__14937),
            .I(N__14917));
    InMux I__3294 (
            .O(N__14936),
            .I(N__14914));
    InMux I__3293 (
            .O(N__14935),
            .I(N__14909));
    InMux I__3292 (
            .O(N__14934),
            .I(N__14909));
    InMux I__3291 (
            .O(N__14931),
            .I(N__14902));
    InMux I__3290 (
            .O(N__14930),
            .I(N__14899));
    CascadeMux I__3289 (
            .O(N__14929),
            .I(N__14895));
    LocalMux I__3288 (
            .O(N__14926),
            .I(N__14892));
    InMux I__3287 (
            .O(N__14925),
            .I(N__14889));
    InMux I__3286 (
            .O(N__14924),
            .I(N__14886));
    InMux I__3285 (
            .O(N__14923),
            .I(N__14883));
    InMux I__3284 (
            .O(N__14922),
            .I(N__14880));
    InMux I__3283 (
            .O(N__14921),
            .I(N__14877));
    InMux I__3282 (
            .O(N__14920),
            .I(N__14874));
    LocalMux I__3281 (
            .O(N__14917),
            .I(N__14870));
    LocalMux I__3280 (
            .O(N__14914),
            .I(N__14865));
    LocalMux I__3279 (
            .O(N__14909),
            .I(N__14865));
    InMux I__3278 (
            .O(N__14908),
            .I(N__14862));
    InMux I__3277 (
            .O(N__14907),
            .I(N__14859));
    InMux I__3276 (
            .O(N__14906),
            .I(N__14856));
    CascadeMux I__3275 (
            .O(N__14905),
            .I(N__14851));
    LocalMux I__3274 (
            .O(N__14902),
            .I(N__14844));
    LocalMux I__3273 (
            .O(N__14899),
            .I(N__14841));
    CascadeMux I__3272 (
            .O(N__14898),
            .I(N__14838));
    InMux I__3271 (
            .O(N__14895),
            .I(N__14835));
    Span4Mux_v I__3270 (
            .O(N__14892),
            .I(N__14832));
    LocalMux I__3269 (
            .O(N__14889),
            .I(N__14825));
    LocalMux I__3268 (
            .O(N__14886),
            .I(N__14825));
    LocalMux I__3267 (
            .O(N__14883),
            .I(N__14825));
    LocalMux I__3266 (
            .O(N__14880),
            .I(N__14820));
    LocalMux I__3265 (
            .O(N__14877),
            .I(N__14820));
    LocalMux I__3264 (
            .O(N__14874),
            .I(N__14817));
    InMux I__3263 (
            .O(N__14873),
            .I(N__14814));
    Span4Mux_h I__3262 (
            .O(N__14870),
            .I(N__14803));
    Span4Mux_v I__3261 (
            .O(N__14865),
            .I(N__14803));
    LocalMux I__3260 (
            .O(N__14862),
            .I(N__14803));
    LocalMux I__3259 (
            .O(N__14859),
            .I(N__14803));
    LocalMux I__3258 (
            .O(N__14856),
            .I(N__14803));
    InMux I__3257 (
            .O(N__14855),
            .I(N__14800));
    InMux I__3256 (
            .O(N__14854),
            .I(N__14797));
    InMux I__3255 (
            .O(N__14851),
            .I(N__14794));
    InMux I__3254 (
            .O(N__14850),
            .I(N__14787));
    InMux I__3253 (
            .O(N__14849),
            .I(N__14787));
    InMux I__3252 (
            .O(N__14848),
            .I(N__14787));
    InMux I__3251 (
            .O(N__14847),
            .I(N__14784));
    Span4Mux_h I__3250 (
            .O(N__14844),
            .I(N__14779));
    Span4Mux_h I__3249 (
            .O(N__14841),
            .I(N__14779));
    InMux I__3248 (
            .O(N__14838),
            .I(N__14776));
    LocalMux I__3247 (
            .O(N__14835),
            .I(N__14769));
    Span4Mux_s2_h I__3246 (
            .O(N__14832),
            .I(N__14769));
    Span4Mux_v I__3245 (
            .O(N__14825),
            .I(N__14769));
    Span4Mux_h I__3244 (
            .O(N__14820),
            .I(N__14760));
    Span4Mux_h I__3243 (
            .O(N__14817),
            .I(N__14760));
    LocalMux I__3242 (
            .O(N__14814),
            .I(N__14760));
    Span4Mux_v I__3241 (
            .O(N__14803),
            .I(N__14760));
    LocalMux I__3240 (
            .O(N__14800),
            .I(beamYZ0Z_1));
    LocalMux I__3239 (
            .O(N__14797),
            .I(beamYZ0Z_1));
    LocalMux I__3238 (
            .O(N__14794),
            .I(beamYZ0Z_1));
    LocalMux I__3237 (
            .O(N__14787),
            .I(beamYZ0Z_1));
    LocalMux I__3236 (
            .O(N__14784),
            .I(beamYZ0Z_1));
    Odrv4 I__3235 (
            .O(N__14779),
            .I(beamYZ0Z_1));
    LocalMux I__3234 (
            .O(N__14776),
            .I(beamYZ0Z_1));
    Odrv4 I__3233 (
            .O(N__14769),
            .I(beamYZ0Z_1));
    Odrv4 I__3232 (
            .O(N__14760),
            .I(beamYZ0Z_1));
    CascadeMux I__3231 (
            .O(N__14741),
            .I(un116_pixel_6_1_1_cascade_));
    InMux I__3230 (
            .O(N__14738),
            .I(N__14735));
    LocalMux I__3229 (
            .O(N__14735),
            .I(N__14732));
    Odrv4 I__3228 (
            .O(N__14732),
            .I(N_17));
    InMux I__3227 (
            .O(N__14729),
            .I(N__14726));
    LocalMux I__3226 (
            .O(N__14726),
            .I(N__14719));
    InMux I__3225 (
            .O(N__14725),
            .I(N__14714));
    InMux I__3224 (
            .O(N__14724),
            .I(N__14714));
    InMux I__3223 (
            .O(N__14723),
            .I(N__14711));
    InMux I__3222 (
            .O(N__14722),
            .I(N__14708));
    Span4Mux_h I__3221 (
            .O(N__14719),
            .I(N__14703));
    LocalMux I__3220 (
            .O(N__14714),
            .I(N__14703));
    LocalMux I__3219 (
            .O(N__14711),
            .I(N__14700));
    LocalMux I__3218 (
            .O(N__14708),
            .I(N_321));
    Odrv4 I__3217 (
            .O(N__14703),
            .I(N_321));
    Odrv4 I__3216 (
            .O(N__14700),
            .I(N_321));
    InMux I__3215 (
            .O(N__14693),
            .I(N__14690));
    LocalMux I__3214 (
            .O(N__14690),
            .I(un116_pixel_2_bmZ0Z_1));
    CascadeMux I__3213 (
            .O(N__14687),
            .I(beamY_RNI4NRC8D1Z0Z_0_cascade_));
    InMux I__3212 (
            .O(N__14684),
            .I(N__14681));
    LocalMux I__3211 (
            .O(N__14681),
            .I(beamY_RNII25UDD3Z0Z_0));
    InMux I__3210 (
            .O(N__14678),
            .I(N__14675));
    LocalMux I__3209 (
            .O(N__14675),
            .I(N_14));
    CascadeMux I__3208 (
            .O(N__14672),
            .I(un116_pixel_2_ns_1_6_cascade_));
    InMux I__3207 (
            .O(N__14669),
            .I(N__14666));
    LocalMux I__3206 (
            .O(N__14666),
            .I(beamY_RNIH01F2SZ0Z_0));
    InMux I__3205 (
            .O(N__14663),
            .I(N__14660));
    LocalMux I__3204 (
            .O(N__14660),
            .I(un116_pixel_2_ns_1Z0Z_5));
    CascadeMux I__3203 (
            .O(N__14657),
            .I(N_276_0_cascade_));
    InMux I__3202 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__3201 (
            .O(N__14651),
            .I(N__14648));
    Odrv4 I__3200 (
            .O(N__14648),
            .I(beamY_RNII25UDD3_3Z0Z_0));
    InMux I__3199 (
            .O(N__14645),
            .I(N__14642));
    LocalMux I__3198 (
            .O(N__14642),
            .I(m7));
    CascadeMux I__3197 (
            .O(N__14639),
            .I(m7_cascade_));
    InMux I__3196 (
            .O(N__14636),
            .I(N__14633));
    LocalMux I__3195 (
            .O(N__14633),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3));
    InMux I__3194 (
            .O(N__14630),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2));
    CascadeMux I__3193 (
            .O(N__14627),
            .I(N__14624));
    InMux I__3192 (
            .O(N__14624),
            .I(N__14621));
    LocalMux I__3191 (
            .O(N__14621),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0));
    InMux I__3190 (
            .O(N__14618),
            .I(N__14609));
    InMux I__3189 (
            .O(N__14617),
            .I(N__14609));
    InMux I__3188 (
            .O(N__14616),
            .I(N__14609));
    LocalMux I__3187 (
            .O(N__14609),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO));
    InMux I__3186 (
            .O(N__14606),
            .I(N__14603));
    LocalMux I__3185 (
            .O(N__14603),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO));
    CascadeMux I__3184 (
            .O(N__14600),
            .I(N__14596));
    CascadeMux I__3183 (
            .O(N__14599),
            .I(N__14593));
    InMux I__3182 (
            .O(N__14596),
            .I(N__14588));
    InMux I__3181 (
            .O(N__14593),
            .I(N__14588));
    LocalMux I__3180 (
            .O(N__14588),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803));
    InMux I__3179 (
            .O(N__14585),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4));
    InMux I__3178 (
            .O(N__14582),
            .I(N__14575));
    InMux I__3177 (
            .O(N__14581),
            .I(N__14572));
    InMux I__3176 (
            .O(N__14580),
            .I(N__14565));
    InMux I__3175 (
            .O(N__14579),
            .I(N__14565));
    InMux I__3174 (
            .O(N__14578),
            .I(N__14565));
    LocalMux I__3173 (
            .O(N__14575),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    LocalMux I__3172 (
            .O(N__14572),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    LocalMux I__3171 (
            .O(N__14565),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3));
    InMux I__3170 (
            .O(N__14558),
            .I(N__14555));
    LocalMux I__3169 (
            .O(N__14555),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3));
    CascadeMux I__3168 (
            .O(N__14552),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_));
    CascadeMux I__3167 (
            .O(N__14549),
            .I(N__14546));
    InMux I__3166 (
            .O(N__14546),
            .I(N__14540));
    InMux I__3165 (
            .O(N__14545),
            .I(N__14540));
    LocalMux I__3164 (
            .O(N__14540),
            .I(un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1));
    InMux I__3163 (
            .O(N__14537),
            .I(N__14528));
    InMux I__3162 (
            .O(N__14536),
            .I(N__14525));
    InMux I__3161 (
            .O(N__14535),
            .I(N__14518));
    InMux I__3160 (
            .O(N__14534),
            .I(N__14518));
    InMux I__3159 (
            .O(N__14533),
            .I(N__14518));
    InMux I__3158 (
            .O(N__14532),
            .I(N__14513));
    InMux I__3157 (
            .O(N__14531),
            .I(N__14513));
    LocalMux I__3156 (
            .O(N__14528),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__3155 (
            .O(N__14525),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__3154 (
            .O(N__14518),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__3153 (
            .O(N__14513),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    InMux I__3152 (
            .O(N__14504),
            .I(N__14494));
    InMux I__3151 (
            .O(N__14503),
            .I(N__14487));
    InMux I__3150 (
            .O(N__14502),
            .I(N__14487));
    InMux I__3149 (
            .O(N__14501),
            .I(N__14487));
    InMux I__3148 (
            .O(N__14500),
            .I(N__14484));
    InMux I__3147 (
            .O(N__14499),
            .I(N__14481));
    InMux I__3146 (
            .O(N__14498),
            .I(N__14478));
    CascadeMux I__3145 (
            .O(N__14497),
            .I(N__14471));
    LocalMux I__3144 (
            .O(N__14494),
            .I(N__14466));
    LocalMux I__3143 (
            .O(N__14487),
            .I(N__14466));
    LocalMux I__3142 (
            .O(N__14484),
            .I(N__14461));
    LocalMux I__3141 (
            .O(N__14481),
            .I(N__14461));
    LocalMux I__3140 (
            .O(N__14478),
            .I(N__14458));
    InMux I__3139 (
            .O(N__14477),
            .I(N__14455));
    CascadeMux I__3138 (
            .O(N__14476),
            .I(N__14452));
    InMux I__3137 (
            .O(N__14475),
            .I(N__14447));
    InMux I__3136 (
            .O(N__14474),
            .I(N__14447));
    InMux I__3135 (
            .O(N__14471),
            .I(N__14444));
    Span12Mux_s6_h I__3134 (
            .O(N__14466),
            .I(N__14441));
    Span4Mux_v I__3133 (
            .O(N__14461),
            .I(N__14438));
    Span12Mux_s10_v I__3132 (
            .O(N__14458),
            .I(N__14435));
    LocalMux I__3131 (
            .O(N__14455),
            .I(N__14432));
    InMux I__3130 (
            .O(N__14452),
            .I(N__14429));
    LocalMux I__3129 (
            .O(N__14447),
            .I(beamXZ0Z_0));
    LocalMux I__3128 (
            .O(N__14444),
            .I(beamXZ0Z_0));
    Odrv12 I__3127 (
            .O(N__14441),
            .I(beamXZ0Z_0));
    Odrv4 I__3126 (
            .O(N__14438),
            .I(beamXZ0Z_0));
    Odrv12 I__3125 (
            .O(N__14435),
            .I(beamXZ0Z_0));
    Odrv4 I__3124 (
            .O(N__14432),
            .I(beamXZ0Z_0));
    LocalMux I__3123 (
            .O(N__14429),
            .I(beamXZ0Z_0));
    InMux I__3122 (
            .O(N__14414),
            .I(N__14409));
    InMux I__3121 (
            .O(N__14413),
            .I(N__14406));
    InMux I__3120 (
            .O(N__14412),
            .I(N__14403));
    LocalMux I__3119 (
            .O(N__14409),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__3118 (
            .O(N__14406),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    LocalMux I__3117 (
            .O(N__14403),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1));
    CascadeMux I__3116 (
            .O(N__14396),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_));
    InMux I__3115 (
            .O(N__14393),
            .I(N__14390));
    LocalMux I__3114 (
            .O(N__14390),
            .I(un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1));
    CascadeMux I__3113 (
            .O(N__14387),
            .I(m15_cascade_));
    InMux I__3112 (
            .O(N__14384),
            .I(N__14377));
    InMux I__3111 (
            .O(N__14383),
            .I(N__14372));
    InMux I__3110 (
            .O(N__14382),
            .I(N__14372));
    InMux I__3109 (
            .O(N__14381),
            .I(N__14369));
    InMux I__3108 (
            .O(N__14380),
            .I(N__14366));
    LocalMux I__3107 (
            .O(N__14377),
            .I(N__14363));
    LocalMux I__3106 (
            .O(N__14372),
            .I(N__14360));
    LocalMux I__3105 (
            .O(N__14369),
            .I(un114_pixel_0_1__N_6_mux));
    LocalMux I__3104 (
            .O(N__14366),
            .I(un114_pixel_0_1__N_6_mux));
    Odrv4 I__3103 (
            .O(N__14363),
            .I(un114_pixel_0_1__N_6_mux));
    Odrv4 I__3102 (
            .O(N__14360),
            .I(un114_pixel_0_1__N_6_mux));
    InMux I__3101 (
            .O(N__14351),
            .I(N__14347));
    InMux I__3100 (
            .O(N__14350),
            .I(N__14342));
    LocalMux I__3099 (
            .O(N__14347),
            .I(N__14339));
    InMux I__3098 (
            .O(N__14346),
            .I(N__14336));
    CascadeMux I__3097 (
            .O(N__14345),
            .I(N__14331));
    LocalMux I__3096 (
            .O(N__14342),
            .I(N__14326));
    Span4Mux_v I__3095 (
            .O(N__14339),
            .I(N__14321));
    LocalMux I__3094 (
            .O(N__14336),
            .I(N__14321));
    InMux I__3093 (
            .O(N__14335),
            .I(N__14316));
    InMux I__3092 (
            .O(N__14334),
            .I(N__14316));
    InMux I__3091 (
            .O(N__14331),
            .I(N__14313));
    InMux I__3090 (
            .O(N__14330),
            .I(N__14310));
    InMux I__3089 (
            .O(N__14329),
            .I(N__14307));
    Span4Mux_h I__3088 (
            .O(N__14326),
            .I(N__14304));
    Span4Mux_h I__3087 (
            .O(N__14321),
            .I(N__14301));
    LocalMux I__3086 (
            .O(N__14316),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__3085 (
            .O(N__14313),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__3084 (
            .O(N__14310),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__3083 (
            .O(N__14307),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3082 (
            .O(N__14304),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__3081 (
            .O(N__14301),
            .I(charx_if_generate_plus_mult1_un40_sum));
    InMux I__3080 (
            .O(N__14288),
            .I(N__14285));
    LocalMux I__3079 (
            .O(N__14285),
            .I(charx_if_generate_plus_mult1_un40_sum_i));
    InMux I__3078 (
            .O(N__14282),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1));
    InMux I__3077 (
            .O(N__14279),
            .I(N__14267));
    InMux I__3076 (
            .O(N__14278),
            .I(N__14262));
    CascadeMux I__3075 (
            .O(N__14277),
            .I(N__14259));
    CascadeMux I__3074 (
            .O(N__14276),
            .I(N__14256));
    CascadeMux I__3073 (
            .O(N__14275),
            .I(N__14253));
    InMux I__3072 (
            .O(N__14274),
            .I(N__14247));
    InMux I__3071 (
            .O(N__14273),
            .I(N__14242));
    InMux I__3070 (
            .O(N__14272),
            .I(N__14242));
    CascadeMux I__3069 (
            .O(N__14271),
            .I(N__14239));
    InMux I__3068 (
            .O(N__14270),
            .I(N__14233));
    LocalMux I__3067 (
            .O(N__14267),
            .I(N__14230));
    InMux I__3066 (
            .O(N__14266),
            .I(N__14227));
    CascadeMux I__3065 (
            .O(N__14265),
            .I(N__14223));
    LocalMux I__3064 (
            .O(N__14262),
            .I(N__14218));
    InMux I__3063 (
            .O(N__14259),
            .I(N__14215));
    InMux I__3062 (
            .O(N__14256),
            .I(N__14210));
    InMux I__3061 (
            .O(N__14253),
            .I(N__14210));
    CascadeMux I__3060 (
            .O(N__14252),
            .I(N__14207));
    CascadeMux I__3059 (
            .O(N__14251),
            .I(N__14204));
    IoInMux I__3058 (
            .O(N__14250),
            .I(N__14201));
    LocalMux I__3057 (
            .O(N__14247),
            .I(N__14196));
    LocalMux I__3056 (
            .O(N__14242),
            .I(N__14196));
    InMux I__3055 (
            .O(N__14239),
            .I(N__14191));
    InMux I__3054 (
            .O(N__14238),
            .I(N__14191));
    InMux I__3053 (
            .O(N__14237),
            .I(N__14188));
    InMux I__3052 (
            .O(N__14236),
            .I(N__14185));
    LocalMux I__3051 (
            .O(N__14233),
            .I(N__14181));
    Span4Mux_v I__3050 (
            .O(N__14230),
            .I(N__14176));
    LocalMux I__3049 (
            .O(N__14227),
            .I(N__14176));
    InMux I__3048 (
            .O(N__14226),
            .I(N__14173));
    InMux I__3047 (
            .O(N__14223),
            .I(N__14168));
    InMux I__3046 (
            .O(N__14222),
            .I(N__14168));
    InMux I__3045 (
            .O(N__14221),
            .I(N__14165));
    Span4Mux_v I__3044 (
            .O(N__14218),
            .I(N__14158));
    LocalMux I__3043 (
            .O(N__14215),
            .I(N__14158));
    LocalMux I__3042 (
            .O(N__14210),
            .I(N__14158));
    InMux I__3041 (
            .O(N__14207),
            .I(N__14155));
    InMux I__3040 (
            .O(N__14204),
            .I(N__14152));
    LocalMux I__3039 (
            .O(N__14201),
            .I(N__14149));
    Span4Mux_v I__3038 (
            .O(N__14196),
            .I(N__14140));
    LocalMux I__3037 (
            .O(N__14191),
            .I(N__14140));
    LocalMux I__3036 (
            .O(N__14188),
            .I(N__14140));
    LocalMux I__3035 (
            .O(N__14185),
            .I(N__14140));
    InMux I__3034 (
            .O(N__14184),
            .I(N__14137));
    Span4Mux_v I__3033 (
            .O(N__14181),
            .I(N__14126));
    Span4Mux_h I__3032 (
            .O(N__14176),
            .I(N__14126));
    LocalMux I__3031 (
            .O(N__14173),
            .I(N__14126));
    LocalMux I__3030 (
            .O(N__14168),
            .I(N__14126));
    LocalMux I__3029 (
            .O(N__14165),
            .I(N__14126));
    Span4Mux_v I__3028 (
            .O(N__14158),
            .I(N__14119));
    LocalMux I__3027 (
            .O(N__14155),
            .I(N__14119));
    LocalMux I__3026 (
            .O(N__14152),
            .I(N__14119));
    IoSpan4Mux I__3025 (
            .O(N__14149),
            .I(N__14116));
    Span4Mux_h I__3024 (
            .O(N__14140),
            .I(N__14111));
    LocalMux I__3023 (
            .O(N__14137),
            .I(N__14111));
    Span4Mux_v I__3022 (
            .O(N__14126),
            .I(N__14108));
    Span4Mux_h I__3021 (
            .O(N__14119),
            .I(N__14103));
    Span4Mux_s1_v I__3020 (
            .O(N__14116),
            .I(N__14103));
    Odrv4 I__3019 (
            .O(N__14111),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3018 (
            .O(N__14108),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3017 (
            .O(N__14103),
            .I(CONSTANT_ONE_NET));
    InMux I__3016 (
            .O(N__14096),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2));
    InMux I__3015 (
            .O(N__14093),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3));
    InMux I__3014 (
            .O(N__14090),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4));
    InMux I__3013 (
            .O(N__14087),
            .I(N__14084));
    LocalMux I__3012 (
            .O(N__14084),
            .I(N__14081));
    Odrv4 I__3011 (
            .O(N__14081),
            .I(un114_pixel_6_1_5__g2_0_1));
    InMux I__3010 (
            .O(N__14078),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1));
    CascadeMux I__3009 (
            .O(N__14075),
            .I(N__14071));
    CascadeMux I__3008 (
            .O(N__14074),
            .I(N__14068));
    InMux I__3007 (
            .O(N__14071),
            .I(N__14063));
    InMux I__3006 (
            .O(N__14068),
            .I(N__14063));
    LocalMux I__3005 (
            .O(N__14063),
            .I(charx_if_generate_plus_mult1_un33_sum_i_5));
    InMux I__3004 (
            .O(N__14060),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__3003 (
            .O(N__14057),
            .I(N__14054));
    LocalMux I__3002 (
            .O(N__14054),
            .I(charx_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__3001 (
            .O(N__14051),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__3000 (
            .O(N__14048),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1));
    CascadeMux I__2999 (
            .O(N__14045),
            .I(N__14042));
    InMux I__2998 (
            .O(N__14042),
            .I(N__14039));
    LocalMux I__2997 (
            .O(N__14039),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0));
    InMux I__2996 (
            .O(N__14036),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__2995 (
            .O(N__14033),
            .I(N__14030));
    LocalMux I__2994 (
            .O(N__14030),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1));
    InMux I__2993 (
            .O(N__14027),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__2992 (
            .O(N__14024),
            .I(N__14021));
    LocalMux I__2991 (
            .O(N__14021),
            .I(charx_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__2990 (
            .O(N__14018),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__2989 (
            .O(N__14015),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_));
    InMux I__2988 (
            .O(N__14012),
            .I(N__14007));
    InMux I__2987 (
            .O(N__14011),
            .I(N__14002));
    InMux I__2986 (
            .O(N__14010),
            .I(N__14002));
    LocalMux I__2985 (
            .O(N__14007),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    LocalMux I__2984 (
            .O(N__14002),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1));
    CascadeMux I__2983 (
            .O(N__13997),
            .I(N__13993));
    CascadeMux I__2982 (
            .O(N__13996),
            .I(N__13990));
    InMux I__2981 (
            .O(N__13993),
            .I(N__13985));
    InMux I__2980 (
            .O(N__13990),
            .I(N__13985));
    LocalMux I__2979 (
            .O(N__13985),
            .I(charx_if_generate_plus_mult1_un40_sum_i_5));
    InMux I__2978 (
            .O(N__13982),
            .I(N__13979));
    LocalMux I__2977 (
            .O(N__13979),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328));
    InMux I__2976 (
            .O(N__13976),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2));
    CascadeMux I__2975 (
            .O(N__13973),
            .I(N__13970));
    InMux I__2974 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__2973 (
            .O(N__13967),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538));
    InMux I__2972 (
            .O(N__13964),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_3));
    CascadeMux I__2971 (
            .O(N__13961),
            .I(N__13949));
    InMux I__2970 (
            .O(N__13960),
            .I(N__13940));
    InMux I__2969 (
            .O(N__13959),
            .I(N__13940));
    InMux I__2968 (
            .O(N__13958),
            .I(N__13937));
    InMux I__2967 (
            .O(N__13957),
            .I(N__13934));
    InMux I__2966 (
            .O(N__13956),
            .I(N__13931));
    InMux I__2965 (
            .O(N__13955),
            .I(N__13922));
    InMux I__2964 (
            .O(N__13954),
            .I(N__13922));
    InMux I__2963 (
            .O(N__13953),
            .I(N__13922));
    InMux I__2962 (
            .O(N__13952),
            .I(N__13922));
    InMux I__2961 (
            .O(N__13949),
            .I(N__13919));
    InMux I__2960 (
            .O(N__13948),
            .I(N__13909));
    InMux I__2959 (
            .O(N__13947),
            .I(N__13909));
    InMux I__2958 (
            .O(N__13946),
            .I(N__13909));
    InMux I__2957 (
            .O(N__13945),
            .I(N__13909));
    LocalMux I__2956 (
            .O(N__13940),
            .I(N__13906));
    LocalMux I__2955 (
            .O(N__13937),
            .I(N__13901));
    LocalMux I__2954 (
            .O(N__13934),
            .I(N__13901));
    LocalMux I__2953 (
            .O(N__13931),
            .I(N__13894));
    LocalMux I__2952 (
            .O(N__13922),
            .I(N__13894));
    LocalMux I__2951 (
            .O(N__13919),
            .I(N__13894));
    CascadeMux I__2950 (
            .O(N__13918),
            .I(N__13883));
    LocalMux I__2949 (
            .O(N__13909),
            .I(N__13880));
    Span4Mux_v I__2948 (
            .O(N__13906),
            .I(N__13875));
    Span4Mux_v I__2947 (
            .O(N__13901),
            .I(N__13875));
    Span4Mux_v I__2946 (
            .O(N__13894),
            .I(N__13872));
    InMux I__2945 (
            .O(N__13893),
            .I(N__13857));
    InMux I__2944 (
            .O(N__13892),
            .I(N__13857));
    InMux I__2943 (
            .O(N__13891),
            .I(N__13857));
    InMux I__2942 (
            .O(N__13890),
            .I(N__13857));
    InMux I__2941 (
            .O(N__13889),
            .I(N__13857));
    InMux I__2940 (
            .O(N__13888),
            .I(N__13857));
    InMux I__2939 (
            .O(N__13887),
            .I(N__13857));
    InMux I__2938 (
            .O(N__13886),
            .I(N__13852));
    InMux I__2937 (
            .O(N__13883),
            .I(N__13852));
    Odrv4 I__2936 (
            .O(N__13880),
            .I(CO3_0));
    Odrv4 I__2935 (
            .O(N__13875),
            .I(CO3_0));
    Odrv4 I__2934 (
            .O(N__13872),
            .I(CO3_0));
    LocalMux I__2933 (
            .O(N__13857),
            .I(CO3_0));
    LocalMux I__2932 (
            .O(N__13852),
            .I(CO3_0));
    InMux I__2931 (
            .O(N__13841),
            .I(N__13838));
    LocalMux I__2930 (
            .O(N__13838),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO));
    InMux I__2929 (
            .O(N__13835),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__2928 (
            .O(N__13832),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_));
    InMux I__2927 (
            .O(N__13829),
            .I(N__13820));
    InMux I__2926 (
            .O(N__13828),
            .I(N__13820));
    InMux I__2925 (
            .O(N__13827),
            .I(N__13820));
    LocalMux I__2924 (
            .O(N__13820),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    CascadeMux I__2923 (
            .O(N__13817),
            .I(N__13813));
    CascadeMux I__2922 (
            .O(N__13816),
            .I(N__13810));
    InMux I__2921 (
            .O(N__13813),
            .I(N__13805));
    InMux I__2920 (
            .O(N__13810),
            .I(N__13805));
    LocalMux I__2919 (
            .O(N__13805),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    InMux I__2918 (
            .O(N__13802),
            .I(N__13799));
    LocalMux I__2917 (
            .O(N__13799),
            .I(N__13796));
    Odrv12 I__2916 (
            .O(N__13796),
            .I(charx_if_generate_plus_mult1_un33_sum_i));
    InMux I__2915 (
            .O(N__13793),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1));
    InMux I__2914 (
            .O(N__13790),
            .I(N__13786));
    InMux I__2913 (
            .O(N__13789),
            .I(N__13783));
    LocalMux I__2912 (
            .O(N__13786),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    LocalMux I__2911 (
            .O(N__13783),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0));
    CascadeMux I__2910 (
            .O(N__13778),
            .I(N__13775));
    InMux I__2909 (
            .O(N__13775),
            .I(N__13772));
    LocalMux I__2908 (
            .O(N__13772),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0));
    InMux I__2907 (
            .O(N__13769),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__2906 (
            .O(N__13766),
            .I(N__13763));
    LocalMux I__2905 (
            .O(N__13763),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0));
    InMux I__2904 (
            .O(N__13760),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6));
    CascadeMux I__2903 (
            .O(N__13757),
            .I(N__13753));
    InMux I__2902 (
            .O(N__13756),
            .I(N__13745));
    InMux I__2901 (
            .O(N__13753),
            .I(N__13745));
    InMux I__2900 (
            .O(N__13752),
            .I(N__13745));
    LocalMux I__2899 (
            .O(N__13745),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0));
    InMux I__2898 (
            .O(N__13742),
            .I(N__13739));
    LocalMux I__2897 (
            .O(N__13739),
            .I(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx));
    InMux I__2896 (
            .O(N__13736),
            .I(N__13733));
    LocalMux I__2895 (
            .O(N__13733),
            .I(N__13730));
    Odrv4 I__2894 (
            .O(N__13730),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0));
    InMux I__2893 (
            .O(N__13727),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__2892 (
            .O(N__13724),
            .I(N__13721));
    InMux I__2891 (
            .O(N__13721),
            .I(N__13718));
    LocalMux I__2890 (
            .O(N__13718),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0));
    InMux I__2889 (
            .O(N__13715),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__2888 (
            .O(N__13712),
            .I(N__13709));
    LocalMux I__2887 (
            .O(N__13709),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__2886 (
            .O(N__13706),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__2885 (
            .O(N__13703),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7));
    InMux I__2884 (
            .O(N__13700),
            .I(N__13697));
    LocalMux I__2883 (
            .O(N__13697),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO));
    InMux I__2882 (
            .O(N__13694),
            .I(N__13690));
    CascadeMux I__2881 (
            .O(N__13693),
            .I(N__13687));
    LocalMux I__2880 (
            .O(N__13690),
            .I(N__13679));
    InMux I__2879 (
            .O(N__13687),
            .I(N__13675));
    CascadeMux I__2878 (
            .O(N__13686),
            .I(N__13672));
    CascadeMux I__2877 (
            .O(N__13685),
            .I(N__13668));
    InMux I__2876 (
            .O(N__13684),
            .I(N__13661));
    InMux I__2875 (
            .O(N__13683),
            .I(N__13661));
    InMux I__2874 (
            .O(N__13682),
            .I(N__13658));
    Span4Mux_v I__2873 (
            .O(N__13679),
            .I(N__13655));
    InMux I__2872 (
            .O(N__13678),
            .I(N__13652));
    LocalMux I__2871 (
            .O(N__13675),
            .I(N__13649));
    InMux I__2870 (
            .O(N__13672),
            .I(N__13644));
    InMux I__2869 (
            .O(N__13671),
            .I(N__13644));
    InMux I__2868 (
            .O(N__13668),
            .I(N__13639));
    InMux I__2867 (
            .O(N__13667),
            .I(N__13639));
    InMux I__2866 (
            .O(N__13666),
            .I(N__13636));
    LocalMux I__2865 (
            .O(N__13661),
            .I(N__13631));
    LocalMux I__2864 (
            .O(N__13658),
            .I(N__13631));
    Odrv4 I__2863 (
            .O(N__13655),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2862 (
            .O(N__13652),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2861 (
            .O(N__13649),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2860 (
            .O(N__13644),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2859 (
            .O(N__13639),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2858 (
            .O(N__13636),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv12 I__2857 (
            .O(N__13631),
            .I(charx_if_generate_plus_mult1_un33_sum));
    CascadeMux I__2856 (
            .O(N__13616),
            .I(N__13610));
    InMux I__2855 (
            .O(N__13615),
            .I(N__13606));
    InMux I__2854 (
            .O(N__13614),
            .I(N__13602));
    InMux I__2853 (
            .O(N__13613),
            .I(N__13599));
    InMux I__2852 (
            .O(N__13610),
            .I(N__13596));
    InMux I__2851 (
            .O(N__13609),
            .I(N__13593));
    LocalMux I__2850 (
            .O(N__13606),
            .I(N__13588));
    InMux I__2849 (
            .O(N__13605),
            .I(N__13585));
    LocalMux I__2848 (
            .O(N__13602),
            .I(N__13578));
    LocalMux I__2847 (
            .O(N__13599),
            .I(N__13578));
    LocalMux I__2846 (
            .O(N__13596),
            .I(N__13578));
    LocalMux I__2845 (
            .O(N__13593),
            .I(N__13575));
    InMux I__2844 (
            .O(N__13592),
            .I(N__13570));
    InMux I__2843 (
            .O(N__13591),
            .I(N__13570));
    Span4Mux_v I__2842 (
            .O(N__13588),
            .I(N__13565));
    LocalMux I__2841 (
            .O(N__13585),
            .I(N__13565));
    Span4Mux_v I__2840 (
            .O(N__13578),
            .I(N__13562));
    Odrv4 I__2839 (
            .O(N__13575),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__2838 (
            .O(N__13570),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2837 (
            .O(N__13565),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2836 (
            .O(N__13562),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum));
    CascadeMux I__2835 (
            .O(N__13553),
            .I(N__13547));
    InMux I__2834 (
            .O(N__13552),
            .I(N__13543));
    CascadeMux I__2833 (
            .O(N__13551),
            .I(N__13539));
    CascadeMux I__2832 (
            .O(N__13550),
            .I(N__13536));
    InMux I__2831 (
            .O(N__13547),
            .I(N__13530));
    InMux I__2830 (
            .O(N__13546),
            .I(N__13530));
    LocalMux I__2829 (
            .O(N__13543),
            .I(N__13527));
    InMux I__2828 (
            .O(N__13542),
            .I(N__13524));
    InMux I__2827 (
            .O(N__13539),
            .I(N__13517));
    InMux I__2826 (
            .O(N__13536),
            .I(N__13517));
    InMux I__2825 (
            .O(N__13535),
            .I(N__13517));
    LocalMux I__2824 (
            .O(N__13530),
            .I(N_520));
    Odrv4 I__2823 (
            .O(N__13527),
            .I(N_520));
    LocalMux I__2822 (
            .O(N__13524),
            .I(N_520));
    LocalMux I__2821 (
            .O(N__13517),
            .I(N_520));
    CascadeMux I__2820 (
            .O(N__13508),
            .I(N__13504));
    InMux I__2819 (
            .O(N__13507),
            .I(N__13501));
    InMux I__2818 (
            .O(N__13504),
            .I(N__13498));
    LocalMux I__2817 (
            .O(N__13501),
            .I(un5_visiblex_i_24));
    LocalMux I__2816 (
            .O(N__13498),
            .I(un5_visiblex_i_24));
    InMux I__2815 (
            .O(N__13493),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1));
    CascadeMux I__2814 (
            .O(N__13490),
            .I(N__13487));
    InMux I__2813 (
            .O(N__13487),
            .I(N__13484));
    LocalMux I__2812 (
            .O(N__13484),
            .I(N__13481));
    Odrv4 I__2811 (
            .O(N__13481),
            .I(column_1_if_generate_plus_mult1_un68_sum_iZ0));
    InMux I__2810 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__2809 (
            .O(N__13475),
            .I(if_generate_plus_mult1_un75_sum_cry_2_s));
    InMux I__2808 (
            .O(N__13472),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__2807 (
            .O(N__13469),
            .I(N__13466));
    LocalMux I__2806 (
            .O(N__13466),
            .I(N__13463));
    Odrv12 I__2805 (
            .O(N__13463),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    CascadeMux I__2804 (
            .O(N__13460),
            .I(N__13457));
    InMux I__2803 (
            .O(N__13457),
            .I(N__13454));
    LocalMux I__2802 (
            .O(N__13454),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__2801 (
            .O(N__13451),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__2800 (
            .O(N__13448),
            .I(N__13445));
    LocalMux I__2799 (
            .O(N__13445),
            .I(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__2798 (
            .O(N__13442),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__2797 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__2796 (
            .O(N__13436),
            .I(N__13433));
    Odrv12 I__2795 (
            .O(N__13433),
            .I(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__2794 (
            .O(N__13430),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__2793 (
            .O(N__13427),
            .I(N__13424));
    LocalMux I__2792 (
            .O(N__13424),
            .I(un116_pixel_2_ns_1_2));
    CascadeMux I__2791 (
            .O(N__13421),
            .I(N__13417));
    InMux I__2790 (
            .O(N__13420),
            .I(N__13412));
    InMux I__2789 (
            .O(N__13417),
            .I(N__13412));
    LocalMux I__2788 (
            .O(N__13412),
            .I(N__13409));
    Odrv12 I__2787 (
            .O(N__13409),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    InMux I__2786 (
            .O(N__13406),
            .I(N__13403));
    LocalMux I__2785 (
            .O(N__13403),
            .I(if_generate_plus_mult1_un75_sum_axb_4_l_fx));
    InMux I__2784 (
            .O(N__13400),
            .I(N__13397));
    LocalMux I__2783 (
            .O(N__13397),
            .I(N__13394));
    Odrv12 I__2782 (
            .O(N__13394),
            .I(beamY_RNII25UDD3_0Z0Z_0));
    CascadeMux I__2781 (
            .O(N__13391),
            .I(un116_pixel_7_ns_1_6_cascade_));
    InMux I__2780 (
            .O(N__13388),
            .I(N__13382));
    InMux I__2779 (
            .O(N__13387),
            .I(N__13382));
    LocalMux I__2778 (
            .O(N__13382),
            .I(N__13368));
    InMux I__2777 (
            .O(N__13381),
            .I(N__13365));
    InMux I__2776 (
            .O(N__13380),
            .I(N__13360));
    InMux I__2775 (
            .O(N__13379),
            .I(N__13360));
    InMux I__2774 (
            .O(N__13378),
            .I(N__13353));
    InMux I__2773 (
            .O(N__13377),
            .I(N__13353));
    InMux I__2772 (
            .O(N__13376),
            .I(N__13353));
    InMux I__2771 (
            .O(N__13375),
            .I(N__13350));
    InMux I__2770 (
            .O(N__13374),
            .I(N__13343));
    InMux I__2769 (
            .O(N__13373),
            .I(N__13343));
    InMux I__2768 (
            .O(N__13372),
            .I(N__13343));
    InMux I__2767 (
            .O(N__13371),
            .I(N__13340));
    Odrv4 I__2766 (
            .O(N__13368),
            .I(font_un3_pixel_29));
    LocalMux I__2765 (
            .O(N__13365),
            .I(font_un3_pixel_29));
    LocalMux I__2764 (
            .O(N__13360),
            .I(font_un3_pixel_29));
    LocalMux I__2763 (
            .O(N__13353),
            .I(font_un3_pixel_29));
    LocalMux I__2762 (
            .O(N__13350),
            .I(font_un3_pixel_29));
    LocalMux I__2761 (
            .O(N__13343),
            .I(font_un3_pixel_29));
    LocalMux I__2760 (
            .O(N__13340),
            .I(font_un3_pixel_29));
    CascadeMux I__2759 (
            .O(N__13325),
            .I(N__13322));
    InMux I__2758 (
            .O(N__13322),
            .I(N__13319));
    LocalMux I__2757 (
            .O(N__13319),
            .I(beamY_RNIBHJ7AMZ0Z_0));
    CascadeMux I__2756 (
            .O(N__13316),
            .I(N__13313));
    InMux I__2755 (
            .O(N__13313),
            .I(N__13310));
    LocalMux I__2754 (
            .O(N__13310),
            .I(N__13307));
    Odrv4 I__2753 (
            .O(N__13307),
            .I(column_1_if_generate_plus_mult1_un75_sum_iZ0));
    InMux I__2752 (
            .O(N__13304),
            .I(N__13301));
    LocalMux I__2751 (
            .O(N__13301),
            .I(G_340));
    InMux I__2750 (
            .O(N__13298),
            .I(N__13295));
    LocalMux I__2749 (
            .O(N__13295),
            .I(G_341));
    InMux I__2748 (
            .O(N__13292),
            .I(column_1_if_generate_plus_mult1_un82_sum_cry_4));
    CascadeMux I__2747 (
            .O(N__13289),
            .I(un5_rowlto0_cascade_));
    InMux I__2746 (
            .O(N__13286),
            .I(N__13283));
    LocalMux I__2745 (
            .O(N__13283),
            .I(beamY_RNIJ720T72Z0Z_0));
    InMux I__2744 (
            .O(N__13280),
            .I(N__13277));
    LocalMux I__2743 (
            .O(N__13277),
            .I(un116_pixel_5_ns_1_2));
    InMux I__2742 (
            .O(N__13274),
            .I(N__13271));
    LocalMux I__2741 (
            .O(N__13271),
            .I(beamY_RNIJDHE4C2Z0Z_1));
    CascadeMux I__2740 (
            .O(N__13268),
            .I(font_un126_pixel_6_am_cascade_));
    InMux I__2739 (
            .O(N__13265),
            .I(N__13262));
    LocalMux I__2738 (
            .O(N__13262),
            .I(font_un126_pixel_2_am));
    InMux I__2737 (
            .O(N__13259),
            .I(N__13256));
    LocalMux I__2736 (
            .O(N__13256),
            .I(beamX_RNIQ6MATS2Z0Z_0));
    InMux I__2735 (
            .O(N__13253),
            .I(N__13250));
    LocalMux I__2734 (
            .O(N__13250),
            .I(N__13244));
    InMux I__2733 (
            .O(N__13249),
            .I(N__13241));
    InMux I__2732 (
            .O(N__13248),
            .I(N__13238));
    InMux I__2731 (
            .O(N__13247),
            .I(N__13235));
    Odrv4 I__2730 (
            .O(N__13244),
            .I(un114_pixel_7_1_7__N_11_i_1));
    LocalMux I__2729 (
            .O(N__13241),
            .I(un114_pixel_7_1_7__N_11_i_1));
    LocalMux I__2728 (
            .O(N__13238),
            .I(un114_pixel_7_1_7__N_11_i_1));
    LocalMux I__2727 (
            .O(N__13235),
            .I(un114_pixel_7_1_7__N_11_i_1));
    CascadeMux I__2726 (
            .O(N__13226),
            .I(N_37_cascade_));
    CascadeMux I__2725 (
            .O(N__13223),
            .I(beamY_RNI05CI5A3_1Z0Z_0_cascade_));
    InMux I__2724 (
            .O(N__13220),
            .I(N__13217));
    LocalMux I__2723 (
            .O(N__13217),
            .I(beamY_RNI05CI5A3Z0Z_0));
    InMux I__2722 (
            .O(N__13214),
            .I(N__13211));
    LocalMux I__2721 (
            .O(N__13211),
            .I(beamY_RNII25UDD3_1Z0Z_0));
    CascadeMux I__2720 (
            .O(N__13208),
            .I(un116_pixel_7_ns_1_4_cascade_));
    InMux I__2719 (
            .O(N__13205),
            .I(N__13202));
    LocalMux I__2718 (
            .O(N__13202),
            .I(N__13199));
    Odrv4 I__2717 (
            .O(N__13199),
            .I(beamY_RNIFHEQCT1Z0Z_0));
    CascadeMux I__2716 (
            .O(N__13196),
            .I(beamY_RNIA4V0NM1Z0Z_0_cascade_));
    InMux I__2715 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__2714 (
            .O(N__13190),
            .I(Pixel_1_r_sn));
    CascadeMux I__2713 (
            .O(N__13187),
            .I(Pixel_1_r_rn_0_cascade_));
    InMux I__2712 (
            .O(N__13184),
            .I(N__13181));
    LocalMux I__2711 (
            .O(N__13181),
            .I(N_396));
    IoInMux I__2710 (
            .O(N__13178),
            .I(N__13174));
    IoInMux I__2709 (
            .O(N__13177),
            .I(N__13171));
    LocalMux I__2708 (
            .O(N__13174),
            .I(N__13168));
    LocalMux I__2707 (
            .O(N__13171),
            .I(N__13165));
    Span4Mux_s2_v I__2706 (
            .O(N__13168),
            .I(N__13162));
    Span4Mux_s3_v I__2705 (
            .O(N__13165),
            .I(N__13159));
    Span4Mux_v I__2704 (
            .O(N__13162),
            .I(N__13156));
    Span4Mux_h I__2703 (
            .O(N__13159),
            .I(N__13153));
    Odrv4 I__2702 (
            .O(N__13156),
            .I(Pixel_c));
    Odrv4 I__2701 (
            .O(N__13153),
            .I(Pixel_c));
    ClkMux I__2700 (
            .O(N__13148),
            .I(N__13103));
    ClkMux I__2699 (
            .O(N__13147),
            .I(N__13103));
    ClkMux I__2698 (
            .O(N__13146),
            .I(N__13103));
    ClkMux I__2697 (
            .O(N__13145),
            .I(N__13103));
    ClkMux I__2696 (
            .O(N__13144),
            .I(N__13103));
    ClkMux I__2695 (
            .O(N__13143),
            .I(N__13103));
    ClkMux I__2694 (
            .O(N__13142),
            .I(N__13103));
    ClkMux I__2693 (
            .O(N__13141),
            .I(N__13103));
    ClkMux I__2692 (
            .O(N__13140),
            .I(N__13103));
    ClkMux I__2691 (
            .O(N__13139),
            .I(N__13103));
    ClkMux I__2690 (
            .O(N__13138),
            .I(N__13103));
    ClkMux I__2689 (
            .O(N__13137),
            .I(N__13103));
    ClkMux I__2688 (
            .O(N__13136),
            .I(N__13103));
    ClkMux I__2687 (
            .O(N__13135),
            .I(N__13103));
    ClkMux I__2686 (
            .O(N__13134),
            .I(N__13103));
    GlobalMux I__2685 (
            .O(N__13103),
            .I(N__13100));
    gio2CtrlBuf I__2684 (
            .O(N__13100),
            .I(PixelClock_g));
    InMux I__2683 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__2682 (
            .O(N__13094),
            .I(m6Z0Z_1));
    InMux I__2681 (
            .O(N__13091),
            .I(N__13088));
    LocalMux I__2680 (
            .O(N__13088),
            .I(N__13085));
    Span4Mux_h I__2679 (
            .O(N__13085),
            .I(N__13082));
    Odrv4 I__2678 (
            .O(N__13082),
            .I(G_7_0_m2_1));
    CascadeMux I__2677 (
            .O(N__13079),
            .I(beamX_RNI1M3Q1V2Z0Z_0_cascade_));
    InMux I__2676 (
            .O(N__13076),
            .I(N__13073));
    LocalMux I__2675 (
            .O(N__13073),
            .I(N_1039_0_0));
    CascadeMux I__2674 (
            .O(N__13070),
            .I(font_un3_pixel_29_cascade_));
    CascadeMux I__2673 (
            .O(N__13067),
            .I(G_7_0_m4_2_1_1_cascade_));
    InMux I__2672 (
            .O(N__13064),
            .I(N__13061));
    LocalMux I__2671 (
            .O(N__13061),
            .I(G_7_0_m4_2_1));
    InMux I__2670 (
            .O(N__13058),
            .I(N__13055));
    LocalMux I__2669 (
            .O(N__13055),
            .I(N__13052));
    Odrv4 I__2668 (
            .O(N__13052),
            .I(beamY_RNINIKJ5A3Z0Z_1));
    CascadeMux I__2667 (
            .O(N__13049),
            .I(beamY_RNI7OTDJ61Z0Z_1_cascade_));
    InMux I__2666 (
            .O(N__13046),
            .I(N__13040));
    InMux I__2665 (
            .O(N__13045),
            .I(N__13040));
    LocalMux I__2664 (
            .O(N__13040),
            .I(N__13036));
    InMux I__2663 (
            .O(N__13039),
            .I(N__13033));
    Odrv4 I__2662 (
            .O(N__13036),
            .I(un4_row));
    LocalMux I__2661 (
            .O(N__13033),
            .I(un4_row));
    InMux I__2660 (
            .O(N__13028),
            .I(N__13025));
    LocalMux I__2659 (
            .O(N__13025),
            .I(N__13022));
    Span4Mux_h I__2658 (
            .O(N__13022),
            .I(N__13019));
    Odrv4 I__2657 (
            .O(N__13019),
            .I(beamY_RNIPG1SS93Z0Z_2));
    InMux I__2656 (
            .O(N__13016),
            .I(N__13013));
    LocalMux I__2655 (
            .O(N__13013),
            .I(N_23_0));
    InMux I__2654 (
            .O(N__13010),
            .I(N__13007));
    LocalMux I__2653 (
            .O(N__13007),
            .I(N_15_0));
    InMux I__2652 (
            .O(N__13004),
            .I(N__13001));
    LocalMux I__2651 (
            .O(N__13001),
            .I(N_342_0_0));
    CascadeMux I__2650 (
            .O(N__12998),
            .I(N_1045_0_cascade_));
    CascadeMux I__2649 (
            .O(N__12995),
            .I(N__12992));
    InMux I__2648 (
            .O(N__12992),
            .I(N__12989));
    LocalMux I__2647 (
            .O(N__12989),
            .I(column_1_if_generate_plus_mult1_un61_sum_iZ0));
    InMux I__2646 (
            .O(N__12986),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_1));
    CascadeMux I__2645 (
            .O(N__12983),
            .I(N__12980));
    InMux I__2644 (
            .O(N__12980),
            .I(N__12977));
    LocalMux I__2643 (
            .O(N__12977),
            .I(N__12974));
    Span4Mux_h I__2642 (
            .O(N__12974),
            .I(N__12971));
    Odrv4 I__2641 (
            .O(N__12971),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__2640 (
            .O(N__12968),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__2639 (
            .O(N__12965),
            .I(N__12959));
    InMux I__2638 (
            .O(N__12964),
            .I(N__12959));
    LocalMux I__2637 (
            .O(N__12959),
            .I(un5_rowlto3_i));
    CascadeMux I__2636 (
            .O(N__12956),
            .I(N__12953));
    InMux I__2635 (
            .O(N__12953),
            .I(N__12950));
    LocalMux I__2634 (
            .O(N__12950),
            .I(N__12947));
    Odrv4 I__2633 (
            .O(N__12947),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__2632 (
            .O(N__12944),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__2631 (
            .O(N__12941),
            .I(N__12938));
    LocalMux I__2630 (
            .O(N__12938),
            .I(N__12935));
    Odrv4 I__2629 (
            .O(N__12935),
            .I(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__2628 (
            .O(N__12932),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__2627 (
            .O(N__12929),
            .I(N__12926));
    LocalMux I__2626 (
            .O(N__12926),
            .I(Pixel_3_sqmuxa));
    InMux I__2625 (
            .O(N__12923),
            .I(N__12920));
    LocalMux I__2624 (
            .O(N__12920),
            .I(un114_pixel_6_1_5__font_un126_pixel_m_4));
    CascadeMux I__2623 (
            .O(N__12917),
            .I(N__12914));
    InMux I__2622 (
            .O(N__12914),
            .I(N__12911));
    LocalMux I__2621 (
            .O(N__12911),
            .I(N__12908));
    Span4Mux_h I__2620 (
            .O(N__12908),
            .I(N__12905));
    Odrv4 I__2619 (
            .O(N__12905),
            .I(un1_beamy_0_0));
    CascadeMux I__2618 (
            .O(N__12902),
            .I(un116_pixel_5_amZ0Z_6_cascade_));
    InMux I__2617 (
            .O(N__12899),
            .I(N__12896));
    LocalMux I__2616 (
            .O(N__12896),
            .I(un116_pixel_5_bmZ0Z_6));
    InMux I__2615 (
            .O(N__12893),
            .I(N__12889));
    CascadeMux I__2614 (
            .O(N__12892),
            .I(N__12886));
    LocalMux I__2613 (
            .O(N__12889),
            .I(N__12883));
    InMux I__2612 (
            .O(N__12886),
            .I(N__12880));
    Span4Mux_h I__2611 (
            .O(N__12883),
            .I(N__12877));
    LocalMux I__2610 (
            .O(N__12880),
            .I(un15_beamy));
    Odrv4 I__2609 (
            .O(N__12877),
            .I(un15_beamy));
    InMux I__2608 (
            .O(N__12872),
            .I(N__12869));
    LocalMux I__2607 (
            .O(N__12869),
            .I(N__12866));
    Span4Mux_v I__2606 (
            .O(N__12866),
            .I(N__12863));
    Odrv4 I__2605 (
            .O(N__12863),
            .I(un114_pixel_6_1_5__g0Z0Z_0));
    CascadeMux I__2604 (
            .O(N__12860),
            .I(un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_));
    InMux I__2603 (
            .O(N__12857),
            .I(N__12854));
    LocalMux I__2602 (
            .O(N__12854),
            .I(N__12851));
    Span4Mux_h I__2601 (
            .O(N__12851),
            .I(N__12848));
    Odrv4 I__2600 (
            .O(N__12848),
            .I(un114_pixel_6_1_5__font_un126_pixel_m_4_1_0));
    CascadeMux I__2599 (
            .O(N__12845),
            .I(un114_pixel_6_1_5__g0_2Z0Z_0_cascade_));
    InMux I__2598 (
            .O(N__12842),
            .I(N__12839));
    LocalMux I__2597 (
            .O(N__12839),
            .I(N__12836));
    Span4Mux_v I__2596 (
            .O(N__12836),
            .I(N__12833));
    Odrv4 I__2595 (
            .O(N__12833),
            .I(un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0));
    InMux I__2594 (
            .O(N__12830),
            .I(N__12827));
    LocalMux I__2593 (
            .O(N__12827),
            .I(N__12824));
    Span4Mux_h I__2592 (
            .O(N__12824),
            .I(N__12821));
    Odrv4 I__2591 (
            .O(N__12821),
            .I(un114_pixel_6_1_5__g0_1_0));
    CascadeMux I__2590 (
            .O(N__12818),
            .I(un114_pixel_6_1_5__g1Z0Z_0_cascade_));
    CascadeMux I__2589 (
            .O(N__12815),
            .I(N__12812));
    InMux I__2588 (
            .O(N__12812),
            .I(N__12809));
    LocalMux I__2587 (
            .O(N__12809),
            .I(charx_if_generate_plus_mult1_un26_sum_s_2_sf));
    InMux I__2586 (
            .O(N__12806),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1));
    CascadeMux I__2585 (
            .O(N__12803),
            .I(N__12800));
    InMux I__2584 (
            .O(N__12800),
            .I(N__12797));
    LocalMux I__2583 (
            .O(N__12797),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_2));
    InMux I__2582 (
            .O(N__12794),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__2581 (
            .O(N__12791),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__2580 (
            .O(N__12788),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4));
    CascadeMux I__2579 (
            .O(N__12785),
            .I(N__12782));
    InMux I__2578 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__2577 (
            .O(N__12779),
            .I(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx));
    CascadeMux I__2576 (
            .O(N__12776),
            .I(N__12773));
    InMux I__2575 (
            .O(N__12773),
            .I(N__12770));
    LocalMux I__2574 (
            .O(N__12770),
            .I(un5_visiblex_i_25));
    InMux I__2573 (
            .O(N__12767),
            .I(N__12762));
    InMux I__2572 (
            .O(N__12766),
            .I(N__12759));
    InMux I__2571 (
            .O(N__12765),
            .I(N__12756));
    LocalMux I__2570 (
            .O(N__12762),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    LocalMux I__2569 (
            .O(N__12759),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    LocalMux I__2568 (
            .O(N__12756),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    CascadeMux I__2567 (
            .O(N__12749),
            .I(N__12745));
    CascadeMux I__2566 (
            .O(N__12748),
            .I(N__12742));
    InMux I__2565 (
            .O(N__12745),
            .I(N__12739));
    InMux I__2564 (
            .O(N__12742),
            .I(N__12736));
    LocalMux I__2563 (
            .O(N__12739),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5));
    LocalMux I__2562 (
            .O(N__12736),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5));
    CascadeMux I__2561 (
            .O(N__12731),
            .I(N__12728));
    InMux I__2560 (
            .O(N__12728),
            .I(N__12725));
    LocalMux I__2559 (
            .O(N__12725),
            .I(un114_pixel_6_1_5__un4_rowZ0Z_0));
    CascadeMux I__2558 (
            .O(N__12722),
            .I(N__12719));
    InMux I__2557 (
            .O(N__12719),
            .I(N__12716));
    LocalMux I__2556 (
            .O(N__12716),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i));
    InMux I__2555 (
            .O(N__12713),
            .I(N__12710));
    LocalMux I__2554 (
            .O(N__12710),
            .I(N__12707));
    Odrv4 I__2553 (
            .O(N__12707),
            .I(column_1_if_generate_plus_mult1_un47_sum0_2));
    InMux I__2552 (
            .O(N__12704),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_1));
    InMux I__2551 (
            .O(N__12701),
            .I(N__12698));
    LocalMux I__2550 (
            .O(N__12698),
            .I(column_1_if_generate_plus_mult1_un47_sum0_3));
    InMux I__2549 (
            .O(N__12695),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_2));
    InMux I__2548 (
            .O(N__12692),
            .I(N__12689));
    LocalMux I__2547 (
            .O(N__12689),
            .I(column_1_if_generate_plus_mult1_un47_sum0_4));
    InMux I__2546 (
            .O(N__12686),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_3));
    InMux I__2545 (
            .O(N__12683),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_4));
    InMux I__2544 (
            .O(N__12680),
            .I(N__12677));
    LocalMux I__2543 (
            .O(N__12677),
            .I(if_generate_plus_mult1_un47_sum_0_cry_3_ma));
    InMux I__2542 (
            .O(N__12674),
            .I(N__12671));
    LocalMux I__2541 (
            .O(N__12671),
            .I(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx));
    CascadeMux I__2540 (
            .O(N__12668),
            .I(N__12665));
    InMux I__2539 (
            .O(N__12665),
            .I(N__12662));
    LocalMux I__2538 (
            .O(N__12662),
            .I(N_200_0_i));
    InMux I__2537 (
            .O(N__12659),
            .I(N__12656));
    LocalMux I__2536 (
            .O(N__12656),
            .I(un116_pixel_4_bmZ0Z_1));
    CascadeMux I__2535 (
            .O(N__12653),
            .I(un116_pixel_4_amZ0Z_1_cascade_));
    InMux I__2534 (
            .O(N__12650),
            .I(N__12647));
    LocalMux I__2533 (
            .O(N__12647),
            .I(un116_pixel_3_ns_1_1));
    InMux I__2532 (
            .O(N__12644),
            .I(N__12641));
    LocalMux I__2531 (
            .O(N__12641),
            .I(N__12638));
    Odrv12 I__2530 (
            .O(N__12638),
            .I(beamY_RNIHIRVUS1Z0Z_1));
    InMux I__2529 (
            .O(N__12635),
            .I(N__12632));
    LocalMux I__2528 (
            .O(N__12632),
            .I(un116_pixel_1_bmZ0Z_1));
    InMux I__2527 (
            .O(N__12629),
            .I(N__12626));
    LocalMux I__2526 (
            .O(N__12626),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421));
    InMux I__2525 (
            .O(N__12623),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__2524 (
            .O(N__12620),
            .I(N__12617));
    InMux I__2523 (
            .O(N__12617),
            .I(N__12614));
    LocalMux I__2522 (
            .O(N__12614),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1));
    InMux I__2521 (
            .O(N__12611),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__2520 (
            .O(N__12608),
            .I(N__12605));
    LocalMux I__2519 (
            .O(N__12605),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__2518 (
            .O(N__12602),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__2517 (
            .O(N__12599),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7));
    CascadeMux I__2516 (
            .O(N__12596),
            .I(N__12592));
    InMux I__2515 (
            .O(N__12595),
            .I(N__12588));
    InMux I__2514 (
            .O(N__12592),
            .I(N__12583));
    InMux I__2513 (
            .O(N__12591),
            .I(N__12583));
    LocalMux I__2512 (
            .O(N__12588),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1));
    LocalMux I__2511 (
            .O(N__12583),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1));
    InMux I__2510 (
            .O(N__12578),
            .I(N__12572));
    InMux I__2509 (
            .O(N__12577),
            .I(N__12572));
    LocalMux I__2508 (
            .O(N__12572),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8));
    CascadeMux I__2507 (
            .O(N__12569),
            .I(un114_pixel_3_i_a3_7_cascade_));
    InMux I__2506 (
            .O(N__12566),
            .I(N__12563));
    LocalMux I__2505 (
            .O(N__12563),
            .I(N__12559));
    InMux I__2504 (
            .O(N__12562),
            .I(N__12556));
    Odrv4 I__2503 (
            .O(N__12559),
            .I(column_0001_0));
    LocalMux I__2502 (
            .O(N__12556),
            .I(column_0001_0));
    CascadeMux I__2501 (
            .O(N__12551),
            .I(un116_pixel_3_ns_1_2_cascade_));
    InMux I__2500 (
            .O(N__12548),
            .I(N__12545));
    LocalMux I__2499 (
            .O(N__12545),
            .I(beamY_RNIDVSK5A3Z0Z_1));
    InMux I__2498 (
            .O(N__12542),
            .I(N__12539));
    LocalMux I__2497 (
            .O(N__12539),
            .I(N_13_0));
    InMux I__2496 (
            .O(N__12536),
            .I(N__12533));
    LocalMux I__2495 (
            .O(N__12533),
            .I(N__12530));
    Odrv4 I__2494 (
            .O(N__12530),
            .I(un114_pixel_0_1__N_6_mux_0));
    CascadeMux I__2493 (
            .O(N__12527),
            .I(un116_pixel_1_amZ0Z_1_cascade_));
    CascadeMux I__2492 (
            .O(N__12524),
            .I(un116_pixel_3_bmZ0Z_6_cascade_));
    CascadeMux I__2491 (
            .O(N__12521),
            .I(beamY_RNISJITRQ2Z0Z_1_cascade_));
    InMux I__2490 (
            .O(N__12518),
            .I(N__12515));
    LocalMux I__2489 (
            .O(N__12515),
            .I(N_12_0));
    CascadeMux I__2488 (
            .O(N__12512),
            .I(N_248_0_cascade_));
    InMux I__2487 (
            .O(N__12509),
            .I(N__12506));
    LocalMux I__2486 (
            .O(N__12506),
            .I(un116_pixel_3_ns_1_0_6));
    CascadeMux I__2485 (
            .O(N__12503),
            .I(N__12500));
    InMux I__2484 (
            .O(N__12500),
            .I(N__12497));
    LocalMux I__2483 (
            .O(N__12497),
            .I(N_25_mux));
    InMux I__2482 (
            .O(N__12494),
            .I(N__12491));
    LocalMux I__2481 (
            .O(N__12491),
            .I(N__12488));
    Span4Mux_h I__2480 (
            .O(N__12488),
            .I(N__12485));
    Odrv4 I__2479 (
            .O(N__12485),
            .I(font_un28_pixel_0_0_29));
    CascadeMux I__2478 (
            .O(N__12482),
            .I(un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_));
    InMux I__2477 (
            .O(N__12479),
            .I(N__12476));
    LocalMux I__2476 (
            .O(N__12476),
            .I(N_14_0));
    CascadeMux I__2475 (
            .O(N__12473),
            .I(column_0111_0_cascade_));
    CascadeMux I__2474 (
            .O(N__12470),
            .I(beamY_RNI05CI5A3_0Z0Z_0_cascade_));
    CascadeMux I__2473 (
            .O(N__12467),
            .I(beamY_RNIBABJS01Z0Z_1_cascade_));
    CascadeMux I__2472 (
            .O(N__12464),
            .I(N_21_0_cascade_));
    InMux I__2471 (
            .O(N__12461),
            .I(N__12458));
    LocalMux I__2470 (
            .O(N__12458),
            .I(N_22_0));
    InMux I__2469 (
            .O(N__12455),
            .I(N__12452));
    LocalMux I__2468 (
            .O(N__12452),
            .I(column_0111_0));
    InMux I__2467 (
            .O(N__12449),
            .I(N__12446));
    LocalMux I__2466 (
            .O(N__12446),
            .I(N__12443));
    Odrv4 I__2465 (
            .O(N__12443),
            .I(chessboardpixel_un174_pixel_0_1));
    InMux I__2464 (
            .O(N__12440),
            .I(N__12437));
    LocalMux I__2463 (
            .O(N__12437),
            .I(chessboardpixel_un200_pixel_0_1));
    InMux I__2462 (
            .O(N__12434),
            .I(N__12431));
    LocalMux I__2461 (
            .O(N__12431),
            .I(un114_pixel_6_1_5__un4_row_7Z0Z_1));
    InMux I__2460 (
            .O(N__12428),
            .I(N__12425));
    LocalMux I__2459 (
            .O(N__12425),
            .I(N_357_0));
    CascadeMux I__2458 (
            .O(N__12422),
            .I(N_18_0_cascade_));
    CascadeMux I__2457 (
            .O(N__12419),
            .I(N_7_0_cascade_));
    InMux I__2456 (
            .O(N__12416),
            .I(N__12413));
    LocalMux I__2455 (
            .O(N__12413),
            .I(N__12410));
    Odrv4 I__2454 (
            .O(N__12410),
            .I(if_generate_plus_mult1_un54_sum_axb_4_l_fx));
    CascadeMux I__2453 (
            .O(N__12407),
            .I(N__12404));
    InMux I__2452 (
            .O(N__12404),
            .I(N__12400));
    InMux I__2451 (
            .O(N__12403),
            .I(N__12397));
    LocalMux I__2450 (
            .O(N__12400),
            .I(N__12391));
    LocalMux I__2449 (
            .O(N__12397),
            .I(N__12391));
    InMux I__2448 (
            .O(N__12396),
            .I(N__12388));
    Odrv4 I__2447 (
            .O(N__12391),
            .I(N_571_i));
    LocalMux I__2446 (
            .O(N__12388),
            .I(N_571_i));
    InMux I__2445 (
            .O(N__12383),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2444 (
            .O(N__12380),
            .I(N__12377));
    LocalMux I__2443 (
            .O(N__12377),
            .I(N__12374));
    Odrv4 I__2442 (
            .O(N__12374),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__2441 (
            .O(N__12371),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__2440 (
            .O(N__12368),
            .I(if_generate_plus_mult1_un54_sum_s_5_cascade_));
    InMux I__2439 (
            .O(N__12365),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__2438 (
            .O(N__12362),
            .I(N__12357));
    InMux I__2437 (
            .O(N__12361),
            .I(N__12354));
    InMux I__2436 (
            .O(N__12360),
            .I(N__12351));
    LocalMux I__2435 (
            .O(N__12357),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__2434 (
            .O(N__12354),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__2433 (
            .O(N__12351),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    CascadeMux I__2432 (
            .O(N__12344),
            .I(N__12341));
    InMux I__2431 (
            .O(N__12341),
            .I(N__12338));
    LocalMux I__2430 (
            .O(N__12338),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    InMux I__2429 (
            .O(N__12335),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__2428 (
            .O(N__12332),
            .I(N__12326));
    InMux I__2427 (
            .O(N__12331),
            .I(N__12326));
    LocalMux I__2426 (
            .O(N__12326),
            .I(column_1_if_generate_plus_mult1_un54_sum_i_5));
    CascadeMux I__2425 (
            .O(N__12323),
            .I(N__12320));
    InMux I__2424 (
            .O(N__12320),
            .I(N__12317));
    LocalMux I__2423 (
            .O(N__12317),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__2422 (
            .O(N__12314),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__2421 (
            .O(N__12311),
            .I(N__12308));
    LocalMux I__2420 (
            .O(N__12308),
            .I(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__2419 (
            .O(N__12305),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2418 (
            .O(N__12302),
            .I(N__12299));
    InMux I__2417 (
            .O(N__12299),
            .I(N__12296));
    LocalMux I__2416 (
            .O(N__12296),
            .I(N_562_i));
    CascadeMux I__2415 (
            .O(N__12293),
            .I(N__12290));
    InMux I__2414 (
            .O(N__12290),
            .I(N__12287));
    LocalMux I__2413 (
            .O(N__12287),
            .I(N_11_0_i));
    CascadeMux I__2412 (
            .O(N__12284),
            .I(N__12281));
    InMux I__2411 (
            .O(N__12281),
            .I(N__12278));
    LocalMux I__2410 (
            .O(N__12278),
            .I(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx));
    InMux I__2409 (
            .O(N__12275),
            .I(N__12272));
    LocalMux I__2408 (
            .O(N__12272),
            .I(N__12267));
    InMux I__2407 (
            .O(N__12271),
            .I(N__12264));
    InMux I__2406 (
            .O(N__12270),
            .I(N__12261));
    Span4Mux_h I__2405 (
            .O(N__12267),
            .I(N__12251));
    LocalMux I__2404 (
            .O(N__12264),
            .I(N__12248));
    LocalMux I__2403 (
            .O(N__12261),
            .I(N__12245));
    InMux I__2402 (
            .O(N__12260),
            .I(N__12237));
    InMux I__2401 (
            .O(N__12259),
            .I(N__12237));
    InMux I__2400 (
            .O(N__12258),
            .I(N__12237));
    InMux I__2399 (
            .O(N__12257),
            .I(N__12230));
    InMux I__2398 (
            .O(N__12256),
            .I(N__12227));
    InMux I__2397 (
            .O(N__12255),
            .I(N__12224));
    InMux I__2396 (
            .O(N__12254),
            .I(N__12221));
    Span4Mux_h I__2395 (
            .O(N__12251),
            .I(N__12216));
    Span4Mux_h I__2394 (
            .O(N__12248),
            .I(N__12216));
    Span4Mux_v I__2393 (
            .O(N__12245),
            .I(N__12213));
    InMux I__2392 (
            .O(N__12244),
            .I(N__12210));
    LocalMux I__2391 (
            .O(N__12237),
            .I(N__12207));
    InMux I__2390 (
            .O(N__12236),
            .I(N__12198));
    InMux I__2389 (
            .O(N__12235),
            .I(N__12198));
    InMux I__2388 (
            .O(N__12234),
            .I(N__12198));
    InMux I__2387 (
            .O(N__12233),
            .I(N__12198));
    LocalMux I__2386 (
            .O(N__12230),
            .I(N__12191));
    LocalMux I__2385 (
            .O(N__12227),
            .I(N__12191));
    LocalMux I__2384 (
            .O(N__12224),
            .I(N__12191));
    LocalMux I__2383 (
            .O(N__12221),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2382 (
            .O(N__12216),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2381 (
            .O(N__12213),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    LocalMux I__2380 (
            .O(N__12210),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2379 (
            .O(N__12207),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    LocalMux I__2378 (
            .O(N__12198),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv12 I__2377 (
            .O(N__12191),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    InMux I__2376 (
            .O(N__12176),
            .I(N__12170));
    InMux I__2375 (
            .O(N__12175),
            .I(N__12165));
    InMux I__2374 (
            .O(N__12174),
            .I(N__12162));
    CascadeMux I__2373 (
            .O(N__12173),
            .I(N__12159));
    LocalMux I__2372 (
            .O(N__12170),
            .I(N__12155));
    InMux I__2371 (
            .O(N__12169),
            .I(N__12151));
    InMux I__2370 (
            .O(N__12168),
            .I(N__12148));
    LocalMux I__2369 (
            .O(N__12165),
            .I(N__12143));
    LocalMux I__2368 (
            .O(N__12162),
            .I(N__12143));
    InMux I__2367 (
            .O(N__12159),
            .I(N__12138));
    InMux I__2366 (
            .O(N__12158),
            .I(N__12138));
    Span4Mux_h I__2365 (
            .O(N__12155),
            .I(N__12135));
    InMux I__2364 (
            .O(N__12154),
            .I(N__12132));
    LocalMux I__2363 (
            .O(N__12151),
            .I(N__12129));
    LocalMux I__2362 (
            .O(N__12148),
            .I(N__12126));
    Odrv12 I__2361 (
            .O(N__12143),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    LocalMux I__2360 (
            .O(N__12138),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__2359 (
            .O(N__12135),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    LocalMux I__2358 (
            .O(N__12132),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__2357 (
            .O(N__12129),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    Odrv4 I__2356 (
            .O(N__12126),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3));
    InMux I__2355 (
            .O(N__12113),
            .I(N__12109));
    CascadeMux I__2354 (
            .O(N__12112),
            .I(N__12105));
    LocalMux I__2353 (
            .O(N__12109),
            .I(N__12098));
    InMux I__2352 (
            .O(N__12108),
            .I(N__12095));
    InMux I__2351 (
            .O(N__12105),
            .I(N__12092));
    InMux I__2350 (
            .O(N__12104),
            .I(N__12085));
    InMux I__2349 (
            .O(N__12103),
            .I(N__12085));
    InMux I__2348 (
            .O(N__12102),
            .I(N__12077));
    InMux I__2347 (
            .O(N__12101),
            .I(N__12077));
    Span4Mux_h I__2346 (
            .O(N__12098),
            .I(N__12074));
    LocalMux I__2345 (
            .O(N__12095),
            .I(N__12071));
    LocalMux I__2344 (
            .O(N__12092),
            .I(N__12068));
    InMux I__2343 (
            .O(N__12091),
            .I(N__12063));
    InMux I__2342 (
            .O(N__12090),
            .I(N__12063));
    LocalMux I__2341 (
            .O(N__12085),
            .I(N__12055));
    InMux I__2340 (
            .O(N__12084),
            .I(N__12050));
    InMux I__2339 (
            .O(N__12083),
            .I(N__12050));
    InMux I__2338 (
            .O(N__12082),
            .I(N__12047));
    LocalMux I__2337 (
            .O(N__12077),
            .I(N__12044));
    Span4Mux_h I__2336 (
            .O(N__12074),
            .I(N__12041));
    Span4Mux_v I__2335 (
            .O(N__12071),
            .I(N__12034));
    Span4Mux_v I__2334 (
            .O(N__12068),
            .I(N__12034));
    LocalMux I__2333 (
            .O(N__12063),
            .I(N__12034));
    InMux I__2332 (
            .O(N__12062),
            .I(N__12027));
    InMux I__2331 (
            .O(N__12061),
            .I(N__12027));
    InMux I__2330 (
            .O(N__12060),
            .I(N__12027));
    InMux I__2329 (
            .O(N__12059),
            .I(N__12022));
    InMux I__2328 (
            .O(N__12058),
            .I(N__12022));
    Span4Mux_h I__2327 (
            .O(N__12055),
            .I(N__12019));
    LocalMux I__2326 (
            .O(N__12050),
            .I(N__12012));
    LocalMux I__2325 (
            .O(N__12047),
            .I(N__12012));
    Span12Mux_s2_v I__2324 (
            .O(N__12044),
            .I(N__12012));
    Odrv4 I__2323 (
            .O(N__12041),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__2322 (
            .O(N__12034),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__2321 (
            .O(N__12027),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__2320 (
            .O(N__12022),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__2319 (
            .O(N__12019),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv12 I__2318 (
            .O(N__12012),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    CascadeMux I__2317 (
            .O(N__11999),
            .I(N__11996));
    InMux I__2316 (
            .O(N__11996),
            .I(N__11993));
    LocalMux I__2315 (
            .O(N__11993),
            .I(un114_pixel_6_1_5__un4_rowZ0Z_2));
    CascadeMux I__2314 (
            .O(N__11990),
            .I(N__11987));
    InMux I__2313 (
            .O(N__11987),
            .I(N__11984));
    LocalMux I__2312 (
            .O(N__11984),
            .I(if_generate_plus_mult1_un47_sum_m_1));
    InMux I__2311 (
            .O(N__11981),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__2310 (
            .O(N__11978),
            .I(N__11975));
    LocalMux I__2309 (
            .O(N__11975),
            .I(N__11971));
    InMux I__2308 (
            .O(N__11974),
            .I(N__11968));
    Odrv4 I__2307 (
            .O(N__11971),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    LocalMux I__2306 (
            .O(N__11968),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    CascadeMux I__2305 (
            .O(N__11963),
            .I(N__11960));
    InMux I__2304 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__2303 (
            .O(N__11957),
            .I(N__11954));
    Odrv12 I__2302 (
            .O(N__11954),
            .I(if_generate_plus_mult1_un47_sum_m_2));
    InMux I__2301 (
            .O(N__11951),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__2300 (
            .O(N__11948),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_4));
    CascadeMux I__2299 (
            .O(N__11945),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5_cascade_));
    CascadeMux I__2298 (
            .O(N__11942),
            .I(N__11939));
    InMux I__2297 (
            .O(N__11939),
            .I(N__11936));
    LocalMux I__2296 (
            .O(N__11936),
            .I(un5_visiblex_i_0_25));
    InMux I__2295 (
            .O(N__11933),
            .I(N__11930));
    LocalMux I__2294 (
            .O(N__11930),
            .I(charx_if_generate_plus_mult1_un26_sum_axb_3_i));
    CascadeMux I__2293 (
            .O(N__11927),
            .I(N__11924));
    InMux I__2292 (
            .O(N__11924),
            .I(N__11921));
    LocalMux I__2291 (
            .O(N__11921),
            .I(N__11918));
    Odrv4 I__2290 (
            .O(N__11918),
            .I(column_1_if_generate_plus_mult1_un47_sum1_4));
    InMux I__2289 (
            .O(N__11915),
            .I(N__11912));
    LocalMux I__2288 (
            .O(N__11912),
            .I(column_1_if_generate_plus_mult1_un47_sum1_3));
    CascadeMux I__2287 (
            .O(N__11909),
            .I(if_generate_plus_mult1_un47_sum_m_5_cascade_));
    CascadeMux I__2286 (
            .O(N__11906),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_));
    CascadeMux I__2285 (
            .O(N__11903),
            .I(N__11900));
    InMux I__2284 (
            .O(N__11900),
            .I(N__11897));
    LocalMux I__2283 (
            .O(N__11897),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2));
    InMux I__2282 (
            .O(N__11894),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__2281 (
            .O(N__11891),
            .I(N__11888));
    LocalMux I__2280 (
            .O(N__11888),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__2279 (
            .O(N__11885),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__2278 (
            .O(N__11882),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__2277 (
            .O(N__11879),
            .I(N__11874));
    InMux I__2276 (
            .O(N__11878),
            .I(N__11869));
    InMux I__2275 (
            .O(N__11877),
            .I(N__11869));
    LocalMux I__2274 (
            .O(N__11874),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2));
    LocalMux I__2273 (
            .O(N__11869),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2));
    CascadeMux I__2272 (
            .O(N__11864),
            .I(N__11861));
    InMux I__2271 (
            .O(N__11861),
            .I(N__11858));
    LocalMux I__2270 (
            .O(N__11858),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__2269 (
            .O(N__11855),
            .I(N__11849));
    InMux I__2268 (
            .O(N__11854),
            .I(N__11849));
    LocalMux I__2267 (
            .O(N__11849),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__2266 (
            .O(N__11846),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_1));
    InMux I__2265 (
            .O(N__11843),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_2));
    InMux I__2264 (
            .O(N__11840),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_3));
    InMux I__2263 (
            .O(N__11837),
            .I(N__11834));
    LocalMux I__2262 (
            .O(N__11834),
            .I(g1_0_1));
    CascadeMux I__2261 (
            .O(N__11831),
            .I(N__11824));
    CascadeMux I__2260 (
            .O(N__11830),
            .I(N__11819));
    CascadeMux I__2259 (
            .O(N__11829),
            .I(N__11816));
    CascadeMux I__2258 (
            .O(N__11828),
            .I(N__11812));
    InMux I__2257 (
            .O(N__11827),
            .I(N__11805));
    InMux I__2256 (
            .O(N__11824),
            .I(N__11800));
    InMux I__2255 (
            .O(N__11823),
            .I(N__11800));
    InMux I__2254 (
            .O(N__11822),
            .I(N__11797));
    InMux I__2253 (
            .O(N__11819),
            .I(N__11789));
    InMux I__2252 (
            .O(N__11816),
            .I(N__11789));
    InMux I__2251 (
            .O(N__11815),
            .I(N__11786));
    InMux I__2250 (
            .O(N__11812),
            .I(N__11783));
    CascadeMux I__2249 (
            .O(N__11811),
            .I(N__11777));
    InMux I__2248 (
            .O(N__11810),
            .I(N__11773));
    CascadeMux I__2247 (
            .O(N__11809),
            .I(N__11769));
    InMux I__2246 (
            .O(N__11808),
            .I(N__11766));
    LocalMux I__2245 (
            .O(N__11805),
            .I(N__11759));
    LocalMux I__2244 (
            .O(N__11800),
            .I(N__11759));
    LocalMux I__2243 (
            .O(N__11797),
            .I(N__11759));
    InMux I__2242 (
            .O(N__11796),
            .I(N__11756));
    InMux I__2241 (
            .O(N__11795),
            .I(N__11751));
    InMux I__2240 (
            .O(N__11794),
            .I(N__11751));
    LocalMux I__2239 (
            .O(N__11789),
            .I(N__11748));
    LocalMux I__2238 (
            .O(N__11786),
            .I(N__11743));
    LocalMux I__2237 (
            .O(N__11783),
            .I(N__11743));
    InMux I__2236 (
            .O(N__11782),
            .I(N__11740));
    InMux I__2235 (
            .O(N__11781),
            .I(N__11737));
    InMux I__2234 (
            .O(N__11780),
            .I(N__11734));
    InMux I__2233 (
            .O(N__11777),
            .I(N__11729));
    InMux I__2232 (
            .O(N__11776),
            .I(N__11729));
    LocalMux I__2231 (
            .O(N__11773),
            .I(N__11726));
    InMux I__2230 (
            .O(N__11772),
            .I(N__11721));
    InMux I__2229 (
            .O(N__11769),
            .I(N__11721));
    LocalMux I__2228 (
            .O(N__11766),
            .I(N__11718));
    Span4Mux_v I__2227 (
            .O(N__11759),
            .I(N__11715));
    LocalMux I__2226 (
            .O(N__11756),
            .I(N__11698));
    LocalMux I__2225 (
            .O(N__11751),
            .I(N__11698));
    Span4Mux_h I__2224 (
            .O(N__11748),
            .I(N__11698));
    Span4Mux_v I__2223 (
            .O(N__11743),
            .I(N__11698));
    LocalMux I__2222 (
            .O(N__11740),
            .I(N__11698));
    LocalMux I__2221 (
            .O(N__11737),
            .I(N__11698));
    LocalMux I__2220 (
            .O(N__11734),
            .I(N__11698));
    LocalMux I__2219 (
            .O(N__11729),
            .I(N__11698));
    Span4Mux_v I__2218 (
            .O(N__11726),
            .I(N__11693));
    LocalMux I__2217 (
            .O(N__11721),
            .I(N__11693));
    Span4Mux_h I__2216 (
            .O(N__11718),
            .I(N__11686));
    Span4Mux_v I__2215 (
            .O(N__11715),
            .I(N__11686));
    Span4Mux_v I__2214 (
            .O(N__11698),
            .I(N__11686));
    Span4Mux_h I__2213 (
            .O(N__11693),
            .I(N__11683));
    Odrv4 I__2212 (
            .O(N__11686),
            .I(beamYZ0Z_3));
    Odrv4 I__2211 (
            .O(N__11683),
            .I(beamYZ0Z_3));
    InMux I__2210 (
            .O(N__11678),
            .I(N__11674));
    InMux I__2209 (
            .O(N__11677),
            .I(N__11668));
    LocalMux I__2208 (
            .O(N__11674),
            .I(N__11665));
    InMux I__2207 (
            .O(N__11673),
            .I(N__11660));
    InMux I__2206 (
            .O(N__11672),
            .I(N__11660));
    CascadeMux I__2205 (
            .O(N__11671),
            .I(N__11654));
    LocalMux I__2204 (
            .O(N__11668),
            .I(N__11650));
    Span4Mux_h I__2203 (
            .O(N__11665),
            .I(N__11645));
    LocalMux I__2202 (
            .O(N__11660),
            .I(N__11645));
    InMux I__2201 (
            .O(N__11659),
            .I(N__11642));
    InMux I__2200 (
            .O(N__11658),
            .I(N__11633));
    InMux I__2199 (
            .O(N__11657),
            .I(N__11633));
    InMux I__2198 (
            .O(N__11654),
            .I(N__11633));
    InMux I__2197 (
            .O(N__11653),
            .I(N__11633));
    Span12Mux_s4_v I__2196 (
            .O(N__11650),
            .I(N__11630));
    Span4Mux_h I__2195 (
            .O(N__11645),
            .I(N__11627));
    LocalMux I__2194 (
            .O(N__11642),
            .I(N__11622));
    LocalMux I__2193 (
            .O(N__11633),
            .I(N__11622));
    Odrv12 I__2192 (
            .O(N__11630),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    Odrv4 I__2191 (
            .O(N__11627),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    Odrv12 I__2190 (
            .O(N__11622),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i));
    InMux I__2189 (
            .O(N__11615),
            .I(N__11612));
    LocalMux I__2188 (
            .O(N__11612),
            .I(g2));
    InMux I__2187 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__2186 (
            .O(N__11606),
            .I(m511_0_o2_1));
    InMux I__2185 (
            .O(N__11603),
            .I(N__11597));
    InMux I__2184 (
            .O(N__11602),
            .I(N__11597));
    LocalMux I__2183 (
            .O(N__11597),
            .I(N__11594));
    Span4Mux_v I__2182 (
            .O(N__11594),
            .I(N__11585));
    InMux I__2181 (
            .O(N__11593),
            .I(N__11582));
    InMux I__2180 (
            .O(N__11592),
            .I(N__11579));
    InMux I__2179 (
            .O(N__11591),
            .I(N__11570));
    InMux I__2178 (
            .O(N__11590),
            .I(N__11570));
    InMux I__2177 (
            .O(N__11589),
            .I(N__11570));
    InMux I__2176 (
            .O(N__11588),
            .I(N__11570));
    Odrv4 I__2175 (
            .O(N__11585),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2174 (
            .O(N__11582),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2173 (
            .O(N__11579),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    LocalMux I__2172 (
            .O(N__11570),
            .I(chary_if_generate_plus_mult1_un68_sum_axbxc5_0));
    InMux I__2171 (
            .O(N__11561),
            .I(N__11558));
    LocalMux I__2170 (
            .O(N__11558),
            .I(N_80_i));
    CEMux I__2169 (
            .O(N__11555),
            .I(N__11550));
    CEMux I__2168 (
            .O(N__11554),
            .I(N__11547));
    InMux I__2167 (
            .O(N__11553),
            .I(N__11539));
    LocalMux I__2166 (
            .O(N__11550),
            .I(N__11534));
    LocalMux I__2165 (
            .O(N__11547),
            .I(N__11534));
    CEMux I__2164 (
            .O(N__11546),
            .I(N__11531));
    CEMux I__2163 (
            .O(N__11545),
            .I(N__11527));
    CEMux I__2162 (
            .O(N__11544),
            .I(N__11524));
    CEMux I__2161 (
            .O(N__11543),
            .I(N__11521));
    InMux I__2160 (
            .O(N__11542),
            .I(N__11518));
    LocalMux I__2159 (
            .O(N__11539),
            .I(N__11515));
    Span4Mux_v I__2158 (
            .O(N__11534),
            .I(N__11510));
    LocalMux I__2157 (
            .O(N__11531),
            .I(N__11510));
    CEMux I__2156 (
            .O(N__11530),
            .I(N__11504));
    LocalMux I__2155 (
            .O(N__11527),
            .I(N__11501));
    LocalMux I__2154 (
            .O(N__11524),
            .I(N__11496));
    LocalMux I__2153 (
            .O(N__11521),
            .I(N__11496));
    LocalMux I__2152 (
            .O(N__11518),
            .I(N__11491));
    Span4Mux_v I__2151 (
            .O(N__11515),
            .I(N__11491));
    Span4Mux_v I__2150 (
            .O(N__11510),
            .I(N__11488));
    InMux I__2149 (
            .O(N__11509),
            .I(N__11485));
    InMux I__2148 (
            .O(N__11508),
            .I(N__11482));
    InMux I__2147 (
            .O(N__11507),
            .I(N__11479));
    LocalMux I__2146 (
            .O(N__11504),
            .I(N__11476));
    Span12Mux_s6_v I__2145 (
            .O(N__11501),
            .I(N__11473));
    Span4Mux_v I__2144 (
            .O(N__11496),
            .I(N__11466));
    Span4Mux_v I__2143 (
            .O(N__11491),
            .I(N__11466));
    Span4Mux_v I__2142 (
            .O(N__11488),
            .I(N__11466));
    LocalMux I__2141 (
            .O(N__11485),
            .I(un3_beamx_0));
    LocalMux I__2140 (
            .O(N__11482),
            .I(un3_beamx_0));
    LocalMux I__2139 (
            .O(N__11479),
            .I(un3_beamx_0));
    Odrv4 I__2138 (
            .O(N__11476),
            .I(un3_beamx_0));
    Odrv12 I__2137 (
            .O(N__11473),
            .I(un3_beamx_0));
    Odrv4 I__2136 (
            .O(N__11466),
            .I(un3_beamx_0));
    InMux I__2135 (
            .O(N__11453),
            .I(N__11450));
    LocalMux I__2134 (
            .O(N__11450),
            .I(N__11443));
    InMux I__2133 (
            .O(N__11449),
            .I(N__11440));
    InMux I__2132 (
            .O(N__11448),
            .I(N__11437));
    InMux I__2131 (
            .O(N__11447),
            .I(N__11434));
    InMux I__2130 (
            .O(N__11446),
            .I(N__11431));
    Span12Mux_s3_h I__2129 (
            .O(N__11443),
            .I(N__11422));
    LocalMux I__2128 (
            .O(N__11440),
            .I(N__11422));
    LocalMux I__2127 (
            .O(N__11437),
            .I(N__11419));
    LocalMux I__2126 (
            .O(N__11434),
            .I(N__11416));
    LocalMux I__2125 (
            .O(N__11431),
            .I(N__11413));
    InMux I__2124 (
            .O(N__11430),
            .I(N__11404));
    InMux I__2123 (
            .O(N__11429),
            .I(N__11404));
    InMux I__2122 (
            .O(N__11428),
            .I(N__11404));
    InMux I__2121 (
            .O(N__11427),
            .I(N__11404));
    Span12Mux_s8_h I__2120 (
            .O(N__11422),
            .I(N__11401));
    Span4Mux_h I__2119 (
            .O(N__11419),
            .I(N__11396));
    Span4Mux_s3_h I__2118 (
            .O(N__11416),
            .I(N__11396));
    Span4Mux_s3_h I__2117 (
            .O(N__11413),
            .I(N__11393));
    LocalMux I__2116 (
            .O(N__11404),
            .I(N__11390));
    Odrv12 I__2115 (
            .O(N__11401),
            .I(un5_beamx_0));
    Odrv4 I__2114 (
            .O(N__11396),
            .I(un5_beamx_0));
    Odrv4 I__2113 (
            .O(N__11393),
            .I(un5_beamx_0));
    Odrv4 I__2112 (
            .O(N__11390),
            .I(un5_beamx_0));
    CascadeMux I__2111 (
            .O(N__11381),
            .I(N__11371));
    InMux I__2110 (
            .O(N__11380),
            .I(N__11362));
    InMux I__2109 (
            .O(N__11379),
            .I(N__11359));
    InMux I__2108 (
            .O(N__11378),
            .I(N__11356));
    InMux I__2107 (
            .O(N__11377),
            .I(N__11353));
    InMux I__2106 (
            .O(N__11376),
            .I(N__11348));
    InMux I__2105 (
            .O(N__11375),
            .I(N__11348));
    InMux I__2104 (
            .O(N__11374),
            .I(N__11345));
    InMux I__2103 (
            .O(N__11371),
            .I(N__11342));
    InMux I__2102 (
            .O(N__11370),
            .I(N__11337));
    InMux I__2101 (
            .O(N__11369),
            .I(N__11337));
    InMux I__2100 (
            .O(N__11368),
            .I(N__11334));
    InMux I__2099 (
            .O(N__11367),
            .I(N__11325));
    InMux I__2098 (
            .O(N__11366),
            .I(N__11322));
    InMux I__2097 (
            .O(N__11365),
            .I(N__11318));
    LocalMux I__2096 (
            .O(N__11362),
            .I(N__11315));
    LocalMux I__2095 (
            .O(N__11359),
            .I(N__11312));
    LocalMux I__2094 (
            .O(N__11356),
            .I(N__11307));
    LocalMux I__2093 (
            .O(N__11353),
            .I(N__11307));
    LocalMux I__2092 (
            .O(N__11348),
            .I(N__11304));
    LocalMux I__2091 (
            .O(N__11345),
            .I(N__11295));
    LocalMux I__2090 (
            .O(N__11342),
            .I(N__11295));
    LocalMux I__2089 (
            .O(N__11337),
            .I(N__11295));
    LocalMux I__2088 (
            .O(N__11334),
            .I(N__11295));
    InMux I__2087 (
            .O(N__11333),
            .I(N__11288));
    InMux I__2086 (
            .O(N__11332),
            .I(N__11288));
    InMux I__2085 (
            .O(N__11331),
            .I(N__11288));
    InMux I__2084 (
            .O(N__11330),
            .I(N__11285));
    InMux I__2083 (
            .O(N__11329),
            .I(N__11280));
    InMux I__2082 (
            .O(N__11328),
            .I(N__11280));
    LocalMux I__2081 (
            .O(N__11325),
            .I(N__11277));
    LocalMux I__2080 (
            .O(N__11322),
            .I(N__11274));
    InMux I__2079 (
            .O(N__11321),
            .I(N__11271));
    LocalMux I__2078 (
            .O(N__11318),
            .I(N__11268));
    Span4Mux_v I__2077 (
            .O(N__11315),
            .I(N__11255));
    Span4Mux_v I__2076 (
            .O(N__11312),
            .I(N__11255));
    Span4Mux_v I__2075 (
            .O(N__11307),
            .I(N__11255));
    Span4Mux_v I__2074 (
            .O(N__11304),
            .I(N__11255));
    Span4Mux_v I__2073 (
            .O(N__11295),
            .I(N__11255));
    LocalMux I__2072 (
            .O(N__11288),
            .I(N__11255));
    LocalMux I__2071 (
            .O(N__11285),
            .I(N__11250));
    LocalMux I__2070 (
            .O(N__11280),
            .I(N__11250));
    Span4Mux_v I__2069 (
            .O(N__11277),
            .I(N__11245));
    Span4Mux_v I__2068 (
            .O(N__11274),
            .I(N__11245));
    LocalMux I__2067 (
            .O(N__11271),
            .I(N__11242));
    Span4Mux_h I__2066 (
            .O(N__11268),
            .I(N__11237));
    Span4Mux_h I__2065 (
            .O(N__11255),
            .I(N__11237));
    Span4Mux_h I__2064 (
            .O(N__11250),
            .I(N__11234));
    Odrv4 I__2063 (
            .O(N__11245),
            .I(beamYZ0Z_2));
    Odrv4 I__2062 (
            .O(N__11242),
            .I(beamYZ0Z_2));
    Odrv4 I__2061 (
            .O(N__11237),
            .I(beamYZ0Z_2));
    Odrv4 I__2060 (
            .O(N__11234),
            .I(beamYZ0Z_2));
    InMux I__2059 (
            .O(N__11225),
            .I(N__11222));
    LocalMux I__2058 (
            .O(N__11222),
            .I(N__11219));
    Odrv12 I__2057 (
            .O(N__11219),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0));
    InMux I__2056 (
            .O(N__11216),
            .I(N__11212));
    InMux I__2055 (
            .O(N__11215),
            .I(N__11209));
    LocalMux I__2054 (
            .O(N__11212),
            .I(beamY_RNIJH2N2PZ0Z_3));
    LocalMux I__2053 (
            .O(N__11209),
            .I(beamY_RNIJH2N2PZ0Z_3));
    CascadeMux I__2052 (
            .O(N__11204),
            .I(N__11201));
    InMux I__2051 (
            .O(N__11201),
            .I(N__11198));
    LocalMux I__2050 (
            .O(N__11198),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1));
    InMux I__2049 (
            .O(N__11195),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2048 (
            .O(N__11192),
            .I(N__11185));
    InMux I__2047 (
            .O(N__11191),
            .I(N__11185));
    InMux I__2046 (
            .O(N__11190),
            .I(N__11182));
    LocalMux I__2045 (
            .O(N__11185),
            .I(N__11179));
    LocalMux I__2044 (
            .O(N__11182),
            .I(un1_beamx_2));
    Odrv4 I__2043 (
            .O(N__11179),
            .I(un1_beamx_2));
    InMux I__2042 (
            .O(N__11174),
            .I(N__11163));
    InMux I__2041 (
            .O(N__11173),
            .I(N__11163));
    InMux I__2040 (
            .O(N__11172),
            .I(N__11163));
    InMux I__2039 (
            .O(N__11171),
            .I(N__11159));
    InMux I__2038 (
            .O(N__11170),
            .I(N__11156));
    LocalMux I__2037 (
            .O(N__11163),
            .I(N__11153));
    InMux I__2036 (
            .O(N__11162),
            .I(N__11150));
    LocalMux I__2035 (
            .O(N__11159),
            .I(beamXZ0Z_7));
    LocalMux I__2034 (
            .O(N__11156),
            .I(beamXZ0Z_7));
    Odrv4 I__2033 (
            .O(N__11153),
            .I(beamXZ0Z_7));
    LocalMux I__2032 (
            .O(N__11150),
            .I(beamXZ0Z_7));
    CascadeMux I__2031 (
            .O(N__11141),
            .I(N__11135));
    CascadeMux I__2030 (
            .O(N__11140),
            .I(N__11132));
    CascadeMux I__2029 (
            .O(N__11139),
            .I(N__11129));
    InMux I__2028 (
            .O(N__11138),
            .I(N__11126));
    InMux I__2027 (
            .O(N__11135),
            .I(N__11123));
    InMux I__2026 (
            .O(N__11132),
            .I(N__11120));
    InMux I__2025 (
            .O(N__11129),
            .I(N__11117));
    LocalMux I__2024 (
            .O(N__11126),
            .I(beamXZ0Z_10));
    LocalMux I__2023 (
            .O(N__11123),
            .I(beamXZ0Z_10));
    LocalMux I__2022 (
            .O(N__11120),
            .I(beamXZ0Z_10));
    LocalMux I__2021 (
            .O(N__11117),
            .I(beamXZ0Z_10));
    InMux I__2020 (
            .O(N__11108),
            .I(N__11105));
    LocalMux I__2019 (
            .O(N__11105),
            .I(un1_beamxlt10_0));
    IoInMux I__2018 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__2017 (
            .O(N__11099),
            .I(N__11095));
    IoInMux I__2016 (
            .O(N__11098),
            .I(N__11092));
    Span4Mux_s1_v I__2015 (
            .O(N__11095),
            .I(N__11089));
    LocalMux I__2014 (
            .O(N__11092),
            .I(N__11086));
    Sp12to4 I__2013 (
            .O(N__11089),
            .I(N__11083));
    Span4Mux_s3_v I__2012 (
            .O(N__11086),
            .I(N__11080));
    Span12Mux_s6_h I__2011 (
            .O(N__11083),
            .I(N__11077));
    Span4Mux_v I__2010 (
            .O(N__11080),
            .I(N__11074));
    Odrv12 I__2009 (
            .O(N__11077),
            .I(HSync_c));
    Odrv4 I__2008 (
            .O(N__11074),
            .I(HSync_c));
    InMux I__2007 (
            .O(N__11069),
            .I(N__11066));
    LocalMux I__2006 (
            .O(N__11066),
            .I(N__11063));
    Odrv4 I__2005 (
            .O(N__11063),
            .I(un114_pixel_6_1_5__un4_rowZ0Z_5));
    InMux I__2004 (
            .O(N__11060),
            .I(N__11056));
    InMux I__2003 (
            .O(N__11059),
            .I(N__11053));
    LocalMux I__2002 (
            .O(N__11056),
            .I(N__11044));
    LocalMux I__2001 (
            .O(N__11053),
            .I(N__11044));
    InMux I__2000 (
            .O(N__11052),
            .I(N__11035));
    InMux I__1999 (
            .O(N__11051),
            .I(N__11035));
    InMux I__1998 (
            .O(N__11050),
            .I(N__11035));
    InMux I__1997 (
            .O(N__11049),
            .I(N__11035));
    Span4Mux_v I__1996 (
            .O(N__11044),
            .I(N__11032));
    LocalMux I__1995 (
            .O(N__11035),
            .I(N__11029));
    Odrv4 I__1994 (
            .O(N__11032),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    Odrv4 I__1993 (
            .O(N__11029),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    CascadeMux I__1992 (
            .O(N__11024),
            .I(N__11021));
    InMux I__1991 (
            .O(N__11021),
            .I(N__11018));
    LocalMux I__1990 (
            .O(N__11018),
            .I(N__11014));
    InMux I__1989 (
            .O(N__11017),
            .I(N__11011));
    Span4Mux_v I__1988 (
            .O(N__11014),
            .I(N__11005));
    LocalMux I__1987 (
            .O(N__11011),
            .I(N__11002));
    InMux I__1986 (
            .O(N__11010),
            .I(N__10997));
    InMux I__1985 (
            .O(N__11009),
            .I(N__10997));
    InMux I__1984 (
            .O(N__11008),
            .I(N__10994));
    Odrv4 I__1983 (
            .O(N__11005),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1));
    Odrv4 I__1982 (
            .O(N__11002),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1));
    LocalMux I__1981 (
            .O(N__10997),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1));
    LocalMux I__1980 (
            .O(N__10994),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1));
    InMux I__1979 (
            .O(N__10985),
            .I(N__10982));
    LocalMux I__1978 (
            .O(N__10982),
            .I(N__10979));
    Span4Mux_h I__1977 (
            .O(N__10979),
            .I(N__10976));
    Odrv4 I__1976 (
            .O(N__10976),
            .I(if_generate_plus_mult1_un75_sum_axbxc5));
    InMux I__1975 (
            .O(N__10973),
            .I(N__10970));
    LocalMux I__1974 (
            .O(N__10970),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3));
    CascadeMux I__1973 (
            .O(N__10967),
            .I(un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_));
    InMux I__1972 (
            .O(N__10964),
            .I(N__10961));
    LocalMux I__1971 (
            .O(N__10961),
            .I(N__10958));
    Odrv4 I__1970 (
            .O(N__10958),
            .I(un114_pixel_6_1_5__un4_rowZ0Z_1));
    InMux I__1969 (
            .O(N__10955),
            .I(N__10952));
    LocalMux I__1968 (
            .O(N__10952),
            .I(N__10949));
    Span4Mux_h I__1967 (
            .O(N__10949),
            .I(N__10943));
    InMux I__1966 (
            .O(N__10948),
            .I(N__10938));
    InMux I__1965 (
            .O(N__10947),
            .I(N__10938));
    InMux I__1964 (
            .O(N__10946),
            .I(N__10935));
    Odrv4 I__1963 (
            .O(N__10943),
            .I(beamY_i_2));
    LocalMux I__1962 (
            .O(N__10938),
            .I(beamY_i_2));
    LocalMux I__1961 (
            .O(N__10935),
            .I(beamY_i_2));
    InMux I__1960 (
            .O(N__10928),
            .I(N__10925));
    LocalMux I__1959 (
            .O(N__10925),
            .I(N__10922));
    Span4Mux_v I__1958 (
            .O(N__10922),
            .I(N__10919));
    Odrv4 I__1957 (
            .O(N__10919),
            .I(un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1));
    InMux I__1956 (
            .O(N__10916),
            .I(N__10910));
    InMux I__1955 (
            .O(N__10915),
            .I(N__10910));
    LocalMux I__1954 (
            .O(N__10910),
            .I(N__10907));
    Span4Mux_h I__1953 (
            .O(N__10907),
            .I(N__10904));
    Span4Mux_h I__1952 (
            .O(N__10904),
            .I(N__10900));
    InMux I__1951 (
            .O(N__10903),
            .I(N__10897));
    Odrv4 I__1950 (
            .O(N__10900),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0));
    LocalMux I__1949 (
            .O(N__10897),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0));
    InMux I__1948 (
            .O(N__10892),
            .I(N__10889));
    LocalMux I__1947 (
            .O(N__10889),
            .I(N__10886));
    Span12Mux_s9_v I__1946 (
            .O(N__10886),
            .I(N__10883));
    Odrv12 I__1945 (
            .O(N__10883),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0));
    CascadeMux I__1944 (
            .O(N__10880),
            .I(chessboardpixel_un200_pixellt10_cascade_));
    InMux I__1943 (
            .O(N__10877),
            .I(N__10874));
    LocalMux I__1942 (
            .O(N__10874),
            .I(N__10871));
    Span4Mux_h I__1941 (
            .O(N__10871),
            .I(N__10868));
    Odrv4 I__1940 (
            .O(N__10868),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5));
    InMux I__1939 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__1938 (
            .O(N__10862),
            .I(N__10856));
    InMux I__1937 (
            .O(N__10861),
            .I(N__10846));
    InMux I__1936 (
            .O(N__10860),
            .I(N__10846));
    InMux I__1935 (
            .O(N__10859),
            .I(N__10846));
    Span4Mux_h I__1934 (
            .O(N__10856),
            .I(N__10843));
    InMux I__1933 (
            .O(N__10855),
            .I(N__10838));
    InMux I__1932 (
            .O(N__10854),
            .I(N__10838));
    InMux I__1931 (
            .O(N__10853),
            .I(N__10835));
    LocalMux I__1930 (
            .O(N__10846),
            .I(N__10832));
    Odrv4 I__1929 (
            .O(N__10843),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0));
    LocalMux I__1928 (
            .O(N__10838),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0));
    LocalMux I__1927 (
            .O(N__10835),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0));
    Odrv4 I__1926 (
            .O(N__10832),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0));
    CascadeMux I__1925 (
            .O(N__10823),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_));
    InMux I__1924 (
            .O(N__10820),
            .I(N__10817));
    LocalMux I__1923 (
            .O(N__10817),
            .I(un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1));
    InMux I__1922 (
            .O(N__10814),
            .I(N__10811));
    LocalMux I__1921 (
            .O(N__10811),
            .I(N__10807));
    InMux I__1920 (
            .O(N__10810),
            .I(N__10804));
    Odrv4 I__1919 (
            .O(N__10807),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0));
    LocalMux I__1918 (
            .O(N__10804),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0));
    CascadeMux I__1917 (
            .O(N__10799),
            .I(N__10796));
    InMux I__1916 (
            .O(N__10796),
            .I(N__10793));
    LocalMux I__1915 (
            .O(N__10793),
            .I(N__10790));
    Odrv4 I__1914 (
            .O(N__10790),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0));
    InMux I__1913 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__1912 (
            .O(N__10784),
            .I(un4_beamy_0));
    CascadeMux I__1911 (
            .O(N__10781),
            .I(un13_beamylt10_0_cascade_));
    CascadeMux I__1910 (
            .O(N__10778),
            .I(N__10775));
    InMux I__1909 (
            .O(N__10775),
            .I(N__10768));
    InMux I__1908 (
            .O(N__10774),
            .I(N__10765));
    CascadeMux I__1907 (
            .O(N__10773),
            .I(N__10762));
    InMux I__1906 (
            .O(N__10772),
            .I(N__10759));
    InMux I__1905 (
            .O(N__10771),
            .I(N__10756));
    LocalMux I__1904 (
            .O(N__10768),
            .I(N__10751));
    LocalMux I__1903 (
            .O(N__10765),
            .I(N__10751));
    InMux I__1902 (
            .O(N__10762),
            .I(N__10748));
    LocalMux I__1901 (
            .O(N__10759),
            .I(beamXZ0Z_4));
    LocalMux I__1900 (
            .O(N__10756),
            .I(beamXZ0Z_4));
    Odrv4 I__1899 (
            .O(N__10751),
            .I(beamXZ0Z_4));
    LocalMux I__1898 (
            .O(N__10748),
            .I(beamXZ0Z_4));
    InMux I__1897 (
            .O(N__10739),
            .I(N__10732));
    InMux I__1896 (
            .O(N__10738),
            .I(N__10729));
    CascadeMux I__1895 (
            .O(N__10737),
            .I(N__10726));
    InMux I__1894 (
            .O(N__10736),
            .I(N__10723));
    InMux I__1893 (
            .O(N__10735),
            .I(N__10720));
    LocalMux I__1892 (
            .O(N__10732),
            .I(N__10715));
    LocalMux I__1891 (
            .O(N__10729),
            .I(N__10715));
    InMux I__1890 (
            .O(N__10726),
            .I(N__10712));
    LocalMux I__1889 (
            .O(N__10723),
            .I(beamXZ0Z_3));
    LocalMux I__1888 (
            .O(N__10720),
            .I(beamXZ0Z_3));
    Odrv4 I__1887 (
            .O(N__10715),
            .I(beamXZ0Z_3));
    LocalMux I__1886 (
            .O(N__10712),
            .I(beamXZ0Z_3));
    CascadeMux I__1885 (
            .O(N__10703),
            .I(N__10700));
    InMux I__1884 (
            .O(N__10700),
            .I(N__10697));
    LocalMux I__1883 (
            .O(N__10697),
            .I(un18_beamylt5_0));
    InMux I__1882 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__1881 (
            .O(N__10691),
            .I(N__10683));
    CascadeMux I__1880 (
            .O(N__10690),
            .I(N__10680));
    InMux I__1879 (
            .O(N__10689),
            .I(N__10675));
    InMux I__1878 (
            .O(N__10688),
            .I(N__10675));
    CascadeMux I__1877 (
            .O(N__10687),
            .I(N__10672));
    InMux I__1876 (
            .O(N__10686),
            .I(N__10669));
    Span4Mux_h I__1875 (
            .O(N__10683),
            .I(N__10666));
    InMux I__1874 (
            .O(N__10680),
            .I(N__10663));
    LocalMux I__1873 (
            .O(N__10675),
            .I(N__10660));
    InMux I__1872 (
            .O(N__10672),
            .I(N__10657));
    LocalMux I__1871 (
            .O(N__10669),
            .I(beamXZ0Z_5));
    Odrv4 I__1870 (
            .O(N__10666),
            .I(beamXZ0Z_5));
    LocalMux I__1869 (
            .O(N__10663),
            .I(beamXZ0Z_5));
    Odrv4 I__1868 (
            .O(N__10660),
            .I(beamXZ0Z_5));
    LocalMux I__1867 (
            .O(N__10657),
            .I(beamXZ0Z_5));
    CascadeMux I__1866 (
            .O(N__10646),
            .I(un18_beamylt5_0_cascade_));
    InMux I__1865 (
            .O(N__10643),
            .I(N__10640));
    LocalMux I__1864 (
            .O(N__10640),
            .I(un114_pixel_6_1_5__un15_beamyZ0Z_0));
    InMux I__1863 (
            .O(N__10637),
            .I(N__10630));
    InMux I__1862 (
            .O(N__10636),
            .I(N__10627));
    CascadeMux I__1861 (
            .O(N__10635),
            .I(N__10624));
    InMux I__1860 (
            .O(N__10634),
            .I(N__10621));
    InMux I__1859 (
            .O(N__10633),
            .I(N__10618));
    LocalMux I__1858 (
            .O(N__10630),
            .I(N__10613));
    LocalMux I__1857 (
            .O(N__10627),
            .I(N__10613));
    InMux I__1856 (
            .O(N__10624),
            .I(N__10610));
    LocalMux I__1855 (
            .O(N__10621),
            .I(beamXZ0Z_8));
    LocalMux I__1854 (
            .O(N__10618),
            .I(beamXZ0Z_8));
    Odrv4 I__1853 (
            .O(N__10613),
            .I(beamXZ0Z_8));
    LocalMux I__1852 (
            .O(N__10610),
            .I(beamXZ0Z_8));
    CascadeMux I__1851 (
            .O(N__10601),
            .I(N__10595));
    InMux I__1850 (
            .O(N__10600),
            .I(N__10591));
    InMux I__1849 (
            .O(N__10599),
            .I(N__10588));
    InMux I__1848 (
            .O(N__10598),
            .I(N__10585));
    InMux I__1847 (
            .O(N__10595),
            .I(N__10582));
    InMux I__1846 (
            .O(N__10594),
            .I(N__10579));
    LocalMux I__1845 (
            .O(N__10591),
            .I(beamXZ0Z_9));
    LocalMux I__1844 (
            .O(N__10588),
            .I(beamXZ0Z_9));
    LocalMux I__1843 (
            .O(N__10585),
            .I(beamXZ0Z_9));
    LocalMux I__1842 (
            .O(N__10582),
            .I(beamXZ0Z_9));
    LocalMux I__1841 (
            .O(N__10579),
            .I(beamXZ0Z_9));
    InMux I__1840 (
            .O(N__10568),
            .I(N__10560));
    InMux I__1839 (
            .O(N__10567),
            .I(N__10555));
    InMux I__1838 (
            .O(N__10566),
            .I(N__10555));
    CascadeMux I__1837 (
            .O(N__10565),
            .I(N__10552));
    InMux I__1836 (
            .O(N__10564),
            .I(N__10549));
    InMux I__1835 (
            .O(N__10563),
            .I(N__10546));
    LocalMux I__1834 (
            .O(N__10560),
            .I(N__10541));
    LocalMux I__1833 (
            .O(N__10555),
            .I(N__10541));
    InMux I__1832 (
            .O(N__10552),
            .I(N__10538));
    LocalMux I__1831 (
            .O(N__10549),
            .I(beamXZ0Z_6));
    LocalMux I__1830 (
            .O(N__10546),
            .I(beamXZ0Z_6));
    Odrv4 I__1829 (
            .O(N__10541),
            .I(beamXZ0Z_6));
    LocalMux I__1828 (
            .O(N__10538),
            .I(beamXZ0Z_6));
    InMux I__1827 (
            .O(N__10529),
            .I(N__10526));
    LocalMux I__1826 (
            .O(N__10526),
            .I(un114_pixel_6_1_5__un18_beamylto9Z0Z_2));
    InMux I__1825 (
            .O(N__10523),
            .I(N__10520));
    LocalMux I__1824 (
            .O(N__10520),
            .I(N__10514));
    CascadeMux I__1823 (
            .O(N__10519),
            .I(N__10511));
    InMux I__1822 (
            .O(N__10518),
            .I(N__10508));
    InMux I__1821 (
            .O(N__10517),
            .I(N__10505));
    Span4Mux_v I__1820 (
            .O(N__10514),
            .I(N__10502));
    InMux I__1819 (
            .O(N__10511),
            .I(N__10499));
    LocalMux I__1818 (
            .O(N__10508),
            .I(beamXZ0Z_2));
    LocalMux I__1817 (
            .O(N__10505),
            .I(beamXZ0Z_2));
    Odrv4 I__1816 (
            .O(N__10502),
            .I(beamXZ0Z_2));
    LocalMux I__1815 (
            .O(N__10499),
            .I(beamXZ0Z_2));
    InMux I__1814 (
            .O(N__10490),
            .I(N__10483));
    CascadeMux I__1813 (
            .O(N__10489),
            .I(N__10480));
    InMux I__1812 (
            .O(N__10488),
            .I(N__10477));
    InMux I__1811 (
            .O(N__10487),
            .I(N__10474));
    InMux I__1810 (
            .O(N__10486),
            .I(N__10471));
    LocalMux I__1809 (
            .O(N__10483),
            .I(N__10468));
    InMux I__1808 (
            .O(N__10480),
            .I(N__10465));
    LocalMux I__1807 (
            .O(N__10477),
            .I(beamXZ0Z_1));
    LocalMux I__1806 (
            .O(N__10474),
            .I(beamXZ0Z_1));
    LocalMux I__1805 (
            .O(N__10471),
            .I(beamXZ0Z_1));
    Odrv4 I__1804 (
            .O(N__10468),
            .I(beamXZ0Z_1));
    LocalMux I__1803 (
            .O(N__10465),
            .I(beamXZ0Z_1));
    CascadeMux I__1802 (
            .O(N__10454),
            .I(N__10451));
    InMux I__1801 (
            .O(N__10451),
            .I(N__10448));
    LocalMux I__1800 (
            .O(N__10448),
            .I(un114_pixel_6_1_5__un13_beamylto2Z0Z_0));
    InMux I__1799 (
            .O(N__10445),
            .I(N__10439));
    InMux I__1798 (
            .O(N__10444),
            .I(N__10439));
    LocalMux I__1797 (
            .O(N__10439),
            .I(un114_pixel_6_1_5__un15_beamyZ0Z_1));
    InMux I__1796 (
            .O(N__10436),
            .I(N__10433));
    LocalMux I__1795 (
            .O(N__10433),
            .I(un4_beamy_0_0));
    CascadeMux I__1794 (
            .O(N__10430),
            .I(N__10427));
    InMux I__1793 (
            .O(N__10427),
            .I(N__10424));
    LocalMux I__1792 (
            .O(N__10424),
            .I(N__10421));
    Odrv4 I__1791 (
            .O(N__10421),
            .I(un114_pixel_6_1_5__g3_0_0_0));
    InMux I__1790 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__1789 (
            .O(N__10415),
            .I(un13_beamylt10_0));
    InMux I__1788 (
            .O(N__10412),
            .I(bfn_6_6_0_));
    InMux I__1787 (
            .O(N__10409),
            .I(un5_visiblex_cry_8));
    InMux I__1786 (
            .O(N__10406),
            .I(N__10403));
    LocalMux I__1785 (
            .O(N__10403),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0));
    InMux I__1784 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__1783 (
            .O(N__10397),
            .I(N__10393));
    InMux I__1782 (
            .O(N__10396),
            .I(N__10390));
    Span4Mux_h I__1781 (
            .O(N__10393),
            .I(N__10387));
    LocalMux I__1780 (
            .O(N__10390),
            .I(N__10384));
    Odrv4 I__1779 (
            .O(N__10387),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    Odrv4 I__1778 (
            .O(N__10384),
            .I(if_generate_plus_mult1_un54_sum_axbxc5));
    InMux I__1777 (
            .O(N__10379),
            .I(N__10376));
    LocalMux I__1776 (
            .O(N__10376),
            .I(N__10373));
    Span4Mux_v I__1775 (
            .O(N__10373),
            .I(N__10369));
    InMux I__1774 (
            .O(N__10372),
            .I(N__10366));
    Odrv4 I__1773 (
            .O(N__10369),
            .I(if_generate_plus_mult1_un61_sum_axbxc5));
    LocalMux I__1772 (
            .O(N__10366),
            .I(if_generate_plus_mult1_un61_sum_axbxc5));
    CascadeMux I__1771 (
            .O(N__10361),
            .I(un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_));
    InMux I__1770 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__1769 (
            .O(N__10355),
            .I(un114_pixel_6_1_5__un3_beamxZ0Z_7));
    CascadeMux I__1768 (
            .O(N__10352),
            .I(N__10349));
    InMux I__1767 (
            .O(N__10349),
            .I(N__10346));
    LocalMux I__1766 (
            .O(N__10346),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i));
    InMux I__1765 (
            .O(N__10343),
            .I(un5_visiblex_cry_0));
    InMux I__1764 (
            .O(N__10340),
            .I(un5_visiblex_cry_1));
    InMux I__1763 (
            .O(N__10337),
            .I(un5_visiblex_cry_2));
    InMux I__1762 (
            .O(N__10334),
            .I(un5_visiblex_cry_3));
    InMux I__1761 (
            .O(N__10331),
            .I(un5_visiblex_cry_4));
    InMux I__1760 (
            .O(N__10328),
            .I(un5_visiblex_cry_5));
    InMux I__1759 (
            .O(N__10325),
            .I(un5_visiblex_cry_6));
    InMux I__1758 (
            .O(N__10322),
            .I(N__10317));
    InMux I__1757 (
            .O(N__10321),
            .I(N__10314));
    CascadeMux I__1756 (
            .O(N__10320),
            .I(N__10311));
    LocalMux I__1755 (
            .O(N__10317),
            .I(N__10307));
    LocalMux I__1754 (
            .O(N__10314),
            .I(N__10302));
    InMux I__1753 (
            .O(N__10311),
            .I(N__10296));
    InMux I__1752 (
            .O(N__10310),
            .I(N__10296));
    Span4Mux_s3_h I__1751 (
            .O(N__10307),
            .I(N__10292));
    InMux I__1750 (
            .O(N__10306),
            .I(N__10287));
    InMux I__1749 (
            .O(N__10305),
            .I(N__10287));
    Span4Mux_s3_h I__1748 (
            .O(N__10302),
            .I(N__10284));
    InMux I__1747 (
            .O(N__10301),
            .I(N__10281));
    LocalMux I__1746 (
            .O(N__10296),
            .I(N__10278));
    InMux I__1745 (
            .O(N__10295),
            .I(N__10275));
    Odrv4 I__1744 (
            .O(N__10292),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1743 (
            .O(N__10287),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    Odrv4 I__1742 (
            .O(N__10284),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1741 (
            .O(N__10281),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    Odrv4 I__1740 (
            .O(N__10278),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1739 (
            .O(N__10275),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    CascadeMux I__1738 (
            .O(N__10262),
            .I(N__10254));
    CascadeMux I__1737 (
            .O(N__10261),
            .I(N__10250));
    InMux I__1736 (
            .O(N__10260),
            .I(N__10244));
    InMux I__1735 (
            .O(N__10259),
            .I(N__10244));
    CascadeMux I__1734 (
            .O(N__10258),
            .I(N__10234));
    InMux I__1733 (
            .O(N__10257),
            .I(N__10231));
    InMux I__1732 (
            .O(N__10254),
            .I(N__10228));
    InMux I__1731 (
            .O(N__10253),
            .I(N__10225));
    InMux I__1730 (
            .O(N__10250),
            .I(N__10222));
    CascadeMux I__1729 (
            .O(N__10249),
            .I(N__10219));
    LocalMux I__1728 (
            .O(N__10244),
            .I(N__10216));
    InMux I__1727 (
            .O(N__10243),
            .I(N__10213));
    InMux I__1726 (
            .O(N__10242),
            .I(N__10208));
    InMux I__1725 (
            .O(N__10241),
            .I(N__10205));
    InMux I__1724 (
            .O(N__10240),
            .I(N__10200));
    InMux I__1723 (
            .O(N__10239),
            .I(N__10200));
    CascadeMux I__1722 (
            .O(N__10238),
            .I(N__10195));
    InMux I__1721 (
            .O(N__10237),
            .I(N__10192));
    InMux I__1720 (
            .O(N__10234),
            .I(N__10189));
    LocalMux I__1719 (
            .O(N__10231),
            .I(N__10186));
    LocalMux I__1718 (
            .O(N__10228),
            .I(N__10183));
    LocalMux I__1717 (
            .O(N__10225),
            .I(N__10180));
    LocalMux I__1716 (
            .O(N__10222),
            .I(N__10177));
    InMux I__1715 (
            .O(N__10219),
            .I(N__10174));
    Span4Mux_v I__1714 (
            .O(N__10216),
            .I(N__10169));
    LocalMux I__1713 (
            .O(N__10213),
            .I(N__10169));
    InMux I__1712 (
            .O(N__10212),
            .I(N__10166));
    InMux I__1711 (
            .O(N__10211),
            .I(N__10163));
    LocalMux I__1710 (
            .O(N__10208),
            .I(N__10160));
    LocalMux I__1709 (
            .O(N__10205),
            .I(N__10155));
    LocalMux I__1708 (
            .O(N__10200),
            .I(N__10155));
    InMux I__1707 (
            .O(N__10199),
            .I(N__10152));
    InMux I__1706 (
            .O(N__10198),
            .I(N__10147));
    InMux I__1705 (
            .O(N__10195),
            .I(N__10147));
    LocalMux I__1704 (
            .O(N__10192),
            .I(N__10142));
    LocalMux I__1703 (
            .O(N__10189),
            .I(N__10142));
    Span4Mux_v I__1702 (
            .O(N__10186),
            .I(N__10137));
    Span4Mux_v I__1701 (
            .O(N__10183),
            .I(N__10137));
    Span4Mux_v I__1700 (
            .O(N__10180),
            .I(N__10128));
    Span4Mux_v I__1699 (
            .O(N__10177),
            .I(N__10128));
    LocalMux I__1698 (
            .O(N__10174),
            .I(N__10128));
    Span4Mux_s1_h I__1697 (
            .O(N__10169),
            .I(N__10128));
    LocalMux I__1696 (
            .O(N__10166),
            .I(N__10119));
    LocalMux I__1695 (
            .O(N__10163),
            .I(N__10119));
    Sp12to4 I__1694 (
            .O(N__10160),
            .I(N__10119));
    Span12Mux_s4_h I__1693 (
            .O(N__10155),
            .I(N__10119));
    LocalMux I__1692 (
            .O(N__10152),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    LocalMux I__1691 (
            .O(N__10147),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1690 (
            .O(N__10142),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1689 (
            .O(N__10137),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1688 (
            .O(N__10128),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv12 I__1687 (
            .O(N__10119),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1686 (
            .O(N__10106),
            .I(N__10101));
    CascadeMux I__1685 (
            .O(N__10105),
            .I(N__10098));
    InMux I__1684 (
            .O(N__10104),
            .I(N__10091));
    InMux I__1683 (
            .O(N__10101),
            .I(N__10087));
    InMux I__1682 (
            .O(N__10098),
            .I(N__10084));
    CascadeMux I__1681 (
            .O(N__10097),
            .I(N__10081));
    CascadeMux I__1680 (
            .O(N__10096),
            .I(N__10078));
    CascadeMux I__1679 (
            .O(N__10095),
            .I(N__10075));
    InMux I__1678 (
            .O(N__10094),
            .I(N__10072));
    LocalMux I__1677 (
            .O(N__10091),
            .I(N__10069));
    InMux I__1676 (
            .O(N__10090),
            .I(N__10066));
    LocalMux I__1675 (
            .O(N__10087),
            .I(N__10063));
    LocalMux I__1674 (
            .O(N__10084),
            .I(N__10060));
    InMux I__1673 (
            .O(N__10081),
            .I(N__10057));
    InMux I__1672 (
            .O(N__10078),
            .I(N__10054));
    InMux I__1671 (
            .O(N__10075),
            .I(N__10051));
    LocalMux I__1670 (
            .O(N__10072),
            .I(N__10044));
    Span4Mux_v I__1669 (
            .O(N__10069),
            .I(N__10044));
    LocalMux I__1668 (
            .O(N__10066),
            .I(N__10044));
    Span4Mux_v I__1667 (
            .O(N__10063),
            .I(N__10037));
    Span4Mux_h I__1666 (
            .O(N__10060),
            .I(N__10037));
    LocalMux I__1665 (
            .O(N__10057),
            .I(N__10037));
    LocalMux I__1664 (
            .O(N__10054),
            .I(N__10034));
    LocalMux I__1663 (
            .O(N__10051),
            .I(N__10029));
    Span4Mux_h I__1662 (
            .O(N__10044),
            .I(N__10029));
    Odrv4 I__1661 (
            .O(N__10037),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1660 (
            .O(N__10034),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1659 (
            .O(N__10029),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    InMux I__1658 (
            .O(N__10022),
            .I(N__10011));
    InMux I__1657 (
            .O(N__10021),
            .I(N__10011));
    InMux I__1656 (
            .O(N__10020),
            .I(N__10008));
    InMux I__1655 (
            .O(N__10019),
            .I(N__10005));
    InMux I__1654 (
            .O(N__10018),
            .I(N__10000));
    InMux I__1653 (
            .O(N__10017),
            .I(N__10000));
    InMux I__1652 (
            .O(N__10016),
            .I(N__9997));
    LocalMux I__1651 (
            .O(N__10011),
            .I(N__9994));
    LocalMux I__1650 (
            .O(N__10008),
            .I(N__9989));
    LocalMux I__1649 (
            .O(N__10005),
            .I(N__9989));
    LocalMux I__1648 (
            .O(N__10000),
            .I(N__9981));
    LocalMux I__1647 (
            .O(N__9997),
            .I(N__9976));
    Span4Mux_h I__1646 (
            .O(N__9994),
            .I(N__9976));
    Span4Mux_h I__1645 (
            .O(N__9989),
            .I(N__9973));
    InMux I__1644 (
            .O(N__9988),
            .I(N__9962));
    InMux I__1643 (
            .O(N__9987),
            .I(N__9962));
    InMux I__1642 (
            .O(N__9986),
            .I(N__9962));
    InMux I__1641 (
            .O(N__9985),
            .I(N__9962));
    InMux I__1640 (
            .O(N__9984),
            .I(N__9962));
    Odrv12 I__1639 (
            .O(N__9981),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    Odrv4 I__1638 (
            .O(N__9976),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    Odrv4 I__1637 (
            .O(N__9973),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    LocalMux I__1636 (
            .O(N__9962),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    InMux I__1635 (
            .O(N__9953),
            .I(N__9948));
    InMux I__1634 (
            .O(N__9952),
            .I(N__9943));
    InMux I__1633 (
            .O(N__9951),
            .I(N__9943));
    LocalMux I__1632 (
            .O(N__9948),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_5));
    LocalMux I__1631 (
            .O(N__9943),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_5));
    CascadeMux I__1630 (
            .O(N__9938),
            .I(chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_));
    InMux I__1629 (
            .O(N__9935),
            .I(N__9932));
    LocalMux I__1628 (
            .O(N__9932),
            .I(beamY_RNIL0E2QG2Z0Z_3));
    InMux I__1627 (
            .O(N__9929),
            .I(N__9926));
    LocalMux I__1626 (
            .O(N__9926),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93));
    InMux I__1625 (
            .O(N__9923),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__1624 (
            .O(N__9920),
            .I(N__9917));
    InMux I__1623 (
            .O(N__9917),
            .I(N__9914));
    LocalMux I__1622 (
            .O(N__9914),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4));
    InMux I__1621 (
            .O(N__9911),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1620 (
            .O(N__9908),
            .I(N__9905));
    LocalMux I__1619 (
            .O(N__9905),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__1618 (
            .O(N__9902),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1617 (
            .O(N__9899),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__1616 (
            .O(N__9896),
            .I(N__9892));
    InMux I__1615 (
            .O(N__9895),
            .I(N__9888));
    InMux I__1614 (
            .O(N__9892),
            .I(N__9883));
    InMux I__1613 (
            .O(N__9891),
            .I(N__9883));
    LocalMux I__1612 (
            .O(N__9888),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36));
    LocalMux I__1611 (
            .O(N__9883),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36));
    CascadeMux I__1610 (
            .O(N__9878),
            .I(N__9875));
    InMux I__1609 (
            .O(N__9875),
            .I(N__9872));
    LocalMux I__1608 (
            .O(N__9872),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__1607 (
            .O(N__9869),
            .I(N__9863));
    InMux I__1606 (
            .O(N__9868),
            .I(N__9863));
    LocalMux I__1605 (
            .O(N__9863),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8));
    InMux I__1604 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1603 (
            .O(N__9857),
            .I(g1));
    CascadeMux I__1602 (
            .O(N__9854),
            .I(N__9848));
    CascadeMux I__1601 (
            .O(N__9853),
            .I(N__9840));
    InMux I__1600 (
            .O(N__9852),
            .I(N__9836));
    InMux I__1599 (
            .O(N__9851),
            .I(N__9833));
    InMux I__1598 (
            .O(N__9848),
            .I(N__9830));
    InMux I__1597 (
            .O(N__9847),
            .I(N__9827));
    InMux I__1596 (
            .O(N__9846),
            .I(N__9822));
    InMux I__1595 (
            .O(N__9845),
            .I(N__9822));
    InMux I__1594 (
            .O(N__9844),
            .I(N__9817));
    InMux I__1593 (
            .O(N__9843),
            .I(N__9817));
    InMux I__1592 (
            .O(N__9840),
            .I(N__9814));
    InMux I__1591 (
            .O(N__9839),
            .I(N__9811));
    LocalMux I__1590 (
            .O(N__9836),
            .I(N__9808));
    LocalMux I__1589 (
            .O(N__9833),
            .I(N__9799));
    LocalMux I__1588 (
            .O(N__9830),
            .I(N__9799));
    LocalMux I__1587 (
            .O(N__9827),
            .I(N__9799));
    LocalMux I__1586 (
            .O(N__9822),
            .I(N__9799));
    LocalMux I__1585 (
            .O(N__9817),
            .I(N__9793));
    LocalMux I__1584 (
            .O(N__9814),
            .I(N__9793));
    LocalMux I__1583 (
            .O(N__9811),
            .I(N__9790));
    Span4Mux_v I__1582 (
            .O(N__9808),
            .I(N__9785));
    Span4Mux_v I__1581 (
            .O(N__9799),
            .I(N__9785));
    InMux I__1580 (
            .O(N__9798),
            .I(N__9782));
    Span4Mux_h I__1579 (
            .O(N__9793),
            .I(N__9779));
    Odrv4 I__1578 (
            .O(N__9790),
            .I(beamYZ0Z_4));
    Odrv4 I__1577 (
            .O(N__9785),
            .I(beamYZ0Z_4));
    LocalMux I__1576 (
            .O(N__9782),
            .I(beamYZ0Z_4));
    Odrv4 I__1575 (
            .O(N__9779),
            .I(beamYZ0Z_4));
    CascadeMux I__1574 (
            .O(N__9770),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_));
    InMux I__1573 (
            .O(N__9767),
            .I(N__9764));
    LocalMux I__1572 (
            .O(N__9764),
            .I(m511_0_x2_1_2));
    CascadeMux I__1571 (
            .O(N__9761),
            .I(G_7_0_m2_1_1_1_cascade_));
    CascadeMux I__1570 (
            .O(N__9758),
            .I(G_7_0_m2_1_1_cascade_));
    InMux I__1569 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__1568 (
            .O(N__9752),
            .I(G_7_0_m2_1_0));
    InMux I__1567 (
            .O(N__9749),
            .I(N__9739));
    InMux I__1566 (
            .O(N__9748),
            .I(N__9739));
    InMux I__1565 (
            .O(N__9747),
            .I(N__9739));
    InMux I__1564 (
            .O(N__9746),
            .I(N__9736));
    LocalMux I__1563 (
            .O(N__9739),
            .I(N__9733));
    LocalMux I__1562 (
            .O(N__9736),
            .I(N__9730));
    Span4Mux_h I__1561 (
            .O(N__9733),
            .I(N__9727));
    Odrv12 I__1560 (
            .O(N__9730),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    Odrv4 I__1559 (
            .O(N__9727),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    InMux I__1558 (
            .O(N__9722),
            .I(N__9718));
    CascadeMux I__1557 (
            .O(N__9721),
            .I(N__9714));
    LocalMux I__1556 (
            .O(N__9718),
            .I(N__9710));
    InMux I__1555 (
            .O(N__9717),
            .I(N__9707));
    InMux I__1554 (
            .O(N__9714),
            .I(N__9702));
    InMux I__1553 (
            .O(N__9713),
            .I(N__9702));
    Odrv4 I__1552 (
            .O(N__9710),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    LocalMux I__1551 (
            .O(N__9707),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    LocalMux I__1550 (
            .O(N__9702),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    CascadeMux I__1549 (
            .O(N__9695),
            .I(un114_pixel_6_1_5__g0_1Z0Z_4_cascade_));
    InMux I__1548 (
            .O(N__9692),
            .I(N__9685));
    InMux I__1547 (
            .O(N__9691),
            .I(N__9682));
    InMux I__1546 (
            .O(N__9690),
            .I(N__9677));
    InMux I__1545 (
            .O(N__9689),
            .I(N__9677));
    InMux I__1544 (
            .O(N__9688),
            .I(N__9674));
    LocalMux I__1543 (
            .O(N__9685),
            .I(N__9665));
    LocalMux I__1542 (
            .O(N__9682),
            .I(N__9665));
    LocalMux I__1541 (
            .O(N__9677),
            .I(N__9660));
    LocalMux I__1540 (
            .O(N__9674),
            .I(N__9660));
    InMux I__1539 (
            .O(N__9673),
            .I(N__9657));
    InMux I__1538 (
            .O(N__9672),
            .I(N__9654));
    InMux I__1537 (
            .O(N__9671),
            .I(N__9651));
    InMux I__1536 (
            .O(N__9670),
            .I(N__9648));
    Span4Mux_v I__1535 (
            .O(N__9665),
            .I(N__9645));
    Span4Mux_v I__1534 (
            .O(N__9660),
            .I(N__9640));
    LocalMux I__1533 (
            .O(N__9657),
            .I(N__9640));
    LocalMux I__1532 (
            .O(N__9654),
            .I(N__9637));
    LocalMux I__1531 (
            .O(N__9651),
            .I(beamYZ0Z_5));
    LocalMux I__1530 (
            .O(N__9648),
            .I(beamYZ0Z_5));
    Odrv4 I__1529 (
            .O(N__9645),
            .I(beamYZ0Z_5));
    Odrv4 I__1528 (
            .O(N__9640),
            .I(beamYZ0Z_5));
    Odrv4 I__1527 (
            .O(N__9637),
            .I(beamYZ0Z_5));
    InMux I__1526 (
            .O(N__9626),
            .I(N__9620));
    InMux I__1525 (
            .O(N__9625),
            .I(N__9617));
    InMux I__1524 (
            .O(N__9624),
            .I(N__9610));
    InMux I__1523 (
            .O(N__9623),
            .I(N__9610));
    LocalMux I__1522 (
            .O(N__9620),
            .I(N__9600));
    LocalMux I__1521 (
            .O(N__9617),
            .I(N__9600));
    InMux I__1520 (
            .O(N__9616),
            .I(N__9595));
    InMux I__1519 (
            .O(N__9615),
            .I(N__9595));
    LocalMux I__1518 (
            .O(N__9610),
            .I(N__9592));
    InMux I__1517 (
            .O(N__9609),
            .I(N__9589));
    InMux I__1516 (
            .O(N__9608),
            .I(N__9585));
    InMux I__1515 (
            .O(N__9607),
            .I(N__9580));
    InMux I__1514 (
            .O(N__9606),
            .I(N__9580));
    InMux I__1513 (
            .O(N__9605),
            .I(N__9577));
    Span4Mux_v I__1512 (
            .O(N__9600),
            .I(N__9574));
    LocalMux I__1511 (
            .O(N__9595),
            .I(N__9567));
    Span4Mux_v I__1510 (
            .O(N__9592),
            .I(N__9567));
    LocalMux I__1509 (
            .O(N__9589),
            .I(N__9567));
    InMux I__1508 (
            .O(N__9588),
            .I(N__9564));
    LocalMux I__1507 (
            .O(N__9585),
            .I(N__9561));
    LocalMux I__1506 (
            .O(N__9580),
            .I(N__9558));
    LocalMux I__1505 (
            .O(N__9577),
            .I(N__9553));
    Span4Mux_v I__1504 (
            .O(N__9574),
            .I(N__9553));
    Span4Mux_h I__1503 (
            .O(N__9567),
            .I(N__9550));
    LocalMux I__1502 (
            .O(N__9564),
            .I(N__9547));
    Span4Mux_v I__1501 (
            .O(N__9561),
            .I(N__9544));
    Span4Mux_s2_h I__1500 (
            .O(N__9558),
            .I(N__9541));
    Odrv4 I__1499 (
            .O(N__9553),
            .I(beamYZ0Z_9));
    Odrv4 I__1498 (
            .O(N__9550),
            .I(beamYZ0Z_9));
    Odrv12 I__1497 (
            .O(N__9547),
            .I(beamYZ0Z_9));
    Odrv4 I__1496 (
            .O(N__9544),
            .I(beamYZ0Z_9));
    Odrv4 I__1495 (
            .O(N__9541),
            .I(beamYZ0Z_9));
    CascadeMux I__1494 (
            .O(N__9530),
            .I(N__9527));
    InMux I__1493 (
            .O(N__9527),
            .I(N__9516));
    InMux I__1492 (
            .O(N__9526),
            .I(N__9516));
    InMux I__1491 (
            .O(N__9525),
            .I(N__9511));
    InMux I__1490 (
            .O(N__9524),
            .I(N__9511));
    InMux I__1489 (
            .O(N__9523),
            .I(N__9507));
    InMux I__1488 (
            .O(N__9522),
            .I(N__9502));
    InMux I__1487 (
            .O(N__9521),
            .I(N__9502));
    LocalMux I__1486 (
            .O(N__9516),
            .I(N__9496));
    LocalMux I__1485 (
            .O(N__9511),
            .I(N__9493));
    InMux I__1484 (
            .O(N__9510),
            .I(N__9488));
    LocalMux I__1483 (
            .O(N__9507),
            .I(N__9483));
    LocalMux I__1482 (
            .O(N__9502),
            .I(N__9483));
    InMux I__1481 (
            .O(N__9501),
            .I(N__9478));
    InMux I__1480 (
            .O(N__9500),
            .I(N__9473));
    InMux I__1479 (
            .O(N__9499),
            .I(N__9473));
    Span4Mux_v I__1478 (
            .O(N__9496),
            .I(N__9468));
    Span4Mux_v I__1477 (
            .O(N__9493),
            .I(N__9468));
    InMux I__1476 (
            .O(N__9492),
            .I(N__9463));
    InMux I__1475 (
            .O(N__9491),
            .I(N__9463));
    LocalMux I__1474 (
            .O(N__9488),
            .I(N__9460));
    Span4Mux_v I__1473 (
            .O(N__9483),
            .I(N__9457));
    InMux I__1472 (
            .O(N__9482),
            .I(N__9452));
    InMux I__1471 (
            .O(N__9481),
            .I(N__9452));
    LocalMux I__1470 (
            .O(N__9478),
            .I(N__9447));
    LocalMux I__1469 (
            .O(N__9473),
            .I(N__9447));
    Span4Mux_h I__1468 (
            .O(N__9468),
            .I(N__9442));
    LocalMux I__1467 (
            .O(N__9463),
            .I(N__9442));
    Odrv12 I__1466 (
            .O(N__9460),
            .I(beamYZ0Z_7));
    Odrv4 I__1465 (
            .O(N__9457),
            .I(beamYZ0Z_7));
    LocalMux I__1464 (
            .O(N__9452),
            .I(beamYZ0Z_7));
    Odrv12 I__1463 (
            .O(N__9447),
            .I(beamYZ0Z_7));
    Odrv4 I__1462 (
            .O(N__9442),
            .I(beamYZ0Z_7));
    CascadeMux I__1461 (
            .O(N__9431),
            .I(N__9427));
    InMux I__1460 (
            .O(N__9430),
            .I(N__9420));
    InMux I__1459 (
            .O(N__9427),
            .I(N__9420));
    InMux I__1458 (
            .O(N__9426),
            .I(N__9417));
    InMux I__1457 (
            .O(N__9425),
            .I(N__9414));
    LocalMux I__1456 (
            .O(N__9420),
            .I(N__9402));
    LocalMux I__1455 (
            .O(N__9417),
            .I(N__9402));
    LocalMux I__1454 (
            .O(N__9414),
            .I(N__9402));
    InMux I__1453 (
            .O(N__9413),
            .I(N__9399));
    InMux I__1452 (
            .O(N__9412),
            .I(N__9396));
    InMux I__1451 (
            .O(N__9411),
            .I(N__9393));
    InMux I__1450 (
            .O(N__9410),
            .I(N__9390));
    InMux I__1449 (
            .O(N__9409),
            .I(N__9387));
    Span4Mux_v I__1448 (
            .O(N__9402),
            .I(N__9382));
    LocalMux I__1447 (
            .O(N__9399),
            .I(N__9382));
    LocalMux I__1446 (
            .O(N__9396),
            .I(N__9377));
    LocalMux I__1445 (
            .O(N__9393),
            .I(N__9377));
    LocalMux I__1444 (
            .O(N__9390),
            .I(beamYZ0Z_6));
    LocalMux I__1443 (
            .O(N__9387),
            .I(beamYZ0Z_6));
    Odrv4 I__1442 (
            .O(N__9382),
            .I(beamYZ0Z_6));
    Odrv4 I__1441 (
            .O(N__9377),
            .I(beamYZ0Z_6));
    InMux I__1440 (
            .O(N__9368),
            .I(N__9365));
    LocalMux I__1439 (
            .O(N__9365),
            .I(N__9362));
    Odrv4 I__1438 (
            .O(N__9362),
            .I(un114_pixel_6_1_5__g0_0Z0Z_4));
    CascadeMux I__1437 (
            .O(N__9359),
            .I(un114_pixel_6_1_5__g0_0Z0Z_3_cascade_));
    CascadeMux I__1436 (
            .O(N__9356),
            .I(un114_pixel_6_1_5__g2_0Z0Z_0_cascade_));
    CascadeMux I__1435 (
            .O(N__9353),
            .I(N__9341));
    InMux I__1434 (
            .O(N__9352),
            .I(N__9337));
    InMux I__1433 (
            .O(N__9351),
            .I(N__9332));
    InMux I__1432 (
            .O(N__9350),
            .I(N__9329));
    InMux I__1431 (
            .O(N__9349),
            .I(N__9325));
    InMux I__1430 (
            .O(N__9348),
            .I(N__9320));
    InMux I__1429 (
            .O(N__9347),
            .I(N__9320));
    InMux I__1428 (
            .O(N__9346),
            .I(N__9315));
    InMux I__1427 (
            .O(N__9345),
            .I(N__9315));
    InMux I__1426 (
            .O(N__9344),
            .I(N__9310));
    InMux I__1425 (
            .O(N__9341),
            .I(N__9310));
    InMux I__1424 (
            .O(N__9340),
            .I(N__9307));
    LocalMux I__1423 (
            .O(N__9337),
            .I(N__9304));
    InMux I__1422 (
            .O(N__9336),
            .I(N__9299));
    InMux I__1421 (
            .O(N__9335),
            .I(N__9299));
    LocalMux I__1420 (
            .O(N__9332),
            .I(N__9290));
    LocalMux I__1419 (
            .O(N__9329),
            .I(N__9290));
    InMux I__1418 (
            .O(N__9328),
            .I(N__9287));
    LocalMux I__1417 (
            .O(N__9325),
            .I(N__9280));
    LocalMux I__1416 (
            .O(N__9320),
            .I(N__9280));
    LocalMux I__1415 (
            .O(N__9315),
            .I(N__9280));
    LocalMux I__1414 (
            .O(N__9310),
            .I(N__9277));
    LocalMux I__1413 (
            .O(N__9307),
            .I(N__9274));
    Span4Mux_v I__1412 (
            .O(N__9304),
            .I(N__9269));
    LocalMux I__1411 (
            .O(N__9299),
            .I(N__9269));
    InMux I__1410 (
            .O(N__9298),
            .I(N__9262));
    InMux I__1409 (
            .O(N__9297),
            .I(N__9262));
    InMux I__1408 (
            .O(N__9296),
            .I(N__9262));
    InMux I__1407 (
            .O(N__9295),
            .I(N__9257));
    Span4Mux_v I__1406 (
            .O(N__9290),
            .I(N__9248));
    LocalMux I__1405 (
            .O(N__9287),
            .I(N__9248));
    Span4Mux_v I__1404 (
            .O(N__9280),
            .I(N__9248));
    Span4Mux_v I__1403 (
            .O(N__9277),
            .I(N__9248));
    Span4Mux_v I__1402 (
            .O(N__9274),
            .I(N__9241));
    Span4Mux_h I__1401 (
            .O(N__9269),
            .I(N__9241));
    LocalMux I__1400 (
            .O(N__9262),
            .I(N__9241));
    InMux I__1399 (
            .O(N__9261),
            .I(N__9238));
    InMux I__1398 (
            .O(N__9260),
            .I(N__9235));
    LocalMux I__1397 (
            .O(N__9257),
            .I(beamYZ0Z_8));
    Odrv4 I__1396 (
            .O(N__9248),
            .I(beamYZ0Z_8));
    Odrv4 I__1395 (
            .O(N__9241),
            .I(beamYZ0Z_8));
    LocalMux I__1394 (
            .O(N__9238),
            .I(beamYZ0Z_8));
    LocalMux I__1393 (
            .O(N__9235),
            .I(beamYZ0Z_8));
    InMux I__1392 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__1391 (
            .O(N__9221),
            .I(N__9218));
    Odrv4 I__1390 (
            .O(N__9218),
            .I(un114_pixel_6_1_5__g0_0_1Z0Z_1));
    CascadeMux I__1389 (
            .O(N__9215),
            .I(un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_));
    CascadeMux I__1388 (
            .O(N__9212),
            .I(un114_pixel_6_1_5__un1_beamylto9_3_cascade_));
    IoInMux I__1387 (
            .O(N__9209),
            .I(N__9206));
    LocalMux I__1386 (
            .O(N__9206),
            .I(N__9203));
    IoSpan4Mux I__1385 (
            .O(N__9203),
            .I(N__9199));
    IoInMux I__1384 (
            .O(N__9202),
            .I(N__9196));
    Span4Mux_s0_v I__1383 (
            .O(N__9199),
            .I(N__9193));
    LocalMux I__1382 (
            .O(N__9196),
            .I(N__9190));
    Span4Mux_v I__1381 (
            .O(N__9193),
            .I(N__9187));
    Span4Mux_s3_v I__1380 (
            .O(N__9190),
            .I(N__9184));
    Span4Mux_v I__1379 (
            .O(N__9187),
            .I(N__9179));
    Span4Mux_v I__1378 (
            .O(N__9184),
            .I(N__9179));
    Odrv4 I__1377 (
            .O(N__9179),
            .I(VSync_c));
    InMux I__1376 (
            .O(N__9176),
            .I(N__9171));
    InMux I__1375 (
            .O(N__9175),
            .I(N__9166));
    InMux I__1374 (
            .O(N__9174),
            .I(N__9166));
    LocalMux I__1373 (
            .O(N__9171),
            .I(un8_beamy_3));
    LocalMux I__1372 (
            .O(N__9166),
            .I(un8_beamy_3));
    CascadeMux I__1371 (
            .O(N__9161),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_));
    InMux I__1370 (
            .O(N__9158),
            .I(N__9155));
    LocalMux I__1369 (
            .O(N__9155),
            .I(N__9152));
    Span4Mux_v I__1368 (
            .O(N__9152),
            .I(N__9145));
    InMux I__1367 (
            .O(N__9151),
            .I(N__9142));
    InMux I__1366 (
            .O(N__9150),
            .I(N__9139));
    InMux I__1365 (
            .O(N__9149),
            .I(N__9134));
    InMux I__1364 (
            .O(N__9148),
            .I(N__9134));
    Odrv4 I__1363 (
            .O(N__9145),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1362 (
            .O(N__9142),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1361 (
            .O(N__9139),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__1360 (
            .O(N__9134),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5));
    CascadeMux I__1359 (
            .O(N__9125),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_));
    CascadeMux I__1358 (
            .O(N__9122),
            .I(N__9117));
    CascadeMux I__1357 (
            .O(N__9121),
            .I(N__9113));
    InMux I__1356 (
            .O(N__9120),
            .I(N__9106));
    InMux I__1355 (
            .O(N__9117),
            .I(N__9101));
    InMux I__1354 (
            .O(N__9116),
            .I(N__9098));
    InMux I__1353 (
            .O(N__9113),
            .I(N__9092));
    InMux I__1352 (
            .O(N__9112),
            .I(N__9085));
    InMux I__1351 (
            .O(N__9111),
            .I(N__9085));
    InMux I__1350 (
            .O(N__9110),
            .I(N__9085));
    InMux I__1349 (
            .O(N__9109),
            .I(N__9082));
    LocalMux I__1348 (
            .O(N__9106),
            .I(N__9079));
    InMux I__1347 (
            .O(N__9105),
            .I(N__9076));
    InMux I__1346 (
            .O(N__9104),
            .I(N__9069));
    LocalMux I__1345 (
            .O(N__9101),
            .I(N__9066));
    LocalMux I__1344 (
            .O(N__9098),
            .I(N__9063));
    InMux I__1343 (
            .O(N__9097),
            .I(N__9055));
    InMux I__1342 (
            .O(N__9096),
            .I(N__9055));
    InMux I__1341 (
            .O(N__9095),
            .I(N__9055));
    LocalMux I__1340 (
            .O(N__9092),
            .I(N__9052));
    LocalMux I__1339 (
            .O(N__9085),
            .I(N__9049));
    LocalMux I__1338 (
            .O(N__9082),
            .I(N__9044));
    Span4Mux_s3_h I__1337 (
            .O(N__9079),
            .I(N__9044));
    LocalMux I__1336 (
            .O(N__9076),
            .I(N__9041));
    InMux I__1335 (
            .O(N__9075),
            .I(N__9032));
    InMux I__1334 (
            .O(N__9074),
            .I(N__9032));
    InMux I__1333 (
            .O(N__9073),
            .I(N__9032));
    InMux I__1332 (
            .O(N__9072),
            .I(N__9032));
    LocalMux I__1331 (
            .O(N__9069),
            .I(N__9029));
    Span4Mux_s2_h I__1330 (
            .O(N__9066),
            .I(N__9026));
    Span4Mux_s2_h I__1329 (
            .O(N__9063),
            .I(N__9023));
    InMux I__1328 (
            .O(N__9062),
            .I(N__9020));
    LocalMux I__1327 (
            .O(N__9055),
            .I(N__9017));
    Span4Mux_h I__1326 (
            .O(N__9052),
            .I(N__9012));
    Span4Mux_s3_h I__1325 (
            .O(N__9049),
            .I(N__9012));
    Span4Mux_v I__1324 (
            .O(N__9044),
            .I(N__9003));
    Span4Mux_s3_h I__1323 (
            .O(N__9041),
            .I(N__9003));
    LocalMux I__1322 (
            .O(N__9032),
            .I(N__9003));
    Span4Mux_s3_h I__1321 (
            .O(N__9029),
            .I(N__9003));
    Span4Mux_v I__1320 (
            .O(N__9026),
            .I(N__8998));
    Span4Mux_v I__1319 (
            .O(N__9023),
            .I(N__8998));
    LocalMux I__1318 (
            .O(N__9020),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1317 (
            .O(N__9017),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1316 (
            .O(N__9012),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1315 (
            .O(N__9003),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1314 (
            .O(N__8998),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    CascadeMux I__1313 (
            .O(N__8987),
            .I(N__8983));
    CascadeMux I__1312 (
            .O(N__8986),
            .I(N__8980));
    InMux I__1311 (
            .O(N__8983),
            .I(N__8975));
    InMux I__1310 (
            .O(N__8980),
            .I(N__8975));
    LocalMux I__1309 (
            .O(N__8975),
            .I(un4_beamylt8_0));
    InMux I__1308 (
            .O(N__8972),
            .I(un8_beamx_cry_6));
    InMux I__1307 (
            .O(N__8969),
            .I(un8_beamx_cry_7));
    InMux I__1306 (
            .O(N__8966),
            .I(bfn_5_7_0_));
    InMux I__1305 (
            .O(N__8963),
            .I(un8_beamx_cry_9));
    InMux I__1304 (
            .O(N__8960),
            .I(N__8957));
    LocalMux I__1303 (
            .O(N__8957),
            .I(row_1_if_generate_plus_mult1_un82_sum_axb4_i));
    InMux I__1302 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__1301 (
            .O(N__8951),
            .I(N__8948));
    Odrv4 I__1300 (
            .O(N__8948),
            .I(un114_pixel_6_1_5__un8_beamylto9Z0Z_0));
    InMux I__1299 (
            .O(N__8945),
            .I(N__8942));
    LocalMux I__1298 (
            .O(N__8942),
            .I(N__8939));
    Span4Mux_h I__1297 (
            .O(N__8939),
            .I(N__8936));
    Odrv4 I__1296 (
            .O(N__8936),
            .I(un8_beamylt9_0));
    InMux I__1295 (
            .O(N__8933),
            .I(N__8930));
    LocalMux I__1294 (
            .O(N__8930),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__1293 (
            .O(N__8927),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__1292 (
            .O(N__8924),
            .I(N__8920));
    InMux I__1291 (
            .O(N__8923),
            .I(N__8915));
    InMux I__1290 (
            .O(N__8920),
            .I(N__8908));
    InMux I__1289 (
            .O(N__8919),
            .I(N__8908));
    InMux I__1288 (
            .O(N__8918),
            .I(N__8908));
    LocalMux I__1287 (
            .O(N__8915),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0));
    LocalMux I__1286 (
            .O(N__8908),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0));
    InMux I__1285 (
            .O(N__8903),
            .I(N__8900));
    LocalMux I__1284 (
            .O(N__8900),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8));
    CascadeMux I__1283 (
            .O(N__8897),
            .I(N__8894));
    InMux I__1282 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__1281 (
            .O(N__8891),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i));
    InMux I__1280 (
            .O(N__8888),
            .I(un8_beamx_cry_1));
    InMux I__1279 (
            .O(N__8885),
            .I(un8_beamx_cry_2));
    InMux I__1278 (
            .O(N__8882),
            .I(un8_beamx_cry_3));
    InMux I__1277 (
            .O(N__8879),
            .I(un8_beamx_cry_4));
    InMux I__1276 (
            .O(N__8876),
            .I(un8_beamx_cry_5));
    InMux I__1275 (
            .O(N__8873),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__1274 (
            .O(N__8870),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1273 (
            .O(N__8867),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__1272 (
            .O(N__8864),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__1271 (
            .O(N__8861),
            .I(N__8855));
    InMux I__1270 (
            .O(N__8860),
            .I(N__8855));
    LocalMux I__1269 (
            .O(N__8855),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__1268 (
            .O(N__8852),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1267 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__1266 (
            .O(N__8846),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6));
    InMux I__1265 (
            .O(N__8843),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5));
    CascadeMux I__1264 (
            .O(N__8840),
            .I(N__8837));
    InMux I__1263 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__1262 (
            .O(N__8834),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9));
    InMux I__1261 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__1260 (
            .O(N__8828),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0));
    InMux I__1259 (
            .O(N__8825),
            .I(N__8822));
    LocalMux I__1258 (
            .O(N__8822),
            .I(N__8819));
    Odrv12 I__1257 (
            .O(N__8819),
            .I(g2_1));
    CascadeMux I__1256 (
            .O(N__8816),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_));
    CascadeMux I__1255 (
            .O(N__8813),
            .I(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_));
    InMux I__1254 (
            .O(N__8810),
            .I(N__8801));
    InMux I__1253 (
            .O(N__8809),
            .I(N__8801));
    InMux I__1252 (
            .O(N__8808),
            .I(N__8798));
    CascadeMux I__1251 (
            .O(N__8807),
            .I(N__8795));
    InMux I__1250 (
            .O(N__8806),
            .I(N__8792));
    LocalMux I__1249 (
            .O(N__8801),
            .I(N__8787));
    LocalMux I__1248 (
            .O(N__8798),
            .I(N__8787));
    InMux I__1247 (
            .O(N__8795),
            .I(N__8783));
    LocalMux I__1246 (
            .O(N__8792),
            .I(N__8780));
    Span4Mux_v I__1245 (
            .O(N__8787),
            .I(N__8777));
    InMux I__1244 (
            .O(N__8786),
            .I(N__8774));
    LocalMux I__1243 (
            .O(N__8783),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    Odrv4 I__1242 (
            .O(N__8780),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    Odrv4 I__1241 (
            .O(N__8777),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    LocalMux I__1240 (
            .O(N__8774),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    InMux I__1239 (
            .O(N__8765),
            .I(N__8759));
    InMux I__1238 (
            .O(N__8764),
            .I(N__8759));
    LocalMux I__1237 (
            .O(N__8759),
            .I(N__8756));
    Odrv4 I__1236 (
            .O(N__8756),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i));
    InMux I__1235 (
            .O(N__8753),
            .I(N__8749));
    InMux I__1234 (
            .O(N__8752),
            .I(N__8746));
    LocalMux I__1233 (
            .O(N__8749),
            .I(N__8741));
    LocalMux I__1232 (
            .O(N__8746),
            .I(N__8741));
    Span4Mux_h I__1231 (
            .O(N__8741),
            .I(N__8737));
    InMux I__1230 (
            .O(N__8740),
            .I(N__8734));
    Odrv4 I__1229 (
            .O(N__8737),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_0));
    LocalMux I__1228 (
            .O(N__8734),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_0));
    InMux I__1227 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__1226 (
            .O(N__8726),
            .I(N__8723));
    Span4Mux_s3_h I__1225 (
            .O(N__8723),
            .I(N__8720));
    Odrv4 I__1224 (
            .O(N__8720),
            .I(chary_if_generate_plus_mult1_un68_sum_c5_0_0));
    CascadeMux I__1223 (
            .O(N__8717),
            .I(un114_pixel_6_1_5__g0_17Z0Z_1_cascade_));
    InMux I__1222 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__1221 (
            .O(N__8711),
            .I(chary_if_generate_plus_mult1_un75_sum_0_5));
    InMux I__1220 (
            .O(N__8708),
            .I(N__8705));
    LocalMux I__1219 (
            .O(N__8705),
            .I(N__8702));
    Odrv4 I__1218 (
            .O(N__8702),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_i));
    CascadeMux I__1217 (
            .O(N__8699),
            .I(N__8696));
    InMux I__1216 (
            .O(N__8696),
            .I(N__8692));
    InMux I__1215 (
            .O(N__8695),
            .I(N__8689));
    LocalMux I__1214 (
            .O(N__8692),
            .I(N__8686));
    LocalMux I__1213 (
            .O(N__8689),
            .I(chary_if_generate_plus_mult1_un61_sum_c4));
    Odrv12 I__1212 (
            .O(N__8686),
            .I(chary_if_generate_plus_mult1_un61_sum_c4));
    InMux I__1211 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__1210 (
            .O(N__8678),
            .I(g1_0_3));
    CascadeMux I__1209 (
            .O(N__8675),
            .I(N__8670));
    CascadeMux I__1208 (
            .O(N__8674),
            .I(N__8667));
    CascadeMux I__1207 (
            .O(N__8673),
            .I(N__8664));
    InMux I__1206 (
            .O(N__8670),
            .I(N__8659));
    InMux I__1205 (
            .O(N__8667),
            .I(N__8659));
    InMux I__1204 (
            .O(N__8664),
            .I(N__8656));
    LocalMux I__1203 (
            .O(N__8659),
            .I(N__8653));
    LocalMux I__1202 (
            .O(N__8656),
            .I(N__8648));
    Span4Mux_h I__1201 (
            .O(N__8653),
            .I(N__8645));
    InMux I__1200 (
            .O(N__8652),
            .I(N__8640));
    InMux I__1199 (
            .O(N__8651),
            .I(N__8640));
    Span4Mux_h I__1198 (
            .O(N__8648),
            .I(N__8637));
    Odrv4 I__1197 (
            .O(N__8645),
            .I(un5_visibley_c5));
    LocalMux I__1196 (
            .O(N__8640),
            .I(un5_visibley_c5));
    Odrv4 I__1195 (
            .O(N__8637),
            .I(un5_visibley_c5));
    InMux I__1194 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__1193 (
            .O(N__8627),
            .I(beamY_RNIP8FF1_2Z0Z_7));
    CascadeMux I__1192 (
            .O(N__8624),
            .I(un4_beamylt6_cascade_));
    InMux I__1191 (
            .O(N__8621),
            .I(N__8615));
    InMux I__1190 (
            .O(N__8620),
            .I(N__8615));
    LocalMux I__1189 (
            .O(N__8615),
            .I(N__8610));
    InMux I__1188 (
            .O(N__8614),
            .I(N__8606));
    InMux I__1187 (
            .O(N__8613),
            .I(N__8603));
    Span4Mux_v I__1186 (
            .O(N__8610),
            .I(N__8600));
    InMux I__1185 (
            .O(N__8609),
            .I(N__8597));
    LocalMux I__1184 (
            .O(N__8606),
            .I(N__8592));
    LocalMux I__1183 (
            .O(N__8603),
            .I(N__8592));
    Span4Mux_h I__1182 (
            .O(N__8600),
            .I(N__8589));
    LocalMux I__1181 (
            .O(N__8597),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    Odrv4 I__1180 (
            .O(N__8592),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    Odrv4 I__1179 (
            .O(N__8589),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    InMux I__1178 (
            .O(N__8582),
            .I(N__8572));
    InMux I__1177 (
            .O(N__8581),
            .I(N__8572));
    InMux I__1176 (
            .O(N__8580),
            .I(N__8566));
    InMux I__1175 (
            .O(N__8579),
            .I(N__8566));
    InMux I__1174 (
            .O(N__8578),
            .I(N__8561));
    InMux I__1173 (
            .O(N__8577),
            .I(N__8561));
    LocalMux I__1172 (
            .O(N__8572),
            .I(N__8558));
    CascadeMux I__1171 (
            .O(N__8571),
            .I(N__8553));
    LocalMux I__1170 (
            .O(N__8566),
            .I(N__8547));
    LocalMux I__1169 (
            .O(N__8561),
            .I(N__8547));
    Span4Mux_h I__1168 (
            .O(N__8558),
            .I(N__8544));
    InMux I__1167 (
            .O(N__8557),
            .I(N__8535));
    InMux I__1166 (
            .O(N__8556),
            .I(N__8535));
    InMux I__1165 (
            .O(N__8553),
            .I(N__8535));
    InMux I__1164 (
            .O(N__8552),
            .I(N__8535));
    Odrv4 I__1163 (
            .O(N__8547),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    Odrv4 I__1162 (
            .O(N__8544),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__1161 (
            .O(N__8535),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    CascadeMux I__1160 (
            .O(N__8528),
            .I(beamY_RNIB6AOI5_0Z0Z_5_cascade_));
    InMux I__1159 (
            .O(N__8525),
            .I(N__8518));
    InMux I__1158 (
            .O(N__8524),
            .I(N__8509));
    InMux I__1157 (
            .O(N__8523),
            .I(N__8509));
    InMux I__1156 (
            .O(N__8522),
            .I(N__8509));
    InMux I__1155 (
            .O(N__8521),
            .I(N__8509));
    LocalMux I__1154 (
            .O(N__8518),
            .I(N__8506));
    LocalMux I__1153 (
            .O(N__8509),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    Odrv4 I__1152 (
            .O(N__8506),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    InMux I__1151 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__1150 (
            .O(N__8498),
            .I(N__8495));
    Span4Mux_v I__1149 (
            .O(N__8495),
            .I(N__8492));
    Odrv4 I__1148 (
            .O(N__8492),
            .I(un5_visibley_c2));
    CascadeMux I__1147 (
            .O(N__8489),
            .I(N__8483));
    CascadeMux I__1146 (
            .O(N__8488),
            .I(N__8476));
    CascadeMux I__1145 (
            .O(N__8487),
            .I(N__8472));
    CascadeMux I__1144 (
            .O(N__8486),
            .I(N__8468));
    InMux I__1143 (
            .O(N__8483),
            .I(N__8465));
    InMux I__1142 (
            .O(N__8482),
            .I(N__8458));
    InMux I__1141 (
            .O(N__8481),
            .I(N__8455));
    InMux I__1140 (
            .O(N__8480),
            .I(N__8448));
    InMux I__1139 (
            .O(N__8479),
            .I(N__8448));
    InMux I__1138 (
            .O(N__8476),
            .I(N__8448));
    InMux I__1137 (
            .O(N__8475),
            .I(N__8443));
    InMux I__1136 (
            .O(N__8472),
            .I(N__8443));
    InMux I__1135 (
            .O(N__8471),
            .I(N__8440));
    InMux I__1134 (
            .O(N__8468),
            .I(N__8437));
    LocalMux I__1133 (
            .O(N__8465),
            .I(N__8434));
    InMux I__1132 (
            .O(N__8464),
            .I(N__8429));
    InMux I__1131 (
            .O(N__8463),
            .I(N__8429));
    InMux I__1130 (
            .O(N__8462),
            .I(N__8426));
    InMux I__1129 (
            .O(N__8461),
            .I(N__8423));
    LocalMux I__1128 (
            .O(N__8458),
            .I(N__8420));
    LocalMux I__1127 (
            .O(N__8455),
            .I(N__8417));
    LocalMux I__1126 (
            .O(N__8448),
            .I(N__8414));
    LocalMux I__1125 (
            .O(N__8443),
            .I(N__8411));
    LocalMux I__1124 (
            .O(N__8440),
            .I(N__8404));
    LocalMux I__1123 (
            .O(N__8437),
            .I(N__8404));
    Span4Mux_s3_h I__1122 (
            .O(N__8434),
            .I(N__8404));
    LocalMux I__1121 (
            .O(N__8429),
            .I(N__8401));
    LocalMux I__1120 (
            .O(N__8426),
            .I(N__8398));
    LocalMux I__1119 (
            .O(N__8423),
            .I(N__8395));
    Span4Mux_s3_h I__1118 (
            .O(N__8420),
            .I(N__8392));
    Span4Mux_s3_h I__1117 (
            .O(N__8417),
            .I(N__8389));
    Span4Mux_v I__1116 (
            .O(N__8414),
            .I(N__8386));
    Span12Mux_s3_h I__1115 (
            .O(N__8411),
            .I(N__8383));
    Span4Mux_v I__1114 (
            .O(N__8404),
            .I(N__8378));
    Span4Mux_s3_h I__1113 (
            .O(N__8401),
            .I(N__8378));
    Span12Mux_s10_v I__1112 (
            .O(N__8398),
            .I(N__8375));
    Span4Mux_s3_h I__1111 (
            .O(N__8395),
            .I(N__8370));
    Span4Mux_v I__1110 (
            .O(N__8392),
            .I(N__8370));
    Odrv4 I__1109 (
            .O(N__8389),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1108 (
            .O(N__8386),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv12 I__1107 (
            .O(N__8383),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1106 (
            .O(N__8378),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv12 I__1105 (
            .O(N__8375),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1104 (
            .O(N__8370),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    InMux I__1103 (
            .O(N__8357),
            .I(N__8351));
    InMux I__1102 (
            .O(N__8356),
            .I(N__8351));
    LocalMux I__1101 (
            .O(N__8351),
            .I(row_1_if_generate_plus_mult1_un75_sum_c5));
    CascadeMux I__1100 (
            .O(N__8348),
            .I(if_generate_plus_mult1_un82_sum_axb4_x1_cascade_));
    InMux I__1099 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__1098 (
            .O(N__8342),
            .I(if_generate_plus_mult1_un82_sum_axb4_x0));
    InMux I__1097 (
            .O(N__8339),
            .I(N__8336));
    LocalMux I__1096 (
            .O(N__8336),
            .I(N__8333));
    Span4Mux_s1_h I__1095 (
            .O(N__8333),
            .I(N__8330));
    Odrv4 I__1094 (
            .O(N__8330),
            .I(beamY_RNIP8FF1_0Z0Z_7));
    CascadeMux I__1093 (
            .O(N__8327),
            .I(un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_));
    CascadeMux I__1092 (
            .O(N__8324),
            .I(un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_));
    CascadeMux I__1091 (
            .O(N__8321),
            .I(beamY_RNIP8FF1Z0Z_7_cascade_));
    InMux I__1090 (
            .O(N__8318),
            .I(N__8312));
    InMux I__1089 (
            .O(N__8317),
            .I(N__8308));
    InMux I__1088 (
            .O(N__8316),
            .I(N__8303));
    InMux I__1087 (
            .O(N__8315),
            .I(N__8300));
    LocalMux I__1086 (
            .O(N__8312),
            .I(N__8297));
    InMux I__1085 (
            .O(N__8311),
            .I(N__8294));
    LocalMux I__1084 (
            .O(N__8308),
            .I(N__8291));
    InMux I__1083 (
            .O(N__8307),
            .I(N__8286));
    InMux I__1082 (
            .O(N__8306),
            .I(N__8286));
    LocalMux I__1081 (
            .O(N__8303),
            .I(N__8279));
    LocalMux I__1080 (
            .O(N__8300),
            .I(N__8279));
    Span4Mux_h I__1079 (
            .O(N__8297),
            .I(N__8279));
    LocalMux I__1078 (
            .O(N__8294),
            .I(un5_visibley_c6));
    Odrv4 I__1077 (
            .O(N__8291),
            .I(un5_visibley_c6));
    LocalMux I__1076 (
            .O(N__8286),
            .I(un5_visibley_c6));
    Odrv4 I__1075 (
            .O(N__8279),
            .I(un5_visibley_c6));
    InMux I__1074 (
            .O(N__8270),
            .I(N__8264));
    InMux I__1073 (
            .O(N__8269),
            .I(N__8264));
    LocalMux I__1072 (
            .O(N__8264),
            .I(N__8260));
    InMux I__1071 (
            .O(N__8263),
            .I(N__8257));
    IoSpan4Mux I__1070 (
            .O(N__8260),
            .I(N__8252));
    LocalMux I__1069 (
            .O(N__8257),
            .I(N__8252));
    Span4Mux_s3_h I__1068 (
            .O(N__8252),
            .I(N__8249));
    Odrv4 I__1067 (
            .O(N__8249),
            .I(chary_if_generate_plus_mult1_un40_sum_c4));
    InMux I__1066 (
            .O(N__8246),
            .I(N__8243));
    LocalMux I__1065 (
            .O(N__8243),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1));
    CascadeMux I__1064 (
            .O(N__8240),
            .I(row_1_if_i4_mux_i_cascade_));
    InMux I__1063 (
            .O(N__8237),
            .I(N__8230));
    InMux I__1062 (
            .O(N__8236),
            .I(N__8225));
    InMux I__1061 (
            .O(N__8235),
            .I(N__8225));
    InMux I__1060 (
            .O(N__8234),
            .I(N__8220));
    InMux I__1059 (
            .O(N__8233),
            .I(N__8220));
    LocalMux I__1058 (
            .O(N__8230),
            .I(N__8215));
    LocalMux I__1057 (
            .O(N__8225),
            .I(N__8215));
    LocalMux I__1056 (
            .O(N__8220),
            .I(N__8212));
    Span4Mux_v I__1055 (
            .O(N__8215),
            .I(N__8209));
    Odrv4 I__1054 (
            .O(N__8212),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3));
    Odrv4 I__1053 (
            .O(N__8209),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3));
    InMux I__1052 (
            .O(N__8204),
            .I(N__8201));
    LocalMux I__1051 (
            .O(N__8201),
            .I(row_1_if_i4_mux_i));
    CascadeMux I__1050 (
            .O(N__8198),
            .I(row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_));
    InMux I__1049 (
            .O(N__8195),
            .I(N__8192));
    LocalMux I__1048 (
            .O(N__8192),
            .I(row_1_if_N_6));
    CascadeMux I__1047 (
            .O(N__8189),
            .I(if_generate_plus_mult1_un75_sum_axbxc3_cascade_));
    InMux I__1046 (
            .O(N__8186),
            .I(N__8182));
    InMux I__1045 (
            .O(N__8185),
            .I(N__8179));
    LocalMux I__1044 (
            .O(N__8182),
            .I(N__8176));
    LocalMux I__1043 (
            .O(N__8179),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0));
    Odrv4 I__1042 (
            .O(N__8176),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0));
    CascadeMux I__1041 (
            .O(N__8171),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_));
    CascadeMux I__1040 (
            .O(N__8168),
            .I(N__8165));
    InMux I__1039 (
            .O(N__8165),
            .I(N__8160));
    InMux I__1038 (
            .O(N__8164),
            .I(N__8155));
    InMux I__1037 (
            .O(N__8163),
            .I(N__8155));
    LocalMux I__1036 (
            .O(N__8160),
            .I(N__8150));
    LocalMux I__1035 (
            .O(N__8155),
            .I(N__8150));
    Odrv4 I__1034 (
            .O(N__8150),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0));
    InMux I__1033 (
            .O(N__8147),
            .I(N__8144));
    LocalMux I__1032 (
            .O(N__8144),
            .I(if_generate_plus_mult1_un75_sum_axbxc3));
    InMux I__1031 (
            .O(N__8141),
            .I(N__8138));
    LocalMux I__1030 (
            .O(N__8138),
            .I(N__8134));
    InMux I__1029 (
            .O(N__8137),
            .I(N__8131));
    Span4Mux_v I__1028 (
            .O(N__8134),
            .I(N__8128));
    LocalMux I__1027 (
            .O(N__8131),
            .I(N__8125));
    Odrv4 I__1026 (
            .O(N__8128),
            .I(un21_beamy_cry_7_c_RNIM7EZ0Z3));
    Odrv12 I__1025 (
            .O(N__8125),
            .I(un21_beamy_cry_7_c_RNIM7EZ0Z3));
    InMux I__1024 (
            .O(N__8120),
            .I(un21_beamy_cry_7));
    InMux I__1023 (
            .O(N__8117),
            .I(bfn_2_13_0_));
    CascadeMux I__1022 (
            .O(N__8114),
            .I(if_generate_plus_mult1_un61_sum_axbxc5_cascade_));
    CascadeMux I__1021 (
            .O(N__8111),
            .I(N__8107));
    InMux I__1020 (
            .O(N__8110),
            .I(N__8104));
    InMux I__1019 (
            .O(N__8107),
            .I(N__8101));
    LocalMux I__1018 (
            .O(N__8104),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5));
    LocalMux I__1017 (
            .O(N__8101),
            .I(row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5));
    CascadeMux I__1016 (
            .O(N__8096),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_));
    CascadeMux I__1015 (
            .O(N__8093),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5_cascade_));
    InMux I__1014 (
            .O(N__8090),
            .I(N__8084));
    InMux I__1013 (
            .O(N__8089),
            .I(N__8084));
    LocalMux I__1012 (
            .O(N__8084),
            .I(N__8081));
    Odrv12 I__1011 (
            .O(N__8081),
            .I(row_1_if_generate_plus_mult1_un61_sum_axb4_i));
    CascadeMux I__1010 (
            .O(N__8078),
            .I(N__8075));
    InMux I__1009 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__1008 (
            .O(N__8072),
            .I(N__8069));
    Odrv12 I__1007 (
            .O(N__8069),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6));
    InMux I__1006 (
            .O(N__8066),
            .I(N__8060));
    InMux I__1005 (
            .O(N__8065),
            .I(N__8060));
    LocalMux I__1004 (
            .O(N__8060),
            .I(N__8057));
    Odrv4 I__1003 (
            .O(N__8057),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    InMux I__1002 (
            .O(N__8054),
            .I(un21_beamy_cry_1));
    InMux I__1001 (
            .O(N__8051),
            .I(N__8048));
    LocalMux I__1000 (
            .O(N__8048),
            .I(N__8044));
    InMux I__999 (
            .O(N__8047),
            .I(N__8041));
    Span4Mux_v I__998 (
            .O(N__8044),
            .I(N__8038));
    LocalMux I__997 (
            .O(N__8041),
            .I(N__8035));
    Odrv4 I__996 (
            .O(N__8038),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    Odrv12 I__995 (
            .O(N__8035),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    InMux I__994 (
            .O(N__8030),
            .I(un21_beamy_cry_2));
    InMux I__993 (
            .O(N__8027),
            .I(N__8023));
    InMux I__992 (
            .O(N__8026),
            .I(N__8020));
    LocalMux I__991 (
            .O(N__8023),
            .I(N__8017));
    LocalMux I__990 (
            .O(N__8020),
            .I(N__8014));
    Odrv12 I__989 (
            .O(N__8017),
            .I(un21_beamy_cry_3_c_RNIERZ0Z93));
    Odrv4 I__988 (
            .O(N__8014),
            .I(un21_beamy_cry_3_c_RNIERZ0Z93));
    InMux I__987 (
            .O(N__8009),
            .I(un21_beamy_cry_3));
    InMux I__986 (
            .O(N__8006),
            .I(N__8003));
    LocalMux I__985 (
            .O(N__8003),
            .I(N__7999));
    InMux I__984 (
            .O(N__8002),
            .I(N__7996));
    Odrv12 I__983 (
            .O(N__7999),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    LocalMux I__982 (
            .O(N__7996),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    InMux I__981 (
            .O(N__7991),
            .I(un21_beamy_cry_4));
    InMux I__980 (
            .O(N__7988),
            .I(N__7985));
    LocalMux I__979 (
            .O(N__7985),
            .I(N__7981));
    InMux I__978 (
            .O(N__7984),
            .I(N__7978));
    Odrv12 I__977 (
            .O(N__7981),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    LocalMux I__976 (
            .O(N__7978),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    InMux I__975 (
            .O(N__7973),
            .I(un21_beamy_cry_5));
    CascadeMux I__974 (
            .O(N__7970),
            .I(N__7967));
    InMux I__973 (
            .O(N__7967),
            .I(N__7961));
    InMux I__972 (
            .O(N__7966),
            .I(N__7961));
    LocalMux I__971 (
            .O(N__7961),
            .I(N__7958));
    Odrv12 I__970 (
            .O(N__7958),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    InMux I__969 (
            .O(N__7955),
            .I(un21_beamy_cry_6));
    InMux I__968 (
            .O(N__7952),
            .I(N__7948));
    InMux I__967 (
            .O(N__7951),
            .I(N__7945));
    LocalMux I__966 (
            .O(N__7948),
            .I(beamY_fastZ0Z_7));
    LocalMux I__965 (
            .O(N__7945),
            .I(beamY_fastZ0Z_7));
    InMux I__964 (
            .O(N__7940),
            .I(N__7932));
    InMux I__963 (
            .O(N__7939),
            .I(N__7932));
    InMux I__962 (
            .O(N__7938),
            .I(N__7929));
    InMux I__961 (
            .O(N__7937),
            .I(N__7926));
    LocalMux I__960 (
            .O(N__7932),
            .I(beamY_fastZ0Z_6));
    LocalMux I__959 (
            .O(N__7929),
            .I(beamY_fastZ0Z_6));
    LocalMux I__958 (
            .O(N__7926),
            .I(beamY_fastZ0Z_6));
    InMux I__957 (
            .O(N__7919),
            .I(N__7910));
    InMux I__956 (
            .O(N__7918),
            .I(N__7910));
    InMux I__955 (
            .O(N__7917),
            .I(N__7910));
    LocalMux I__954 (
            .O(N__7910),
            .I(beamY_fastZ0Z_5));
    CascadeMux I__953 (
            .O(N__7907),
            .I(un5_visibley_ac0_11_0_1_cascade_));
    CascadeMux I__952 (
            .O(N__7904),
            .I(N__7900));
    InMux I__951 (
            .O(N__7903),
            .I(N__7896));
    InMux I__950 (
            .O(N__7900),
            .I(N__7891));
    InMux I__949 (
            .O(N__7899),
            .I(N__7891));
    LocalMux I__948 (
            .O(N__7896),
            .I(beamY_fastZ0Z_4));
    LocalMux I__947 (
            .O(N__7891),
            .I(beamY_fastZ0Z_4));
    CascadeMux I__946 (
            .O(N__7886),
            .I(N__7882));
    CascadeMux I__945 (
            .O(N__7885),
            .I(N__7879));
    InMux I__944 (
            .O(N__7882),
            .I(N__7874));
    InMux I__943 (
            .O(N__7879),
            .I(N__7874));
    LocalMux I__942 (
            .O(N__7874),
            .I(beamY_fastZ0Z_8));
    InMux I__941 (
            .O(N__7871),
            .I(N__7868));
    LocalMux I__940 (
            .O(N__7868),
            .I(un5_visibley_c7));
    InMux I__939 (
            .O(N__7865),
            .I(N__7862));
    LocalMux I__938 (
            .O(N__7862),
            .I(N__7856));
    InMux I__937 (
            .O(N__7861),
            .I(N__7853));
    InMux I__936 (
            .O(N__7860),
            .I(N__7850));
    InMux I__935 (
            .O(N__7859),
            .I(N__7847));
    Odrv4 I__934 (
            .O(N__7856),
            .I(beamY_fastZ0Z_3));
    LocalMux I__933 (
            .O(N__7853),
            .I(beamY_fastZ0Z_3));
    LocalMux I__932 (
            .O(N__7850),
            .I(beamY_fastZ0Z_3));
    LocalMux I__931 (
            .O(N__7847),
            .I(beamY_fastZ0Z_3));
    CascadeMux I__930 (
            .O(N__7838),
            .I(un5_visibley_c2_cascade_));
    InMux I__929 (
            .O(N__7835),
            .I(N__7829));
    InMux I__928 (
            .O(N__7834),
            .I(N__7826));
    InMux I__927 (
            .O(N__7833),
            .I(N__7821));
    InMux I__926 (
            .O(N__7832),
            .I(N__7821));
    LocalMux I__925 (
            .O(N__7829),
            .I(beamY_fastZ0Z_2));
    LocalMux I__924 (
            .O(N__7826),
            .I(beamY_fastZ0Z_2));
    LocalMux I__923 (
            .O(N__7821),
            .I(beamY_fastZ0Z_2));
    CascadeMux I__922 (
            .O(N__7814),
            .I(beamY_fast_RNIT5UFZ0Z_4_cascade_));
    InMux I__921 (
            .O(N__7811),
            .I(N__7808));
    LocalMux I__920 (
            .O(N__7808),
            .I(un5_visibley_ac0_7));
    CascadeMux I__919 (
            .O(N__7805),
            .I(un5_visibley_ac0_7_cascade_));
    CascadeMux I__918 (
            .O(N__7802),
            .I(N__7799));
    InMux I__917 (
            .O(N__7799),
            .I(N__7796));
    LocalMux I__916 (
            .O(N__7796),
            .I(N__7792));
    InMux I__915 (
            .O(N__7795),
            .I(N__7789));
    Odrv4 I__914 (
            .O(N__7792),
            .I(chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux));
    LocalMux I__913 (
            .O(N__7789),
            .I(chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux));
    InMux I__912 (
            .O(N__7784),
            .I(N__7781));
    LocalMux I__911 (
            .O(N__7781),
            .I(N__7778));
    Odrv4 I__910 (
            .O(N__7778),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0));
    CascadeMux I__909 (
            .O(N__7775),
            .I(N__7772));
    InMux I__908 (
            .O(N__7772),
            .I(N__7766));
    InMux I__907 (
            .O(N__7771),
            .I(N__7766));
    LocalMux I__906 (
            .O(N__7766),
            .I(N__7763));
    Span4Mux_v I__905 (
            .O(N__7763),
            .I(N__7760));
    Odrv4 I__904 (
            .O(N__7760),
            .I(chary_if_generate_plus_mult1_un47_sum_axb3));
    InMux I__903 (
            .O(N__7757),
            .I(N__7751));
    InMux I__902 (
            .O(N__7756),
            .I(N__7751));
    LocalMux I__901 (
            .O(N__7751),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0));
    InMux I__900 (
            .O(N__7748),
            .I(N__7742));
    InMux I__899 (
            .O(N__7747),
            .I(N__7742));
    LocalMux I__898 (
            .O(N__7742),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0));
    CascadeMux I__897 (
            .O(N__7739),
            .I(beamY_i_2_cascade_));
    CascadeMux I__896 (
            .O(N__7736),
            .I(N__7733));
    InMux I__895 (
            .O(N__7733),
            .I(N__7730));
    LocalMux I__894 (
            .O(N__7730),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0));
    CascadeMux I__893 (
            .O(N__7727),
            .I(N__7724));
    InMux I__892 (
            .O(N__7724),
            .I(N__7721));
    LocalMux I__891 (
            .O(N__7721),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1));
    InMux I__890 (
            .O(N__7718),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__889 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__888 (
            .O(N__7712),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1));
    CascadeMux I__887 (
            .O(N__7709),
            .I(N__7706));
    InMux I__886 (
            .O(N__7706),
            .I(N__7703));
    LocalMux I__885 (
            .O(N__7703),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1));
    InMux I__884 (
            .O(N__7700),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__883 (
            .O(N__7697),
            .I(N__7694));
    InMux I__882 (
            .O(N__7694),
            .I(N__7691));
    LocalMux I__881 (
            .O(N__7691),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1));
    InMux I__880 (
            .O(N__7688),
            .I(N__7685));
    LocalMux I__879 (
            .O(N__7685),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__878 (
            .O(N__7682),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__877 (
            .O(N__7679),
            .I(N__7674));
    InMux I__876 (
            .O(N__7678),
            .I(N__7669));
    InMux I__875 (
            .O(N__7677),
            .I(N__7669));
    LocalMux I__874 (
            .O(N__7674),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__873 (
            .O(N__7669),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    CascadeMux I__872 (
            .O(N__7664),
            .I(N__7661));
    InMux I__871 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__870 (
            .O(N__7658),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__869 (
            .O(N__7655),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__868 (
            .O(N__7652),
            .I(N__7647));
    CascadeMux I__867 (
            .O(N__7651),
            .I(N__7643));
    InMux I__866 (
            .O(N__7650),
            .I(N__7631));
    InMux I__865 (
            .O(N__7647),
            .I(N__7631));
    InMux I__864 (
            .O(N__7646),
            .I(N__7631));
    InMux I__863 (
            .O(N__7643),
            .I(N__7631));
    InMux I__862 (
            .O(N__7642),
            .I(N__7631));
    LocalMux I__861 (
            .O(N__7631),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9));
    InMux I__860 (
            .O(N__7628),
            .I(N__7625));
    LocalMux I__859 (
            .O(N__7625),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7));
    CascadeMux I__858 (
            .O(N__7622),
            .I(N__7618));
    InMux I__857 (
            .O(N__7621),
            .I(N__7608));
    InMux I__856 (
            .O(N__7618),
            .I(N__7608));
    InMux I__855 (
            .O(N__7617),
            .I(N__7608));
    InMux I__854 (
            .O(N__7616),
            .I(N__7603));
    InMux I__853 (
            .O(N__7615),
            .I(N__7603));
    LocalMux I__852 (
            .O(N__7608),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0));
    LocalMux I__851 (
            .O(N__7603),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0));
    InMux I__850 (
            .O(N__7598),
            .I(N__7595));
    LocalMux I__849 (
            .O(N__7595),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7));
    InMux I__848 (
            .O(N__7592),
            .I(N__7589));
    LocalMux I__847 (
            .O(N__7589),
            .I(N__7586));
    Odrv4 I__846 (
            .O(N__7586),
            .I(if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx));
    InMux I__845 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__844 (
            .O(N__7580),
            .I(beamY_RNIUUEM_0Z0Z_8));
    InMux I__843 (
            .O(N__7577),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__842 (
            .O(N__7574),
            .I(N__7571));
    LocalMux I__841 (
            .O(N__7571),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21));
    InMux I__840 (
            .O(N__7568),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__839 (
            .O(N__7565),
            .I(N__7562));
    LocalMux I__838 (
            .O(N__7562),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21));
    InMux I__837 (
            .O(N__7559),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__836 (
            .O(N__7556),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__835 (
            .O(N__7553),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__834 (
            .O(N__7550),
            .I(N__7544));
    InMux I__833 (
            .O(N__7549),
            .I(N__7544));
    LocalMux I__832 (
            .O(N__7544),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__831 (
            .O(N__7541),
            .I(N__7538));
    LocalMux I__830 (
            .O(N__7538),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0));
    InMux I__829 (
            .O(N__7535),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__828 (
            .O(N__7532),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_));
    InMux I__827 (
            .O(N__7529),
            .I(N__7526));
    LocalMux I__826 (
            .O(N__7526),
            .I(un114_pixel_6_1_5__g0Z0Z_2));
    InMux I__825 (
            .O(N__7523),
            .I(N__7517));
    InMux I__824 (
            .O(N__7522),
            .I(N__7517));
    LocalMux I__823 (
            .O(N__7517),
            .I(N__7514));
    Odrv4 I__822 (
            .O(N__7514),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0));
    CascadeMux I__821 (
            .O(N__7511),
            .I(chary_if_generate_plus_mult1_un61_sum_c4_cascade_));
    InMux I__820 (
            .O(N__7508),
            .I(N__7505));
    LocalMux I__819 (
            .O(N__7505),
            .I(N__7500));
    InMux I__818 (
            .O(N__7504),
            .I(N__7497));
    InMux I__817 (
            .O(N__7503),
            .I(N__7494));
    Odrv4 I__816 (
            .O(N__7500),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    LocalMux I__815 (
            .O(N__7497),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    LocalMux I__814 (
            .O(N__7494),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    CascadeMux I__813 (
            .O(N__7487),
            .I(beamY_RNISDTA58Z0Z_5_cascade_));
    InMux I__812 (
            .O(N__7484),
            .I(N__7481));
    LocalMux I__811 (
            .O(N__7481),
            .I(beamY_RNIJ0797KZ0Z_4));
    InMux I__810 (
            .O(N__7478),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__809 (
            .O(N__7475),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__808 (
            .O(N__7472),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__807 (
            .O(N__7469),
            .I(N__7466));
    LocalMux I__806 (
            .O(N__7466),
            .I(beamY_RNI2B511_0Z0Z_9));
    CascadeMux I__805 (
            .O(N__7463),
            .I(N__7460));
    InMux I__804 (
            .O(N__7460),
            .I(N__7457));
    LocalMux I__803 (
            .O(N__7457),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0));
    CascadeMux I__802 (
            .O(N__7454),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_));
    CascadeMux I__801 (
            .O(N__7451),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_));
    InMux I__800 (
            .O(N__7448),
            .I(N__7445));
    LocalMux I__799 (
            .O(N__7445),
            .I(g1_0_2));
    InMux I__798 (
            .O(N__7442),
            .I(N__7436));
    InMux I__797 (
            .O(N__7441),
            .I(N__7436));
    LocalMux I__796 (
            .O(N__7436),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    CascadeMux I__795 (
            .O(N__7433),
            .I(N__7430));
    InMux I__794 (
            .O(N__7430),
            .I(N__7427));
    LocalMux I__793 (
            .O(N__7427),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_0));
    InMux I__792 (
            .O(N__7424),
            .I(N__7421));
    LocalMux I__791 (
            .O(N__7421),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4_i_0));
    InMux I__790 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__789 (
            .O(N__7415),
            .I(g1_1));
    CascadeMux I__788 (
            .O(N__7412),
            .I(g2_0_cascade_));
    CascadeMux I__787 (
            .O(N__7409),
            .I(beamY_RNIV5SUC3_0Z0Z_9_cascade_));
    CascadeMux I__786 (
            .O(N__7406),
            .I(N__7403));
    InMux I__785 (
            .O(N__7403),
            .I(N__7400));
    LocalMux I__784 (
            .O(N__7400),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0_1));
    CascadeMux I__783 (
            .O(N__7397),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_));
    InMux I__782 (
            .O(N__7394),
            .I(N__7385));
    InMux I__781 (
            .O(N__7393),
            .I(N__7385));
    InMux I__780 (
            .O(N__7392),
            .I(N__7382));
    InMux I__779 (
            .O(N__7391),
            .I(N__7377));
    InMux I__778 (
            .O(N__7390),
            .I(N__7377));
    LocalMux I__777 (
            .O(N__7385),
            .I(beamY_RNIVADQVZ0Z_8));
    LocalMux I__776 (
            .O(N__7382),
            .I(beamY_RNIVADQVZ0Z_8));
    LocalMux I__775 (
            .O(N__7377),
            .I(beamY_RNIVADQVZ0Z_8));
    CascadeMux I__774 (
            .O(N__7370),
            .I(N__7364));
    CascadeMux I__773 (
            .O(N__7369),
            .I(N__7361));
    CascadeMux I__772 (
            .O(N__7368),
            .I(N__7357));
    InMux I__771 (
            .O(N__7367),
            .I(N__7350));
    InMux I__770 (
            .O(N__7364),
            .I(N__7350));
    InMux I__769 (
            .O(N__7361),
            .I(N__7350));
    InMux I__768 (
            .O(N__7360),
            .I(N__7345));
    InMux I__767 (
            .O(N__7357),
            .I(N__7345));
    LocalMux I__766 (
            .O(N__7350),
            .I(N__7342));
    LocalMux I__765 (
            .O(N__7345),
            .I(N__7339));
    Odrv12 I__764 (
            .O(N__7342),
            .I(chary_if_generate_plus_mult1_un47_sum_c4));
    Odrv4 I__763 (
            .O(N__7339),
            .I(chary_if_generate_plus_mult1_un47_sum_c4));
    CascadeMux I__762 (
            .O(N__7334),
            .I(N__7327));
    InMux I__761 (
            .O(N__7333),
            .I(N__7319));
    InMux I__760 (
            .O(N__7332),
            .I(N__7319));
    InMux I__759 (
            .O(N__7331),
            .I(N__7319));
    InMux I__758 (
            .O(N__7330),
            .I(N__7312));
    InMux I__757 (
            .O(N__7327),
            .I(N__7312));
    InMux I__756 (
            .O(N__7326),
            .I(N__7312));
    LocalMux I__755 (
            .O(N__7319),
            .I(N__7308));
    LocalMux I__754 (
            .O(N__7312),
            .I(N__7305));
    InMux I__753 (
            .O(N__7311),
            .I(N__7302));
    Odrv12 I__752 (
            .O(N__7308),
            .I(chary_if_generate_plus_mult1_un47_sum_axb4));
    Odrv4 I__751 (
            .O(N__7305),
            .I(chary_if_generate_plus_mult1_un47_sum_axb4));
    LocalMux I__750 (
            .O(N__7302),
            .I(chary_if_generate_plus_mult1_un47_sum_axb4));
    InMux I__749 (
            .O(N__7295),
            .I(N__7292));
    LocalMux I__748 (
            .O(N__7292),
            .I(beamY_RNIV5SUC3Z0Z_9));
    CascadeMux I__747 (
            .O(N__7289),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_));
    InMux I__746 (
            .O(N__7286),
            .I(N__7283));
    LocalMux I__745 (
            .O(N__7283),
            .I(beamY_RNIP8FF1_1Z0Z_7));
    InMux I__744 (
            .O(N__7280),
            .I(N__7275));
    CascadeMux I__743 (
            .O(N__7279),
            .I(N__7271));
    CascadeMux I__742 (
            .O(N__7278),
            .I(N__7265));
    LocalMux I__741 (
            .O(N__7275),
            .I(N__7262));
    InMux I__740 (
            .O(N__7274),
            .I(N__7257));
    InMux I__739 (
            .O(N__7271),
            .I(N__7257));
    InMux I__738 (
            .O(N__7270),
            .I(N__7254));
    InMux I__737 (
            .O(N__7269),
            .I(N__7249));
    InMux I__736 (
            .O(N__7268),
            .I(N__7249));
    InMux I__735 (
            .O(N__7265),
            .I(N__7246));
    Odrv4 I__734 (
            .O(N__7262),
            .I(beamY_RNI93821Z0Z_9));
    LocalMux I__733 (
            .O(N__7257),
            .I(beamY_RNI93821Z0Z_9));
    LocalMux I__732 (
            .O(N__7254),
            .I(beamY_RNI93821Z0Z_9));
    LocalMux I__731 (
            .O(N__7249),
            .I(beamY_RNI93821Z0Z_9));
    LocalMux I__730 (
            .O(N__7246),
            .I(beamY_RNI93821Z0Z_9));
    CascadeMux I__729 (
            .O(N__7235),
            .I(beamY_RNIBV5E51Z0Z_8_cascade_));
    InMux I__728 (
            .O(N__7232),
            .I(N__7229));
    LocalMux I__727 (
            .O(N__7229),
            .I(beamY_RNIBV5E51_0Z0Z_8));
    InMux I__726 (
            .O(N__7226),
            .I(N__7216));
    InMux I__725 (
            .O(N__7225),
            .I(N__7216));
    InMux I__724 (
            .O(N__7224),
            .I(N__7216));
    InMux I__723 (
            .O(N__7223),
            .I(N__7213));
    LocalMux I__722 (
            .O(N__7216),
            .I(N__7208));
    LocalMux I__721 (
            .O(N__7213),
            .I(N__7208));
    Odrv4 I__720 (
            .O(N__7208),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_2));
    CascadeMux I__719 (
            .O(N__7205),
            .I(N__7200));
    InMux I__718 (
            .O(N__7204),
            .I(N__7190));
    InMux I__717 (
            .O(N__7203),
            .I(N__7190));
    InMux I__716 (
            .O(N__7200),
            .I(N__7190));
    InMux I__715 (
            .O(N__7199),
            .I(N__7190));
    LocalMux I__714 (
            .O(N__7190),
            .I(N__7186));
    InMux I__713 (
            .O(N__7189),
            .I(N__7183));
    Odrv4 I__712 (
            .O(N__7186),
            .I(chary_if_generate_plus_mult1_un47_sum_c5));
    LocalMux I__711 (
            .O(N__7183),
            .I(chary_if_generate_plus_mult1_un47_sum_c5));
    CascadeMux I__710 (
            .O(N__7178),
            .I(beamY_RNIVADQVZ0Z_8_cascade_));
    InMux I__709 (
            .O(N__7175),
            .I(N__7169));
    InMux I__708 (
            .O(N__7174),
            .I(N__7169));
    LocalMux I__707 (
            .O(N__7169),
            .I(chary_if_generate_plus_mult1_un54_sum_ac0_5));
    CascadeMux I__706 (
            .O(N__7166),
            .I(beamY_RNI93821Z0Z_9_cascade_));
    InMux I__705 (
            .O(N__7163),
            .I(N__7160));
    LocalMux I__704 (
            .O(N__7160),
            .I(beamY_RNIM5433_0Z0Z_8));
    InMux I__703 (
            .O(N__7157),
            .I(N__7154));
    LocalMux I__702 (
            .O(N__7154),
            .I(beamY_RNIIR4K3_0Z0Z_7));
    CascadeMux I__701 (
            .O(N__7151),
            .I(beamY_RNIIR4K3_0Z0Z_7_cascade_));
    InMux I__700 (
            .O(N__7148),
            .I(N__7145));
    LocalMux I__699 (
            .O(N__7145),
            .I(beamY_RNIKM9GC_0Z0Z_9));
    CascadeMux I__698 (
            .O(N__7142),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_));
    InMux I__697 (
            .O(N__7139),
            .I(N__7136));
    LocalMux I__696 (
            .O(N__7136),
            .I(N__7133));
    Odrv12 I__695 (
            .O(N__7133),
            .I(beamY_RNI9DSP2_0Z0Z_8));
    CascadeMux I__694 (
            .O(N__7130),
            .I(beamY_RNI41384Z0Z_7_cascade_));
    CascadeMux I__693 (
            .O(N__7127),
            .I(chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_));
    CascadeMux I__692 (
            .O(N__7124),
            .I(un8_beamylt9_0_cascade_));
    CascadeMux I__691 (
            .O(N__7121),
            .I(N__7118));
    InMux I__690 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__689 (
            .O(N__7115),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0));
    CascadeMux I__688 (
            .O(N__7112),
            .I(N__7107));
    CascadeMux I__687 (
            .O(N__7111),
            .I(N__7103));
    InMux I__686 (
            .O(N__7110),
            .I(N__7099));
    InMux I__685 (
            .O(N__7107),
            .I(N__7090));
    InMux I__684 (
            .O(N__7106),
            .I(N__7090));
    InMux I__683 (
            .O(N__7103),
            .I(N__7090));
    InMux I__682 (
            .O(N__7102),
            .I(N__7090));
    LocalMux I__681 (
            .O(N__7099),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0));
    LocalMux I__680 (
            .O(N__7090),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0));
    InMux I__679 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__678 (
            .O(N__7082),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__677 (
            .O(N__7079),
            .I(N__7076));
    LocalMux I__676 (
            .O(N__7076),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__675 (
            .O(N__7073),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__674 (
            .O(N__7070),
            .I(N__7067));
    LocalMux I__673 (
            .O(N__7067),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0));
    CascadeMux I__672 (
            .O(N__7064),
            .I(chary_if_generate_plus_mult1_un47_sum_axb4_cascade_));
    CascadeMux I__671 (
            .O(N__7061),
            .I(beamY_RNIKM9GCZ0Z_9_cascade_));
    InMux I__670 (
            .O(N__7058),
            .I(N__7055));
    LocalMux I__669 (
            .O(N__7055),
            .I(beamY_RNIM5433Z0Z_8));
    CascadeMux I__668 (
            .O(N__7052),
            .I(N__7049));
    InMux I__667 (
            .O(N__7049),
            .I(N__7046));
    LocalMux I__666 (
            .O(N__7046),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3));
    InMux I__665 (
            .O(N__7043),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__664 (
            .O(N__7040),
            .I(N__7037));
    InMux I__663 (
            .O(N__7037),
            .I(N__7034));
    LocalMux I__662 (
            .O(N__7034),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4));
    InMux I__661 (
            .O(N__7031),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__660 (
            .O(N__7028),
            .I(N__7025));
    LocalMux I__659 (
            .O(N__7025),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__658 (
            .O(N__7022),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__657 (
            .O(N__7019),
            .I(N__7014));
    InMux I__656 (
            .O(N__7018),
            .I(N__7009));
    InMux I__655 (
            .O(N__7017),
            .I(N__7000));
    InMux I__654 (
            .O(N__7014),
            .I(N__7000));
    InMux I__653 (
            .O(N__7013),
            .I(N__7000));
    InMux I__652 (
            .O(N__7012),
            .I(N__7000));
    LocalMux I__651 (
            .O(N__7009),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5));
    LocalMux I__650 (
            .O(N__7000),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5));
    InMux I__649 (
            .O(N__6995),
            .I(N__6992));
    LocalMux I__648 (
            .O(N__6992),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__647 (
            .O(N__6989),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__646 (
            .O(N__6986),
            .I(N__6983));
    InMux I__645 (
            .O(N__6983),
            .I(N__6980));
    LocalMux I__644 (
            .O(N__6980),
            .I(N__6977));
    Odrv4 I__643 (
            .O(N__6977),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6));
    InMux I__642 (
            .O(N__6974),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__641 (
            .O(N__6971),
            .I(N__6968));
    LocalMux I__640 (
            .O(N__6968),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9));
    InMux I__639 (
            .O(N__6965),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__638 (
            .O(N__6962),
            .I(N__6958));
    InMux I__637 (
            .O(N__6961),
            .I(N__6949));
    InMux I__636 (
            .O(N__6958),
            .I(N__6949));
    InMux I__635 (
            .O(N__6957),
            .I(N__6949));
    InMux I__634 (
            .O(N__6956),
            .I(N__6946));
    LocalMux I__633 (
            .O(N__6949),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2));
    LocalMux I__632 (
            .O(N__6946),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2));
    CascadeMux I__631 (
            .O(N__6941),
            .I(N__6938));
    InMux I__630 (
            .O(N__6938),
            .I(N__6935));
    LocalMux I__629 (
            .O(N__6935),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1));
    InMux I__628 (
            .O(N__6932),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__627 (
            .O(N__6929),
            .I(N__6926));
    LocalMux I__626 (
            .O(N__6926),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85));
    CascadeMux I__625 (
            .O(N__6923),
            .I(N__6919));
    InMux I__624 (
            .O(N__6922),
            .I(N__6916));
    InMux I__623 (
            .O(N__6919),
            .I(N__6913));
    LocalMux I__622 (
            .O(N__6916),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2));
    LocalMux I__621 (
            .O(N__6913),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2));
    InMux I__620 (
            .O(N__6908),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__619 (
            .O(N__6905),
            .I(N__6902));
    LocalMux I__618 (
            .O(N__6902),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__617 (
            .O(N__6899),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__616 (
            .O(N__6896),
            .I(N__6893));
    InMux I__615 (
            .O(N__6893),
            .I(N__6890));
    LocalMux I__614 (
            .O(N__6890),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0));
    CascadeMux I__613 (
            .O(N__6887),
            .I(N__6884));
    InMux I__612 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__611 (
            .O(N__6881),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__610 (
            .O(N__6878),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__609 (
            .O(N__6875),
            .I(N__6872));
    LocalMux I__608 (
            .O(N__6872),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3));
    InMux I__607 (
            .O(N__6869),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__606 (
            .O(N__6866),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__605 (
            .O(N__6863),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__604 (
            .O(N__6860),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__603 (
            .O(N__6857),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__602 (
            .O(N__6854),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_));
    InMux I__601 (
            .O(N__6851),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__600 (
            .O(N__6848),
            .I(N__6845));
    LocalMux I__599 (
            .O(N__6845),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0));
    InMux I__598 (
            .O(N__6842),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    IoInMux I__597 (
            .O(N__6839),
            .I(N__6836));
    LocalMux I__596 (
            .O(N__6836),
            .I(N__6833));
    IoSpan4Mux I__595 (
            .O(N__6833),
            .I(N__6830));
    Odrv4 I__594 (
            .O(N__6830),
            .I(Clock12MHz_c));
    IoInMux I__593 (
            .O(N__6827),
            .I(N__6824));
    LocalMux I__592 (
            .O(N__6824),
            .I(N__6821));
    IoSpan4Mux I__591 (
            .O(N__6821),
            .I(N__6818));
    IoSpan4Mux I__590 (
            .O(N__6818),
            .I(N__6815));
    IoSpan4Mux I__589 (
            .O(N__6815),
            .I(N__6812));
    Odrv4 I__588 (
            .O(N__6812),
            .I(\Clock50MHz.PixelClock ));
    CascadeMux I__587 (
            .O(N__6809),
            .I(N__6806));
    InMux I__586 (
            .O(N__6806),
            .I(N__6803));
    LocalMux I__585 (
            .O(N__6803),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__584 (
            .O(N__6800),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__6827),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_3_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_3_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8462),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(N__9116),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_1_4_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_1_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_1_4_1 (
            .in0(_gnd_net_),
            .in1(N__7617),
            .in2(N__6809),
            .in3(N__6800),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_1_4_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_1_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_1_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_1_4_2 (
            .in0(_gnd_net_),
            .in1(N__7541),
            .in2(N__7622),
            .in3(N__6866),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68E2_LC_1_4_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68E2_LC_1_4_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68E2_LC_1_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68E2_LC_1_4_3 (
            .in0(_gnd_net_),
            .in1(N__7621),
            .in2(N__7727),
            .in3(N__6863),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC29L5_LC_1_4_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC29L5_LC_1_4_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC29L5_LC_1_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC29L5_LC_1_4_4 (
            .in0(N__6956),
            .in1(N__7598),
            .in2(N__7709),
            .in3(N__6860),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQ2_LC_1_4_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQ2_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQ2_LC_1_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQ2_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(N__7688),
            .in2(_gnd_net_),
            .in3(N__6857),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRU85_LC_1_4_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRU85_LC_1_4_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRU85_LC_1_4_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRU85_LC_1_4_6 (
            .in0(N__6922),
            .in1(_gnd_net_),
            .in2(N__6854),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUUEM_0_8_LC_1_4_7.C_ON=1'b0;
    defparam beamY_RNIUUEM_0_8_LC_1_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIUUEM_0_8_LC_1_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 beamY_RNIUUEM_0_8_LC_1_4_7 (
            .in0(N__12168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_RNIUUEM_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_5_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_5_0 (
            .in0(_gnd_net_),
            .in1(N__10239),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDC3_LC_1_5_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDC3_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDC3_LC_1_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDC3_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__6957),
            .in2(N__6896),
            .in3(N__6851),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PU3_LC_1_5_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PU3_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PU3_LC_1_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PU3_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(N__6848),
            .in2(N__6962),
            .in3(N__6842),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJ4_LC_1_5_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJ4_LC_1_5_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJ4_LC_1_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJ4_LC_1_5_3 (
            .in0(_gnd_net_),
            .in1(N__6961),
            .in2(N__6941),
            .in3(N__6932),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINP5QD_LC_1_5_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINP5QD_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINP5QD_LC_1_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINP5QD_LC_1_5_4 (
            .in0(N__7018),
            .in1(N__6929),
            .in2(N__6923),
            .in3(N__6908),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_LC_1_5_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_LC_1_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_LC_1_5_5 (
            .in0(_gnd_net_),
            .in1(N__6905),
            .in2(_gnd_net_),
            .in3(N__6899),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_5_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9104),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_5_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_5_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_5_7 (
            .in0(N__10240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_6_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(N__10090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8A6_LC_1_6_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8A6_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8A6_LC_1_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8A6_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(N__7013),
            .in2(N__6887),
            .in3(N__6878),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RH9_LC_1_6_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RH9_LC_1_6_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RH9_LC_1_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RH9_LC_1_6_2 (
            .in0(_gnd_net_),
            .in1(N__6875),
            .in2(N__7019),
            .in3(N__6869),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74A_LC_1_6_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74A_LC_1_6_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74A_LC_1_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74A_LC_1_6_3 (
            .in0(_gnd_net_),
            .in1(N__7017),
            .in2(N__7052),
            .in3(N__7043),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIQGGSO_LC_1_6_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIQGGSO_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIQGGSO_LC_1_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIQGGSO_LC_1_6_4 (
            .in0(N__7110),
            .in1(N__6995),
            .in2(N__7040),
            .in3(N__7031),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3E_LC_1_6_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3E_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3E_LC_1_6_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3E_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(N__7028),
            .in2(_gnd_net_),
            .in3(N__7022),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUUEM_8_LC_1_6_6.C_ON=1'b0;
    defparam beamY_RNIUUEM_8_LC_1_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIUUEM_8_LC_1_6_6.LUT_INIT=16'b1010101001010101;
    LogicCell40 beamY_RNIUUEM_8_LC_1_6_6 (
            .in0(N__8315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9261),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_0_LC_1_6_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_0_LC_1_6_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_0_LC_1_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_0_LC_1_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7012),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_7_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_7_0 (
            .in0(_gnd_net_),
            .in1(N__10946),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NE_LC_1_7_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NE_LC_1_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NE_LC_1_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NE_LC_1_7_1 (
            .in0(_gnd_net_),
            .in1(N__7070),
            .in2(N__7111),
            .in3(N__6989),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATK_LC_1_7_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATK_LC_1_7_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATK_LC_1_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATK_LC_1_7_2 (
            .in0(_gnd_net_),
            .in1(N__7106),
            .in2(N__6986),
            .in3(N__6974),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4O_LC_1_7_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4O_LC_1_7_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4O_LC_1_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4O_LC_1_7_3 (
            .in0(_gnd_net_),
            .in1(N__6971),
            .in2(N__7112),
            .in3(N__6965),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_1_7_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_1_7_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_1_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_1_7_4 (
            .in0(_gnd_net_),
            .in1(N__7085),
            .in2(N__7121),
            .in3(N__7102),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CP_LC_1_7_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CP_LC_1_7_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CP_LC_1_7_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CP_LC_1_7_5 (
            .in0(_gnd_net_),
            .in1(N__7079),
            .in2(_gnd_net_),
            .in3(N__7073),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DSP2_0_8_LC_1_7_6.C_ON=1'b0;
    defparam beamY_RNI9DSP2_0_8_LC_1_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DSP2_0_8_LC_1_7_6.LUT_INIT=16'b0000011011111001;
    LogicCell40 beamY_RNI9DSP2_0_8_LC_1_7_6 (
            .in0(N__9295),
            .in1(N__8316),
            .in2(N__12112),
            .in3(N__7270),
            .lcout(beamY_RNI9DSP2_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_1_7_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_1_7_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_1_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_1_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10104),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICLER6_8_LC_1_8_0.C_ON=1'b0;
    defparam beamY_RNICLER6_8_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam beamY_RNICLER6_8_LC_1_8_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 beamY_RNICLER6_8_LC_1_8_0 (
            .in0(N__7163),
            .in1(N__7058),
            .in2(_gnd_net_),
            .in3(N__8306),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axb4),
            .ltout(chary_if_generate_plus_mult1_un47_sum_axb4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKM9GC_9_LC_1_8_1.C_ON=1'b0;
    defparam beamY_RNIKM9GC_9_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIKM9GC_9_LC_1_8_1.LUT_INIT=16'b1111001111010000;
    LogicCell40 beamY_RNIKM9GC_9_LC_1_8_1 (
            .in0(N__12236),
            .in1(N__7269),
            .in2(N__7064),
            .in3(N__7157),
            .lcout(),
            .ltout(beamY_RNIKM9GCZ0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI42CCP_5_LC_1_8_2.C_ON=1'b0;
    defparam beamY_RNI42CCP_5_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI42CCP_5_LC_1_8_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 beamY_RNI42CCP_5_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(N__7148),
            .in2(N__7061),
            .in3(N__8461),
            .lcout(chary_if_generate_plus_mult1_un47_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM5433_8_LC_1_8_3.C_ON=1'b0;
    defparam beamY_RNIM5433_8_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIM5433_8_LC_1_8_3.LUT_INIT=16'b1010010110010110;
    LogicCell40 beamY_RNIM5433_8_LC_1_8_3 (
            .in0(N__12233),
            .in1(N__9298),
            .in2(N__7278),
            .in3(N__12059),
            .lcout(beamY_RNIM5433Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI93821_9_LC_1_8_4.C_ON=1'b0;
    defparam beamY_RNI93821_9_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI93821_9_LC_1_8_4.LUT_INIT=16'b0010001011011101;
    LogicCell40 beamY_RNI93821_9_LC_1_8_4 (
            .in0(N__9296),
            .in1(N__7795),
            .in2(_gnd_net_),
            .in3(N__9608),
            .lcout(beamY_RNI93821Z0Z_9),
            .ltout(beamY_RNI93821Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM5433_0_8_LC_1_8_5.C_ON=1'b0;
    defparam beamY_RNIM5433_0_8_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIM5433_0_8_LC_1_8_5.LUT_INIT=16'b1010010101101001;
    LogicCell40 beamY_RNIM5433_0_8_LC_1_8_5 (
            .in0(N__12234),
            .in1(N__9297),
            .in2(N__7166),
            .in3(N__12058),
            .lcout(beamY_RNIM5433_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIR4K3_0_7_LC_1_8_6.C_ON=1'b0;
    defparam beamY_RNIIR4K3_0_7_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIIR4K3_0_7_LC_1_8_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 beamY_RNIIR4K3_0_7_LC_1_8_6 (
            .in0(N__8339),
            .in1(N__7286),
            .in2(_gnd_net_),
            .in3(N__8307),
            .lcout(beamY_RNIIR4K3_0Z0Z_7),
            .ltout(beamY_RNIIR4K3_0Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKM9GC_0_9_LC_1_8_7.C_ON=1'b0;
    defparam beamY_RNIKM9GC_0_9_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIKM9GC_0_9_LC_1_8_7.LUT_INIT=16'b0111010000110000;
    LogicCell40 beamY_RNIKM9GC_0_9_LC_1_8_7 (
            .in0(N__12235),
            .in1(N__7268),
            .in2(N__7151),
            .in3(N__7311),
            .lcout(beamY_RNIKM9GC_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DSP2_8_LC_1_9_0.C_ON=1'b0;
    defparam beamY_RNI9DSP2_8_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DSP2_8_LC_1_9_0.LUT_INIT=16'b1110000110110100;
    LogicCell40 beamY_RNI9DSP2_8_LC_1_9_0 (
            .in0(N__12061),
            .in1(N__8311),
            .in2(N__7279),
            .in3(N__9344),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axbxc5_2),
            .ltout(chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI41384_7_LC_1_9_1.C_ON=1'b0;
    defparam beamY_RNI41384_7_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI41384_7_LC_1_9_1.LUT_INIT=16'b1111000001101001;
    LogicCell40 beamY_RNI41384_7_LC_1_9_1 (
            .in0(N__9482),
            .in1(N__8652),
            .in2(N__7142),
            .in3(N__12062),
            .lcout(),
            .ltout(beamY_RNI41384Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBDEO7_7_LC_1_9_2.C_ON=1'b0;
    defparam beamY_RNIBDEO7_7_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIBDEO7_7_LC_1_9_2.LUT_INIT=16'b1110001011100010;
    LogicCell40 beamY_RNIBDEO7_7_LC_1_9_2 (
            .in0(N__7139),
            .in1(N__12169),
            .in2(N__7130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIH5LL11_5_LC_1_9_3.C_ON=1'b0;
    defparam beamY_RNIH5LL11_5_LC_1_9_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIH5LL11_5_LC_1_9_3.LUT_INIT=16'b0100100010000100;
    LogicCell40 beamY_RNIH5LL11_5_LC_1_9_3 (
            .in0(N__8464),
            .in1(N__9105),
            .in2(N__7127),
            .in3(N__7189),
            .lcout(chary_if_generate_plus_mult1_un54_sum_ac0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIIGUB_4_LC_1_9_4.C_ON=1'b0;
    defparam beamY_fast_RNIIGUB_4_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIIGUB_4_LC_1_9_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 beamY_fast_RNIIGUB_4_LC_1_9_4 (
            .in0(N__7903),
            .in1(N__7860),
            .in2(_gnd_net_),
            .in3(N__7834),
            .lcout(un8_beamylt9_0),
            .ltout(un8_beamylt9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI0A6L_7_LC_1_9_5.C_ON=1'b0;
    defparam beamY_fast_RNI0A6L_7_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI0A6L_7_LC_1_9_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_fast_RNI0A6L_7_LC_1_9_5 (
            .in0(N__9672),
            .in1(N__7952),
            .in2(N__7124),
            .in3(N__7938),
            .lcout(un5_visibley_c6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIQEC2_9_LC_1_9_6.C_ON=1'b0;
    defparam beamY_RNIIQEC2_9_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIIQEC2_9_LC_1_9_6.LUT_INIT=16'b1000100011101110;
    LogicCell40 beamY_RNIIQEC2_9_LC_1_9_6 (
            .in0(N__7274),
            .in1(N__8463),
            .in2(_gnd_net_),
            .in3(N__12244),
            .lcout(chary_if_generate_plus_mult1_un47_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP8FF1_1_7_LC_1_9_7.C_ON=1'b0;
    defparam beamY_RNIP8FF1_1_7_LC_1_9_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIP8FF1_1_7_LC_1_9_7.LUT_INIT=16'b1001100101101001;
    LogicCell40 beamY_RNIP8FF1_1_7_LC_1_9_7 (
            .in0(N__9481),
            .in1(N__8651),
            .in2(N__9353),
            .in3(N__12060),
            .lcout(beamY_RNIP8FF1_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUFT79_9_LC_1_10_0.C_ON=1'b0;
    defparam beamY_RNIUFT79_9_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIUFT79_9_LC_1_10_0.LUT_INIT=16'b0110110000110110;
    LogicCell40 beamY_RNIUFT79_9_LC_1_10_0 (
            .in0(N__7280),
            .in1(N__7330),
            .in2(N__8488),
            .in3(N__12254),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb4_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2BHS32_9_LC_1_10_1.C_ON=1'b0;
    defparam beamY_RNI2BHS32_9_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI2BHS32_9_LC_1_10_1.LUT_INIT=16'b1001011000101101;
    LogicCell40 beamY_RNI2BHS32_9_LC_1_10_1 (
            .in0(N__8481),
            .in1(N__7392),
            .in2(N__7775),
            .in3(N__7175),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBV5E51_0_8_LC_1_10_2.C_ON=1'b0;
    defparam beamY_RNIBV5E51_0_8_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIBV5E51_0_8_LC_1_10_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIBV5E51_0_8_LC_1_10_2 (
            .in0(N__7224),
            .in1(N__7326),
            .in2(N__7368),
            .in3(N__7203),
            .lcout(beamY_RNIBV5E51_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBV5E51_8_LC_1_10_3.C_ON=1'b0;
    defparam beamY_RNIBV5E51_8_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIBV5E51_8_LC_1_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIBV5E51_8_LC_1_10_3 (
            .in0(N__7204),
            .in1(N__7360),
            .in2(N__7334),
            .in3(N__7225),
            .lcout(),
            .ltout(beamY_RNIBV5E51Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8QGGE2_8_LC_1_10_4.C_ON=1'b0;
    defparam beamY_RNI8QGGE2_8_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI8QGGE2_8_LC_1_10_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNI8QGGE2_8_LC_1_10_4 (
            .in0(_gnd_net_),
            .in1(N__8270),
            .in2(N__7235),
            .in3(N__7232),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRV5601_8_LC_1_10_5.C_ON=1'b0;
    defparam beamY_RNIRV5601_8_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIRV5601_8_LC_1_10_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIRV5601_8_LC_1_10_5 (
            .in0(N__8269),
            .in1(N__8479),
            .in2(N__7205),
            .in3(N__7226),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVADQV_8_LC_1_10_6.C_ON=1'b0;
    defparam beamY_RNIVADQV_8_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIVADQV_8_LC_1_10_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNIVADQV_8_LC_1_10_6 (
            .in0(N__8263),
            .in1(N__7223),
            .in2(_gnd_net_),
            .in3(N__7199),
            .lcout(beamY_RNIVADQVZ0Z_8),
            .ltout(beamY_RNIVADQVZ0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2BHS32_0_9_LC_1_10_7.C_ON=1'b0;
    defparam beamY_RNI2BHS32_0_9_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI2BHS32_0_9_LC_1_10_7.LUT_INIT=16'b0110111100100110;
    LogicCell40 beamY_RNI2BHS32_0_9_LC_1_10_7 (
            .in0(N__7771),
            .in1(N__8480),
            .in2(N__7178),
            .in3(N__7174),
            .lcout(chary_if_generate_plus_mult1_un54_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV5SUC3_0_9_LC_1_11_0.C_ON=1'b0;
    defparam beamY_RNIV5SUC3_0_9_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIV5SUC3_0_9_LC_1_11_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIV5SUC3_0_9_LC_1_11_0 (
            .in0(N__7332),
            .in1(N__7367),
            .in2(N__8571),
            .in3(N__7394),
            .lcout(),
            .ltout(beamY_RNIV5SUC3_0Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0N9QT8_9_LC_1_11_1.C_ON=1'b0;
    defparam beamY_RNI0N9QT8_9_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI0N9QT8_9_LC_1_11_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNI0N9QT8_9_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(N__8740),
            .in2(N__7409),
            .in3(N__7295),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI3SC791_5_LC_1_11_3.C_ON=1'b0;
    defparam beamY_RNI3SC791_5_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI3SC791_5_LC_1_11_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNI3SC791_5_LC_1_11_3 (
            .in0(N__9110),
            .in1(N__7390),
            .in2(N__7369),
            .in3(N__7331),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIURID92_5_LC_1_11_4.C_ON=1'b0;
    defparam beamY_RNIURID92_5_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIURID92_5_LC_1_11_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIURID92_5_LC_1_11_4 (
            .in0(N__7391),
            .in1(N__9111),
            .in2(N__7406),
            .in3(N__8786),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb4_0),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEIALM5_4_LC_1_11_5.C_ON=1'b0;
    defparam beamY_RNIEIALM5_4_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIEIALM5_4_LC_1_11_5.LUT_INIT=16'b0010000000001000;
    LogicCell40 beamY_RNIEIALM5_4_LC_1_11_5 (
            .in0(N__10243),
            .in1(N__7503),
            .in2(N__7397),
            .in3(N__8556),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_7_d),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_13_LC_1_11_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_13_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_13_LC_1_11_6.LUT_INIT=16'b0000100111110000;
    LogicCell40 un114_pixel_6_1_5__g0_13_LC_1_11_6 (
            .in0(N__8557),
            .in1(N__8609),
            .in2(N__8807),
            .in3(N__9112),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV5SUC3_9_LC_1_11_7.C_ON=1'b0;
    defparam beamY_RNIV5SUC3_9_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIV5SUC3_9_LC_1_11_7.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIV5SUC3_9_LC_1_11_7 (
            .in0(N__7393),
            .in1(N__8552),
            .in2(N__7370),
            .in3(N__7333),
            .lcout(beamY_RNIV5SUC3Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIB6AOI5_5_LC_1_12_0.C_ON=1'b0;
    defparam beamY_RNIB6AOI5_5_LC_1_12_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIB6AOI5_5_LC_1_12_0.LUT_INIT=16'b0010110000011100;
    LogicCell40 beamY_RNIB6AOI5_5_LC_1_12_0 (
            .in0(N__8614),
            .in1(N__8806),
            .in2(N__9122),
            .in3(N__8579),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0),
            .ltout(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0797K_4_LC_1_12_1.C_ON=1'b0;
    defparam beamY_RNIJ0797K_4_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0797K_4_LC_1_12_1.LUT_INIT=16'b0011011011001001;
    LogicCell40 beamY_RNIJ0797K_4_LC_1_12_1 (
            .in0(N__8521),
            .in1(N__9984),
            .in2(N__7289),
            .in3(N__9852),
            .lcout(beamY_RNIJ0797KZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g1_0_0_LC_1_12_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g1_0_0_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g1_0_0_LC_1_12_2.LUT_INIT=16'b0110011001101001;
    LogicCell40 un114_pixel_6_1_5__g1_0_0_LC_1_12_2 (
            .in0(N__9988),
            .in1(N__10260),
            .in2(N__7463),
            .in3(N__8524),
            .lcout(g1_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g1_1_0_LC_1_12_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g1_1_0_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g1_1_0_LC_1_12_3.LUT_INIT=16'b0110011010011001;
    LogicCell40 un114_pixel_6_1_5__g1_1_0_LC_1_12_3 (
            .in0(N__10259),
            .in1(N__10321),
            .in2(_gnd_net_),
            .in3(N__9987),
            .lcout(g1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGMN7D3_4_LC_1_12_4.C_ON=1'b0;
    defparam beamY_RNIGMN7D3_4_LC_1_12_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIGMN7D3_4_LC_1_12_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNIGMN7D3_4_LC_1_12_4 (
            .in0(N__10253),
            .in1(N__7504),
            .in2(_gnd_net_),
            .in3(N__8580),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axb4_0),
            .ltout(chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI96MFKN_4_LC_1_12_5.C_ON=1'b0;
    defparam beamY_RNI96MFKN_4_LC_1_12_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI96MFKN_4_LC_1_12_5.LUT_INIT=16'b1110000100011110;
    LogicCell40 beamY_RNI96MFKN_4_LC_1_12_5 (
            .in0(N__8522),
            .in1(N__7441),
            .in2(N__7454),
            .in3(N__9985),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axb4_i),
            .ltout(chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g2_1_LC_1_12_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g2_1_LC_1_12_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g2_1_LC_1_12_6.LUT_INIT=16'b0000011000000000;
    LogicCell40 un114_pixel_6_1_5__g2_1_LC_1_12_6 (
            .in0(N__11377),
            .in1(N__11827),
            .in2(N__7451),
            .in3(N__7448),
            .lcout(g2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_4_LC_1_12_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_4_LC_1_12_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_4_LC_1_12_7.LUT_INIT=16'b1110000100011110;
    LogicCell40 un114_pixel_6_1_5__g0_4_LC_1_12_7 (
            .in0(N__8523),
            .in1(N__7442),
            .in2(N__7433),
            .in3(N__9986),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axb4_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g2_0_LC_1_13_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g2_0_LC_1_13_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g2_0_LC_1_13_0.LUT_INIT=16'b0001001000000000;
    LogicCell40 un114_pixel_6_1_5__g2_0_LC_1_13_0 (
            .in0(N__11376),
            .in1(N__7424),
            .in2(N__11831),
            .in3(N__7418),
            .lcout(),
            .ltout(g2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_7_LC_1_13_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_7_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_7_LC_1_13_1.LUT_INIT=16'b1100100100110110;
    LogicCell40 un114_pixel_6_1_5__g0_7_LC_1_13_1 (
            .in0(N__8729),
            .in1(N__7529),
            .in2(N__7412),
            .in3(N__10322),
            .lcout(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI074AD4_5_LC_1_13_3.C_ON=1'b0;
    defparam beamY_RNI074AD4_5_LC_1_13_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI074AD4_5_LC_1_13_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNI074AD4_5_LC_1_13_3 (
            .in0(_gnd_net_),
            .in1(N__7522),
            .in2(_gnd_net_),
            .in3(N__8578),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb4_i),
            .ltout(chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_2_0_LC_1_13_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_2_0_LC_1_13_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_2_0_LC_1_13_4.LUT_INIT=16'b0110100110010110;
    LogicCell40 un114_pixel_6_1_5__g0_2_0_LC_1_13_4 (
            .in0(N__11823),
            .in1(N__8695),
            .in2(N__7532),
            .in3(N__10016),
            .lcout(un114_pixel_6_1_5__g0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRLTLI4_0_5_LC_1_13_5.C_ON=1'b0;
    defparam beamY_RNIRLTLI4_0_5_LC_1_13_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIRLTLI4_0_5_LC_1_13_5.LUT_INIT=16'b0111000111010100;
    LogicCell40 beamY_RNIRLTLI4_0_5_LC_1_13_5 (
            .in0(N__9120),
            .in1(N__8613),
            .in2(N__10261),
            .in3(N__8577),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c4),
            .ltout(chary_if_generate_plus_mult1_un61_sum_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISDTA58_5_LC_1_13_6.C_ON=1'b0;
    defparam beamY_RNISDTA58_5_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam beamY_RNISDTA58_5_LC_1_13_6.LUT_INIT=16'b0101101010100101;
    LogicCell40 beamY_RNISDTA58_5_LC_1_13_6 (
            .in0(N__7523),
            .in1(_gnd_net_),
            .in2(N__7511),
            .in3(N__7508),
            .lcout(),
            .ltout(beamY_RNISDTA58Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0DLMCS_3_LC_1_13_7.C_ON=1'b0;
    defparam beamY_RNI0DLMCS_3_LC_1_13_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI0DLMCS_3_LC_1_13_7.LUT_INIT=16'b0001000110101111;
    LogicCell40 beamY_RNI0DLMCS_3_LC_1_13_7 (
            .in0(N__11822),
            .in1(N__11375),
            .in2(N__7487),
            .in3(N__7484),
            .lcout(chary_if_generate_plus_mult1_un75_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_2_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_2_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_2_0 (
            .in0(_gnd_net_),
            .in1(N__7592),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVL21_LC_2_2_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVL21_LC_2_2_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVL21_LC_2_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVL21_LC_2_2_1 (
            .in0(_gnd_net_),
            .in1(N__7469),
            .in2(N__14251),
            .in3(N__7478),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1N21_LC_2_2_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1N21_LC_2_2_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1N21_LC_2_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1N21_LC_2_2_2 (
            .in0(_gnd_net_),
            .in1(N__12102),
            .in2(N__14252),
            .in3(N__7475),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_2_2_3.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_2_2_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_2_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_2_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7472),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2B511_0_9_LC_2_2_6.C_ON=1'b0;
    defparam beamY_RNI2B511_0_9_LC_2_2_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI2B511_0_9_LC_2_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNI2B511_0_9_LC_2_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12101),
            .lcout(beamY_RNI2B511_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_3_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_3_0 (
            .in0(_gnd_net_),
            .in1(N__12255),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6U_LC_2_3_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6U_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6U_LC_2_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6U_LC_2_3_1 (
            .in0(_gnd_net_),
            .in1(N__7583),
            .in2(N__14275),
            .in3(N__7577),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEA1_LC_2_3_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEA1_LC_2_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEA1_LC_2_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEA1_LC_2_3_2 (
            .in0(_gnd_net_),
            .in1(N__7574),
            .in2(N__14277),
            .in3(N__7568),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HA1_LC_2_3_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HA1_LC_2_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HA1_LC_2_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HA1_LC_2_3_3 (
            .in0(_gnd_net_),
            .in1(N__7565),
            .in2(N__14276),
            .in3(N__7559),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_2_3_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_2_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_2_3_4 (
            .in0(_gnd_net_),
            .in1(N__7677),
            .in2(_gnd_net_),
            .in3(N__7556),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_2_3_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_2_3_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_2_3_5 (
            .in0(N__7550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7553),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_2_3_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_2_3_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_2_3_6.LUT_INIT=16'b0011001100110011;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_2_3_6 (
            .in0(_gnd_net_),
            .in1(N__7549),
            .in2(_gnd_net_),
            .in3(N__7678),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0 (
            .in0(_gnd_net_),
            .in1(N__8482),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_2_4_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_2_4_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_2_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_2_4_1 (
            .in0(_gnd_net_),
            .in1(N__7784),
            .in2(N__7651),
            .in3(N__7535),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVH1_LC_2_4_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVH1_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVH1_LC_2_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVH1_LC_2_4_2 (
            .in0(_gnd_net_),
            .in1(N__7646),
            .in2(N__7736),
            .in3(N__7718),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8U1_LC_2_4_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8U1_LC_2_4_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8U1_LC_2_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8U1_LC_2_4_3 (
            .in0(_gnd_net_),
            .in1(N__7715),
            .in2(N__7652),
            .in3(N__7700),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINI2Q2_LC_2_4_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINI2Q2_LC_2_4_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINI2Q2_LC_2_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINI2Q2_LC_2_4_4 (
            .in0(N__7616),
            .in1(N__7628),
            .in2(N__7697),
            .in3(N__7682),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_2_4_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_2_4_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_2_4_5 (
            .in0(N__7650),
            .in1(N__7679),
            .in2(N__7664),
            .in3(N__7655),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_2_4_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_2_4_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_2_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_2_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7642),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_2_4_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_2_4_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_2_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_2_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7615),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx_LC_2_5_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx_LC_2_5_0.LUT_INIT=16'b1100110000110011;
    LogicCell40 row_1_if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx_LC_2_5_0 (
            .in0(_gnd_net_),
            .in1(N__9260),
            .in2(_gnd_net_),
            .in3(N__8318),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_5_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_5_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_5_4.LUT_INIT=16'b0100001010010100;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_5_4 (
            .in0(N__12257),
            .in1(N__12154),
            .in2(N__8489),
            .in3(N__12082),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12256),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIM5M02_9_LC_2_6_0.C_ON=1'b0;
    defparam beamY_RNIM5M02_9_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIM5M02_9_LC_2_6_0.LUT_INIT=16'b0101100110100110;
    LogicCell40 beamY_RNIM5M02_9_LC_2_6_0 (
            .in0(N__12259),
            .in1(N__9328),
            .in2(N__7802),
            .in3(N__9588),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_8_LC_2_6_1.C_ON=1'b0;
    defparam beamY_8_LC_2_6_1.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_2_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_8_LC_2_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8141),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13139),
            .ce(N__11545),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_6_LC_2_6_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_6_LC_2_6_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_6_LC_2_6_5.LUT_INIT=16'b0000000011100111;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_6_LC_2_6_5 (
            .in0(N__12084),
            .in1(N__12260),
            .in2(N__12173),
            .in3(N__8475),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_6_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_6_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_6_6.LUT_INIT=16'b0010010001001001;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_6_6 (
            .in0(N__12258),
            .in1(N__12158),
            .in2(N__8487),
            .in3(N__12083),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIF0BK31_LC_2_7_0.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIF0BK31_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIF0BK31_LC_2_7_0.LUT_INIT=16'b1111111110111011;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIF0BK31_LC_2_7_0 (
            .in0(N__7757),
            .in1(N__10947),
            .in2(_gnd_net_),
            .in3(N__7748),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_7_1.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_7_1 (
            .in0(N__10948),
            .in1(N__14278),
            .in2(_gnd_net_),
            .in3(N__11321),
            .lcout(beamY_i_2),
            .ltout(beamY_i_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_1_LC_2_7_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_1_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_1_LC_2_7_2.LUT_INIT=16'b0001100010001000;
    LogicCell40 un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_1_LC_2_7_2 (
            .in0(N__7756),
            .in1(N__7747),
            .in2(N__7739),
            .in3(N__10903),
            .lcout(un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_3_LC_2_7_6.C_ON=1'b0;
    defparam beamY_3_LC_2_7_6.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_2_7_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_3_LC_2_7_6 (
            .in0(_gnd_net_),
            .in1(N__8051),
            .in2(_gnd_net_),
            .in3(N__11446),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13138),
            .ce(N__11530),
            .sr(_gnd_net_));
    defparam beamY_fast_3_LC_2_8_0.C_ON=1'b0;
    defparam beamY_fast_3_LC_2_8_0.SEQ_MODE=4'b1000;
    defparam beamY_fast_3_LC_2_8_0.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_fast_3_LC_2_8_0 (
            .in0(N__8047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(beamY_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_fast_6_LC_2_8_1.C_ON=1'b0;
    defparam beamY_fast_6_LC_2_8_1.SEQ_MODE=4'b1000;
    defparam beamY_fast_6_LC_2_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_6_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7988),
            .lcout(beamY_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_fast_8_LC_2_8_2.C_ON=1'b0;
    defparam beamY_fast_8_LC_2_8_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_8_LC_2_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_8_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8137),
            .lcout(beamY_fastZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_7_LC_2_8_4.C_ON=1'b0;
    defparam beamY_7_LC_2_8_4.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_2_8_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_7_LC_2_8_4 (
            .in0(_gnd_net_),
            .in1(N__7966),
            .in2(_gnd_net_),
            .in3(N__11427),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_fast_7_LC_2_8_5.C_ON=1'b0;
    defparam beamY_fast_7_LC_2_8_5.SEQ_MODE=4'b1000;
    defparam beamY_fast_7_LC_2_8_5.LUT_INIT=16'b0101000001010000;
    LogicCell40 beamY_fast_7_LC_2_8_5 (
            .in0(N__11430),
            .in1(_gnd_net_),
            .in2(N__7970),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_fast_4_LC_2_8_6.C_ON=1'b0;
    defparam beamY_fast_4_LC_2_8_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_4_LC_2_8_6.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_fast_4_LC_2_8_6 (
            .in0(N__8027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11429),
            .lcout(beamY_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13136),
            .ce(N__11543),
            .sr(_gnd_net_));
    defparam beamY_RNID2EU_6_LC_2_9_0.C_ON=1'b0;
    defparam beamY_RNID2EU_6_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam beamY_RNID2EU_6_LC_2_9_0.LUT_INIT=16'b1010101010011001;
    LogicCell40 beamY_RNID2EU_6_LC_2_9_0 (
            .in0(N__9491),
            .in1(N__9411),
            .in2(_gnd_net_),
            .in3(N__7811),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIT5UF_4_LC_2_9_1.C_ON=1'b0;
    defparam beamY_fast_RNIT5UF_4_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIT5UF_4_LC_2_9_1.LUT_INIT=16'b0101010001000100;
    LogicCell40 beamY_fast_RNIT5UF_4_LC_2_9_1 (
            .in0(N__7939),
            .in1(N__7918),
            .in2(N__7904),
            .in3(N__7833),
            .lcout(),
            .ltout(beamY_fast_RNIT5UFZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIKRSR_5_LC_2_9_2.C_ON=1'b0;
    defparam beamY_fast_RNIKRSR_5_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIKRSR_5_LC_2_9_2.LUT_INIT=16'b1111000000100010;
    LogicCell40 beamY_fast_RNIKRSR_5_LC_2_9_2 (
            .in0(N__7919),
            .in1(N__7940),
            .in2(N__7814),
            .in3(N__7861),
            .lcout(un5_visibley_ac0_7),
            .ltout(un5_visibley_ac0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICOMV_6_LC_2_9_3.C_ON=1'b0;
    defparam beamY_RNICOMV_6_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam beamY_RNICOMV_6_LC_2_9_3.LUT_INIT=16'b0000000101010111;
    LogicCell40 beamY_RNICOMV_6_LC_2_9_3 (
            .in0(N__9607),
            .in1(N__9412),
            .in2(N__7805),
            .in3(N__9492),
            .lcout(chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_5_LC_2_9_4.C_ON=1'b0;
    defparam beamY_fast_5_LC_2_9_4.SEQ_MODE=4'b1000;
    defparam beamY_fast_5_LC_2_9_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_fast_5_LC_2_9_4 (
            .in0(N__8006),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13134),
            .ce(N__11555),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI6FUF_7_LC_2_9_5.C_ON=1'b0;
    defparam beamY_fast_RNI6FUF_7_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI6FUF_7_LC_2_9_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_fast_RNI6FUF_7_LC_2_9_5 (
            .in0(N__7951),
            .in1(N__7937),
            .in2(N__7886),
            .in3(N__7917),
            .lcout(),
            .ltout(un5_visibley_ac0_11_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2B511_9_LC_2_9_6.C_ON=1'b0;
    defparam beamY_RNI2B511_9_LC_2_9_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI2B511_9_LC_2_9_6.LUT_INIT=16'b1100110011000011;
    LogicCell40 beamY_RNI2B511_9_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(N__9606),
            .in2(N__7907),
            .in3(N__7871),
            .lcout(chary_if_generate_plus_mult1_un33_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIT5UF_8_LC_2_9_7.C_ON=1'b0;
    defparam beamY_fast_RNIT5UF_8_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIT5UF_8_LC_2_9_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_fast_RNIT5UF_8_LC_2_9_7 (
            .in0(N__7899),
            .in1(N__7859),
            .in2(N__7885),
            .in3(N__7832),
            .lcout(un5_visibley_c7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_2_10_1.C_ON=1'b0;
    defparam beamY_2_LC_2_10_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_2_10_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_2_LC_2_10_1 (
            .in0(N__8065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13135),
            .ce(N__11544),
            .sr(_gnd_net_));
    defparam beamY_4_LC_2_10_3.C_ON=1'b0;
    defparam beamY_4_LC_2_10_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_2_10_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_4_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(N__8026),
            .in2(_gnd_net_),
            .in3(N__11447),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13135),
            .ce(N__11544),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un8_beamylto4_0_LC_2_10_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un8_beamylto4_0_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un8_beamylto4_0_LC_2_10_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 un114_pixel_6_1_5__un8_beamylto4_0_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__7865),
            .in2(_gnd_net_),
            .in3(N__7835),
            .lcout(un5_visibley_c2),
            .ltout(un5_visibley_c2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISKOB_5_LC_2_10_5.C_ON=1'b0;
    defparam beamY_RNISKOB_5_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam beamY_RNISKOB_5_LC_2_10_5.LUT_INIT=16'b1111111111101100;
    LogicCell40 beamY_RNISKOB_5_LC_2_10_5 (
            .in0(N__9798),
            .in1(N__9409),
            .in2(N__7838),
            .in3(N__9670),
            .lcout(un5_visibley_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_2_LC_2_10_7.C_ON=1'b0;
    defparam beamY_fast_2_LC_2_10_7.SEQ_MODE=4'b1000;
    defparam beamY_fast_2_LC_2_10_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_fast_2_LC_2_10_7 (
            .in0(N__8066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13135),
            .ce(N__11544),
            .sr(_gnd_net_));
    defparam beamY_6_LC_2_11_3.C_ON=1'b0;
    defparam beamY_6_LC_2_11_3.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_2_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_6_LC_2_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7984),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13137),
            .ce(N__11554),
            .sr(_gnd_net_));
    defparam beamY_5_LC_2_11_4.C_ON=1'b0;
    defparam beamY_5_LC_2_11_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_2_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_5_LC_2_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8002),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13137),
            .ce(N__11554),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_2_12_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_2_12_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_2_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_2_12_0 (
            .in0(_gnd_net_),
            .in1(N__15132),
            .in2(N__14939),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_RNIAL73_LC_2_12_1.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_2_12_1.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_2_12_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_1_c_RNIAL73_LC_2_12_1 (
            .in0(_gnd_net_),
            .in1(N__11378),
            .in2(_gnd_net_),
            .in3(N__8054),
            .lcout(un21_beamy_cry_1_c_RNIALZ0Z73),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_2_c_RNICO83_LC_2_12_2.C_ON=1'b1;
    defparam un21_beamy_cry_2_c_RNICO83_LC_2_12_2.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_2_c_RNICO83_LC_2_12_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_2_c_RNICO83_LC_2_12_2 (
            .in0(_gnd_net_),
            .in1(N__11810),
            .in2(_gnd_net_),
            .in3(N__8030),
            .lcout(un21_beamy_cry_2_c_RNICOZ0Z83),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_3_c_RNIER93_LC_2_12_3.C_ON=1'b1;
    defparam un21_beamy_cry_3_c_RNIER93_LC_2_12_3.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_3_c_RNIER93_LC_2_12_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_3_c_RNIER93_LC_2_12_3 (
            .in0(_gnd_net_),
            .in1(N__9839),
            .in2(_gnd_net_),
            .in3(N__8009),
            .lcout(un21_beamy_cry_3_c_RNIERZ0Z93),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_2_12_4.C_ON=1'b1;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_2_12_4.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_2_12_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_4_c_RNIGUA3_LC_2_12_4 (
            .in0(_gnd_net_),
            .in1(N__9671),
            .in2(_gnd_net_),
            .in3(N__7991),
            .lcout(un21_beamy_cry_4_c_RNIGUAZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_5_c_RNII1C3_LC_2_12_5.C_ON=1'b1;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_2_12_5.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_2_12_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_5_c_RNII1C3_LC_2_12_5 (
            .in0(_gnd_net_),
            .in1(N__9410),
            .in2(_gnd_net_),
            .in3(N__7973),
            .lcout(un21_beamy_cry_5_c_RNII1CZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_2_12_6.C_ON=1'b1;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_2_12_6.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_2_12_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_6_c_RNIK4D3_LC_2_12_6 (
            .in0(_gnd_net_),
            .in1(N__9510),
            .in2(_gnd_net_),
            .in3(N__7955),
            .lcout(un21_beamy_cry_6_c_RNIK4DZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_2_12_7.C_ON=1'b1;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_2_12_7.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_2_12_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_7_c_RNIM7E3_LC_2_12_7 (
            .in0(_gnd_net_),
            .in1(N__9340),
            .in2(_gnd_net_),
            .in3(N__8120),
            .lcout(un21_beamy_cry_7_c_RNIM7EZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_9_LC_2_13_0.C_ON=1'b0;
    defparam beamY_9_LC_2_13_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_2_13_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_2_13_0 (
            .in0(N__9605),
            .in1(N__11453),
            .in2(_gnd_net_),
            .in3(N__8117),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13140),
            .ce(N__11546),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_5_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_5_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_5_3 (
            .in0(N__14238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9148),
            .lcout(if_generate_plus_mult1_un61_sum_axbxc5),
            .ltout(if_generate_plus_mult1_un61_sum_axbxc5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_5_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_5_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_5_4.LUT_INIT=16'b1000011001111001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_5_4 (
            .in0(N__9097),
            .in1(N__8110),
            .in2(N__8114),
            .in3(N__8234),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_0_LC_4_5_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_0_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_7_0_LC_4_5_6.LUT_INIT=16'b0111010110110010;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_7_0_LC_4_5_6 (
            .in0(N__9096),
            .in1(N__10372),
            .in2(N__8111),
            .in3(N__8233),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_5_LC_4_5_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_5_LC_4_5_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_ac0_5_LC_4_5_7.LUT_INIT=16'b0010100010000010;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_ac0_5_LC_4_5_7 (
            .in0(N__10241),
            .in1(N__9149),
            .in2(N__14271),
            .in3(N__9095),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_d_LC_4_6_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_d_LC_4_6_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_d_LC_4_6_0.LUT_INIT=16'b0100010000000000;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_7_d_LC_4_6_0 (
            .in0(N__8089),
            .in1(N__8235),
            .in2(_gnd_net_),
            .in3(N__9072),
            .lcout(),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_6_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_6_1.LUT_INIT=16'b1111001011110101;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_6_1 (
            .in0(N__8246),
            .in1(N__10396),
            .in2(N__8096),
            .in3(N__8471),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_c5),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m5_i_LC_4_6_2.C_ON=1'b0;
    defparam row_1_if_m5_i_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam row_1_if_m5_i_LC_4_6_2.LUT_INIT=16'b0101101010100101;
    LogicCell40 row_1_if_m5_i_LC_4_6_2 (
            .in0(N__14272),
            .in1(_gnd_net_),
            .in2(N__8093),
            .in3(N__9075),
            .lcout(row_1_if_N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_4_6_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_4_6_3.LUT_INIT=16'b1100100111000011;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_4_6_3 (
            .in0(N__9073),
            .in1(N__8090),
            .in2(N__8078),
            .in3(N__8237),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_1_LC_4_6_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_1_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_1_LC_4_6_4.LUT_INIT=16'b0110011011011101;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_1_LC_4_6_4 (
            .in0(N__12271),
            .in1(N__12174),
            .in2(_gnd_net_),
            .in3(N__12108),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_m5x_LC_4_6_5.C_ON=1'b0;
    defparam row_1_if_m5x_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam row_1_if_m5x_LC_4_6_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_m5x_LC_4_6_5 (
            .in0(N__9074),
            .in1(N__14273),
            .in2(N__10262),
            .in3(N__9150),
            .lcout(row_1_if_i4_mux_i),
            .ltout(row_1_if_i4_mux_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_1_LC_4_6_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_1_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_1_LC_4_6_6.LUT_INIT=16'b0010011010001001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_1_LC_4_6_6 (
            .in0(N__10242),
            .in1(N__8185),
            .in2(N__8240),
            .in3(N__8236),
            .lcout(),
            .ltout(row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_LC_4_6_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_LC_4_6_7.LUT_INIT=16'b0000110010101100;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_LC_4_6_7 (
            .in0(N__10094),
            .in1(N__8204),
            .in2(N__8198),
            .in3(N__8195),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_7_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_7_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_7_0 (
            .in0(N__10257),
            .in1(N__11008),
            .in2(N__10096),
            .in3(N__11049),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc3),
            .ltout(if_generate_plus_mult1_un75_sum_axbxc3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x0_LC_4_7_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x0_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x0_LC_4_7_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axb4_x0_LC_4_7_1 (
            .in0(N__11050),
            .in1(N__8163),
            .in2(N__8189),
            .in3(N__11009),
            .lcout(if_generate_plus_mult1_un82_sum_axb4_x0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_7_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_7_3.LUT_INIT=16'b0110011010011001;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_7_3 (
            .in0(N__14274),
            .in1(N__8186),
            .in2(_gnd_net_),
            .in3(N__9151),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1),
            .ltout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_7_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_7_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_7_4 (
            .in0(N__8164),
            .in1(N__8357),
            .in2(N__8171),
            .in3(N__11052),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x1_LC_4_7_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x1_LC_4_7_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_x1_LC_4_7_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axb4_x1_LC_4_7_5 (
            .in0(N__11051),
            .in1(N__11010),
            .in2(N__8168),
            .in3(N__8147),
            .lcout(),
            .ltout(if_generate_plus_mult1_un82_sum_axb4_x1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_ns_LC_4_7_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_ns_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_ns_LC_4_7_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axb4_ns_LC_4_7_6 (
            .in0(_gnd_net_),
            .in1(N__8356),
            .in2(N__8348),
            .in3(N__8345),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP8FF1_0_7_LC_4_8_1.C_ON=1'b0;
    defparam beamY_RNIP8FF1_0_7_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIP8FF1_0_7_LC_4_8_1.LUT_INIT=16'b1010010110010110;
    LogicCell40 beamY_RNIP8FF1_0_7_LC_4_8_1 (
            .in0(N__9499),
            .in1(N__9335),
            .in2(N__8673),
            .in3(N__12103),
            .lcout(beamY_RNIP8FF1_0Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un5_beamx_3_LC_4_8_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un5_beamx_3_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un5_beamx_3_LC_4_8_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 un114_pixel_6_1_5__un5_beamx_3_LC_4_8_3 (
            .in0(N__9846),
            .in1(N__15170),
            .in2(_gnd_net_),
            .in3(N__9336),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un5_beamx_5_LC_4_8_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un5_beamx_5_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un5_beamx_5_LC_4_8_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_6_1_5__un5_beamx_5_LC_4_8_4 (
            .in0(N__14921),
            .in1(N__9500),
            .in2(N__8327),
            .in3(N__9625),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un5_beamx_LC_4_8_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un5_beamx_LC_4_8_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un5_beamx_LC_4_8_5.LUT_INIT=16'b0000000010000000;
    LogicCell40 un114_pixel_6_1_5__un5_beamx_LC_4_8_5 (
            .in0(N__9176),
            .in1(N__11772),
            .in2(N__8324),
            .in3(N__11329),
            .lcout(un5_beamx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_5_LC_4_8_6.C_ON=1'b0;
    defparam beamY_RNI6125_5_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_5_LC_4_8_6.LUT_INIT=16'b1000000001111111;
    LogicCell40 beamY_RNI6125_5_LC_4_8_6 (
            .in0(N__11328),
            .in1(N__9845),
            .in2(N__11809),
            .in3(N__9691),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_4_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_4_8_7.LUT_INIT=16'b0100110110011011;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_4_8_7 (
            .in0(N__12270),
            .in1(N__12176),
            .in2(N__8486),
            .in3(N__12104),
            .lcout(if_generate_plus_mult1_un54_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP8FF1_7_LC_4_9_0.C_ON=1'b0;
    defparam beamY_RNIP8FF1_7_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIP8FF1_7_LC_4_9_0.LUT_INIT=16'b1100110011101101;
    LogicCell40 beamY_RNIP8FF1_7_LC_4_9_0 (
            .in0(N__9522),
            .in1(N__9346),
            .in2(N__8675),
            .in3(N__12091),
            .lcout(),
            .ltout(beamY_RNIP8FF1Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIR4K3_7_LC_4_9_1.C_ON=1'b0;
    defparam beamY_RNIIR4K3_7_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIIR4K3_7_LC_4_9_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 beamY_RNIIR4K3_7_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(N__8630),
            .in2(N__8321),
            .in3(N__8317),
            .lcout(chary_if_generate_plus_mult1_un40_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP8FF1_2_7_LC_4_9_2.C_ON=1'b0;
    defparam beamY_RNIP8FF1_2_7_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIP8FF1_2_7_LC_4_9_2.LUT_INIT=16'b0011001110110111;
    LogicCell40 beamY_RNIP8FF1_2_7_LC_4_9_2 (
            .in0(N__9521),
            .in1(N__9345),
            .in2(N__8674),
            .in3(N__12090),
            .lcout(beamY_RNIP8FF1_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_4_9_4.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_4_9_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_4_9_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIHUG2_0_3_LC_4_9_4 (
            .in0(_gnd_net_),
            .in1(N__11781),
            .in2(_gnd_net_),
            .in3(N__11366),
            .lcout(),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_beamylto6_LC_4_9_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_beamylto6_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_beamylto6_LC_4_9_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 un114_pixel_6_1_5__un4_beamylto6_LC_4_9_5 (
            .in0(N__9847),
            .in1(N__9426),
            .in2(N__8624),
            .in3(N__9692),
            .lcout(un4_beamylt8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un8_beamylto9_0_LC_4_10_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un8_beamylto9_0_LC_4_10_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un8_beamylto9_0_LC_4_10_4.LUT_INIT=16'b0000000000010001;
    LogicCell40 un114_pixel_6_1_5__un8_beamylto9_0_LC_4_10_4 (
            .in0(N__9350),
            .in1(N__9523),
            .in2(_gnd_net_),
            .in3(N__9609),
            .lcout(un114_pixel_6_1_5__un8_beamylto9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRLTLI4_5_LC_4_11_1.C_ON=1'b0;
    defparam beamY_RNIRLTLI4_5_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIRLTLI4_5_LC_4_11_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIRLTLI4_5_LC_4_11_1 (
            .in0(N__8621),
            .in1(N__9109),
            .in2(N__10249),
            .in3(N__8582),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIB6AOI5_0_5_LC_4_11_5.C_ON=1'b0;
    defparam beamY_RNIB6AOI5_0_5_LC_4_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIB6AOI5_0_5_LC_4_11_5.LUT_INIT=16'b0010110000011100;
    LogicCell40 beamY_RNIB6AOI5_0_5_LC_4_11_5 (
            .in0(N__8620),
            .in1(N__8808),
            .in2(N__9121),
            .in3(N__8581),
            .lcout(),
            .ltout(beamY_RNIB6AOI5_0Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPOKD9B_5_LC_4_11_6.C_ON=1'b0;
    defparam beamY_RNIPOKD9B_5_LC_4_11_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIPOKD9B_5_LC_4_11_6.LUT_INIT=16'b1111111111110000;
    LogicCell40 beamY_RNIPOKD9B_5_LC_4_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8528),
            .in3(N__8525),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISKOB_0_5_LC_4_11_7.C_ON=1'b0;
    defparam beamY_RNISKOB_0_5_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam beamY_RNISKOB_0_5_LC_4_11_7.LUT_INIT=16'b1100110010010011;
    LogicCell40 beamY_RNISKOB_0_5_LC_4_11_7 (
            .in0(N__8501),
            .in1(N__9413),
            .in2(N__9853),
            .in3(N__9673),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI3GESM7_4_LC_4_12_2.C_ON=1'b0;
    defparam beamY_RNI3GESM7_4_LC_4_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI3GESM7_4_LC_4_12_2.LUT_INIT=16'b1000101000101010;
    LogicCell40 beamY_RNI3GESM7_4_LC_4_12_2 (
            .in0(N__8764),
            .in1(N__8809),
            .in2(N__10238),
            .in3(N__8752),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c5_0),
            .ltout(chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_11_LC_4_12_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_11_LC_4_12_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_11_LC_4_12_3.LUT_INIT=16'b1100100100110110;
    LogicCell40 un114_pixel_6_1_5__g0_11_LC_4_12_3 (
            .in0(N__8825),
            .in1(N__11815),
            .in2(N__8816),
            .in3(N__11593),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_5_LC_4_12_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_5_LC_4_12_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_5_LC_4_12_4.LUT_INIT=16'b0110110110111100;
    LogicCell40 un114_pixel_6_1_5__g0_0_5_LC_4_12_4 (
            .in0(N__8714),
            .in1(N__14920),
            .in2(N__8813),
            .in3(N__11367),
            .lcout(un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILT8E7K_3_LC_4_12_6.C_ON=1'b0;
    defparam beamY_RNILT8E7K_3_LC_4_12_6.SEQ_MODE=4'b0000;
    defparam beamY_RNILT8E7K_3_LC_4_12_6.LUT_INIT=16'b0111000111010100;
    LogicCell40 beamY_RNILT8E7K_3_LC_4_12_6 (
            .in0(N__10198),
            .in1(N__10301),
            .in2(N__10105),
            .in3(N__10020),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI3GESM7_0_4_LC_4_12_7.C_ON=1'b0;
    defparam beamY_RNI3GESM7_0_4_LC_4_12_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI3GESM7_0_4_LC_4_12_7.LUT_INIT=16'b1000110001001100;
    LogicCell40 beamY_RNI3GESM7_0_4_LC_4_12_7 (
            .in0(N__8810),
            .in1(N__8765),
            .in2(N__10258),
            .in3(N__8753),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c5_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_17_1_LC_4_13_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_17_1_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_17_1_LC_4_13_0.LUT_INIT=16'b0101010111101010;
    LogicCell40 un114_pixel_6_1_5__g0_17_1_LC_4_13_0 (
            .in0(N__10853),
            .in1(N__8681),
            .in2(N__10106),
            .in3(N__11677),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g0_17Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_17_LC_4_13_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_17_LC_4_13_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_17_LC_4_13_1.LUT_INIT=16'b0110100110010110;
    LogicCell40 un114_pixel_6_1_5__g0_17_LC_4_13_1 (
            .in0(N__9717),
            .in1(N__11592),
            .in2(N__8717),
            .in3(N__9746),
            .lcout(chary_if_generate_plus_mult1_un75_sum_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKC087T_5_LC_4_13_3.C_ON=1'b0;
    defparam beamY_RNIKC087T_5_LC_4_13_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIKC087T_5_LC_4_13_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIKC087T_5_LC_4_13_3 (
            .in0(N__8708),
            .in1(N__10310),
            .in2(N__8699),
            .in3(N__10021),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axbxc5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4VNB7K_0_4_LC_4_13_4.C_ON=1'b0;
    defparam beamY_RNI4VNB7K_0_4_LC_4_13_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI4VNB7K_0_4_LC_4_13_4.LUT_INIT=16'b0101101010100101;
    LogicCell40 beamY_RNI4VNB7K_0_4_LC_4_13_4 (
            .in0(N__10022),
            .in1(_gnd_net_),
            .in2(N__10320),
            .in3(N__10237),
            .lcout(g1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0 (
            .in0(_gnd_net_),
            .in1(N__15279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_5_4_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_5_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_5_4_1 (
            .in0(_gnd_net_),
            .in1(N__8860),
            .in2(N__10352),
            .in3(N__8873),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_5_4_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_5_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_5_4_2 (
            .in0(_gnd_net_),
            .in1(N__9929),
            .in2(N__9896),
            .in3(N__8870),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_5_4_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_5_4_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_5_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_5_4_3 (
            .in0(N__8923),
            .in1(N__8861),
            .in2(N__9920),
            .in3(N__8867),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_5_4_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_5_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__9908),
            .in2(_gnd_net_),
            .in3(N__8864),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_5_4_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_5_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_5_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9891),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_5_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_5_0 (
            .in0(_gnd_net_),
            .in1(N__16131),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_5_5_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_5_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_5_5_1 (
            .in0(_gnd_net_),
            .in1(N__8903),
            .in2(N__8897),
            .in3(N__8852),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_5_5_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_5_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_5_5_2 (
            .in0(_gnd_net_),
            .in1(N__8849),
            .in2(N__8924),
            .in3(N__8843),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_5_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_5_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_5_3 (
            .in0(_gnd_net_),
            .in1(N__8831),
            .in2(N__8840),
            .in3(N__8919),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_5_5_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_5_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_5_5_4 (
            .in0(_gnd_net_),
            .in1(N__8933),
            .in2(_gnd_net_),
            .in3(N__8927),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_5_5_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_5_5_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_5_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8918),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_5_6.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_5_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_5_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15280),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_5_6_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_5_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_5_6_0 (
            .in0(_gnd_net_),
            .in1(N__10487),
            .in2(N__14497),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_5_6_1.C_ON=1'b1;
    defparam beamX_2_LC_5_6_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_5_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_5_6_1 (
            .in0(_gnd_net_),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__8888),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_5_6_2.C_ON=1'b1;
    defparam beamX_3_LC_5_6_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_5_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_5_6_2 (
            .in0(_gnd_net_),
            .in1(N__10736),
            .in2(_gnd_net_),
            .in3(N__8885),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_5_6_3.C_ON=1'b1;
    defparam beamX_4_LC_5_6_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_5_6_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_5_6_3 (
            .in0(N__11509),
            .in1(N__10772),
            .in2(_gnd_net_),
            .in3(N__8882),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_5_6_4.C_ON=1'b1;
    defparam beamX_5_LC_5_6_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_5_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_5_6_4 (
            .in0(_gnd_net_),
            .in1(N__10686),
            .in2(_gnd_net_),
            .in3(N__8879),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_5_6_5.C_ON=1'b1;
    defparam beamX_6_LC_5_6_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_5_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_5_6_5 (
            .in0(_gnd_net_),
            .in1(N__10564),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_5_6_6.C_ON=1'b1;
    defparam beamX_7_LC_5_6_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_5_6_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_5_6_6 (
            .in0(_gnd_net_),
            .in1(N__11171),
            .in2(_gnd_net_),
            .in3(N__8972),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_5_6_7.C_ON=1'b1;
    defparam beamX_8_LC_5_6_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_5_6_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_5_6_7 (
            .in0(_gnd_net_),
            .in1(N__10634),
            .in2(_gnd_net_),
            .in3(N__8969),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__13145),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_5_7_0.C_ON=1'b1;
    defparam beamX_9_LC_5_7_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_5_7_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(N__8966),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__13142),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_5_7_1.C_ON=1'b0;
    defparam beamX_10_LC_5_7_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_5_7_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_5_7_1 (
            .in0(N__11138),
            .in1(N__11508),
            .in2(_gnd_net_),
            .in3(N__8963),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13142),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_1_LC_5_7_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_1_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_1_LC_5_7_3.LUT_INIT=16'b0000010101000101;
    LogicCell40 un114_pixel_6_1_5__un4_row_1_LC_5_7_3 (
            .in0(N__8960),
            .in1(N__11808),
            .in2(N__10095),
            .in3(N__11365),
            .lcout(un114_pixel_6_1_5__un4_rowZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un3_beamx_LC_5_7_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un3_beamx_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un3_beamx_LC_5_7_7.LUT_INIT=16'b0000001000000000;
    LogicCell40 un114_pixel_6_1_5__un3_beamx_LC_5_7_7 (
            .in0(N__11190),
            .in1(N__11170),
            .in2(N__10690),
            .in3(N__10358),
            .lcout(un3_beamx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un15_beamy_0_LC_5_8_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un15_beamy_0_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un15_beamy_0_LC_5_8_1.LUT_INIT=16'b0000110100001111;
    LogicCell40 un114_pixel_6_1_5__un15_beamy_0_LC_5_8_1 (
            .in0(N__8954),
            .in1(N__8945),
            .in2(N__11139),
            .in3(N__9174),
            .lcout(un114_pixel_6_1_5__un15_beamyZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un1_beamxlto6_LC_5_8_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un1_beamxlto6_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un1_beamxlto6_LC_5_8_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_6_1_5__un1_beamxlto6_LC_5_8_3 (
            .in0(N__10739),
            .in1(N__10694),
            .in2(N__10778),
            .in3(N__10568),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un1_beamylto9_0_LC_5_8_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un1_beamylto9_0_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un1_beamylto9_0_LC_5_8_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 un114_pixel_6_1_5__un1_beamylto9_0_LC_5_8_4 (
            .in0(N__9851),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11796),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un1_beamylto9_3_0_LC_5_8_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un1_beamylto9_3_0_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un1_beamylto9_3_0_LC_5_8_5.LUT_INIT=16'b0000000001110000;
    LogicCell40 un114_pixel_6_1_5__un1_beamylto9_3_0_LC_5_8_5 (
            .in0(N__11330),
            .in1(N__14922),
            .in2(N__9215),
            .in3(N__9501),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un1_beamylto9_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_5_8_6.C_ON=1'b0;
    defparam VSync_1_LC_5_8_6.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_5_8_6.LUT_INIT=16'b1111111111011111;
    LogicCell40 VSync_1_LC_5_8_6 (
            .in0(N__9175),
            .in1(N__9349),
            .in2(N__9212),
            .in3(N__9626),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13141),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un3_beamx_2_LC_5_8_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un3_beamx_2_LC_5_8_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un3_beamx_2_LC_5_8_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_6_1_5__un3_beamx_2_LC_5_8_7 (
            .in0(_gnd_net_),
            .in1(N__10598),
            .in2(_gnd_net_),
            .in3(N__10637),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_20_LC_5_9_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_20_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_20_LC_5_9_0.LUT_INIT=16'b1010101010101000;
    LogicCell40 un114_pixel_6_1_5__g0_20_LC_5_9_0 (
            .in0(N__9624),
            .in1(N__9525),
            .in2(N__8987),
            .in3(N__9348),
            .lcout(un4_beamy_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un5_beamx_4_LC_5_9_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un5_beamx_4_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un5_beamx_4_LC_5_9_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_6_1_5__un5_beamx_4_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(N__9425),
            .in2(_gnd_net_),
            .in3(N__9688),
            .lcout(un8_beamy_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_5_9_3.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_5_9_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_5_9_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_3_LC_5_9_3 (
            .in0(_gnd_net_),
            .in1(N__11780),
            .in2(_gnd_net_),
            .in3(N__11368),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_1_LC_5_9_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_1_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_1_LC_5_9_4.LUT_INIT=16'b0001011101001101;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_1_LC_5_9_4 (
            .in0(N__10212),
            .in1(N__11017),
            .in2(N__9161),
            .in3(N__11059),
            .lcout(),
            .ltout(row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_LC_5_9_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_LC_5_9_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_LC_5_9_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_LC_5_9_5 (
            .in0(N__14279),
            .in1(N__9158),
            .in2(N__9125),
            .in3(N__9062),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_beamylto9_LC_5_9_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_beamylto9_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_beamylto9_LC_5_9_6.LUT_INIT=16'b1010101010101000;
    LogicCell40 un114_pixel_6_1_5__un4_beamylto9_LC_5_9_6 (
            .in0(N__9623),
            .in1(N__9524),
            .in2(N__8986),
            .in3(N__9347),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_1_4_LC_5_10_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_1_4_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_1_4_LC_5_10_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 un114_pixel_6_1_5__g0_1_4_LC_5_10_1 (
            .in0(N__9689),
            .in1(N__9526),
            .in2(N__9431),
            .in3(N__11794),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g0_1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_1_LC_5_10_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_1_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_1_LC_5_10_2.LUT_INIT=16'b1011111100000000;
    LogicCell40 un114_pixel_6_1_5__g0_0_1_LC_5_10_2 (
            .in0(N__9616),
            .in1(N__9224),
            .in2(N__9695),
            .in3(N__14499),
            .lcout(un114_pixel_6_1_5__g0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_4_LC_5_10_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_4_LC_5_10_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_4_LC_5_10_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 un114_pixel_6_1_5__g0_0_4_LC_5_10_5 (
            .in0(N__9690),
            .in1(N__9351),
            .in2(N__9854),
            .in3(N__9615),
            .lcout(un114_pixel_6_1_5__g0_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_3_LC_5_10_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_3_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_3_LC_5_10_6.LUT_INIT=16'b0000000000000101;
    LogicCell40 un114_pixel_6_1_5__g0_0_3_LC_5_10_6 (
            .in0(N__11795),
            .in1(_gnd_net_),
            .in2(N__9530),
            .in3(N__9430),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g0_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_8_LC_5_10_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_8_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_8_LC_5_10_7.LUT_INIT=16'b0010000010100000;
    LogicCell40 un114_pixel_6_1_5__g0_8_LC_5_10_7 (
            .in0(N__9368),
            .in1(N__14854),
            .in2(N__9359),
            .in3(N__11374),
            .lcout(un1_beamy_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g2_0_0_LC_5_11_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g2_0_0_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g2_0_0_LC_5_11_1.LUT_INIT=16'b0000000001100110;
    LogicCell40 un114_pixel_6_1_5__g2_0_0_LC_5_11_1 (
            .in0(N__11332),
            .in1(N__11782),
            .in2(_gnd_net_),
            .in3(N__11672),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g2_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJH2N2P_0_3_LC_5_11_2.C_ON=1'b0;
    defparam beamY_RNIJH2N2P_0_3_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIJH2N2P_0_3_LC_5_11_2.LUT_INIT=16'b0001010111101010;
    LogicCell40 beamY_RNIJH2N2P_0_3_LC_5_11_2 (
            .in0(N__10854),
            .in1(N__9860),
            .in2(N__9356),
            .in3(N__9767),
            .lcout(N_80_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ3MRIJ1_3_LC_5_11_3.C_ON=1'b0;
    defparam beamY_RNIQ3MRIJ1_3_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ3MRIJ1_3_LC_5_11_3.LUT_INIT=16'b0011110000011110;
    LogicCell40 beamY_RNIQ3MRIJ1_3_LC_5_11_3 (
            .in0(N__9953),
            .in1(N__10855),
            .in2(N__11811),
            .in3(N__11673),
            .lcout(m511_0_o2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_1_1_LC_5_11_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_1_1_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_1_1_LC_5_11_4.LUT_INIT=16'b0000000000010101;
    LogicCell40 un114_pixel_6_1_5__g0_0_1_1_LC_5_11_4 (
            .in0(N__9844),
            .in1(N__11333),
            .in2(N__14898),
            .in3(N__9352),
            .lcout(un114_pixel_6_1_5__g0_0_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4VNB7K_1_4_LC_5_11_5.C_ON=1'b0;
    defparam beamY_RNI4VNB7K_1_4_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI4VNB7K_1_4_LC_5_11_5.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI4VNB7K_1_4_LC_5_11_5 (
            .in0(N__10199),
            .in1(N__10305),
            .in2(_gnd_net_),
            .in3(N__10017),
            .lcout(g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_4_LC_5_11_6.C_ON=1'b0;
    defparam beamY_RNIBFP3_4_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_4_LC_5_11_6.LUT_INIT=16'b0110011010101010;
    LogicCell40 beamY_RNIBFP3_4_LC_5_11_6 (
            .in0(N__9843),
            .in1(N__11776),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4VNB7K_4_LC_5_11_7.C_ON=1'b0;
    defparam beamY_RNI4VNB7K_4_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI4VNB7K_4_LC_5_11_7.LUT_INIT=16'b0011110011000011;
    LogicCell40 beamY_RNI4VNB7K_4_LC_5_11_7 (
            .in0(_gnd_net_),
            .in1(N__10306),
            .in2(N__9770),
            .in3(N__10018),
            .lcout(g1_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIITKSF53_3_LC_5_12_0.C_ON=1'b0;
    defparam beamY_RNIITKSF53_3_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIITKSF53_3_LC_5_12_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIITKSF53_3_LC_5_12_0 (
            .in0(N__11589),
            .in1(N__9713),
            .in2(N__11671),
            .in3(N__9747),
            .lcout(m511_0_x2_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ3MRIJ1_0_3_LC_5_12_1.C_ON=1'b0;
    defparam beamY_RNIQ3MRIJ1_0_3_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ3MRIJ1_0_3_LC_5_12_1.LUT_INIT=16'b0100101101011010;
    LogicCell40 beamY_RNIQ3MRIJ1_0_3_LC_5_12_1 (
            .in0(N__10861),
            .in1(N__11658),
            .in2(N__11828),
            .in3(N__9952),
            .lcout(G_7_0_m2_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1KDQIJ1_3_LC_5_12_2.C_ON=1'b0;
    defparam beamY_RNI1KDQIJ1_3_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI1KDQIJ1_3_LC_5_12_2.LUT_INIT=16'b0011001111101110;
    LogicCell40 beamY_RNI1KDQIJ1_3_LC_5_12_2 (
            .in0(N__9951),
            .in1(N__10860),
            .in2(_gnd_net_),
            .in3(N__11659),
            .lcout(),
            .ltout(G_7_0_m2_1_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIABC7E1_3_LC_5_12_3.C_ON=1'b0;
    defparam beamY_RNIABC7E1_3_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIABC7E1_3_LC_5_12_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIABC7E1_3_LC_5_12_3 (
            .in0(N__9749),
            .in1(N__9722),
            .in2(N__9761),
            .in3(N__11590),
            .lcout(),
            .ltout(G_7_0_m2_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGABC8I2_2_LC_5_12_4.C_ON=1'b0;
    defparam beamY_RNIGABC8I2_2_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIGABC8I2_2_LC_5_12_4.LUT_INIT=16'b0001100000100100;
    LogicCell40 beamY_RNIGABC8I2_2_LC_5_12_4 (
            .in0(N__11591),
            .in1(N__11380),
            .in2(N__9758),
            .in3(N__9755),
            .lcout(G_7_0_m2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJH2N2P_3_LC_5_12_5.C_ON=1'b0;
    defparam beamY_RNIJH2N2P_3_LC_5_12_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIJH2N2P_3_LC_5_12_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIJH2N2P_3_LC_5_12_5 (
            .in0(N__9748),
            .in1(N__11657),
            .in2(N__9721),
            .in3(N__9935),
            .lcout(beamY_RNIJH2N2PZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILT8E7K_0_3_LC_5_12_6.C_ON=1'b0;
    defparam beamY_RNILT8E7K_0_3_LC_5_12_6.SEQ_MODE=4'b0000;
    defparam beamY_RNILT8E7K_0_3_LC_5_12_6.LUT_INIT=16'b0110000010010000;
    LogicCell40 beamY_RNILT8E7K_0_3_LC_5_12_6 (
            .in0(N__10295),
            .in1(N__10211),
            .in2(N__10097),
            .in3(N__10019),
            .lcout(chary_if_generate_plus_mult1_un68_sum_ac0_5),
            .ltout(chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIL0E2QG2_3_LC_5_12_7.C_ON=1'b0;
    defparam beamY_RNIL0E2QG2_3_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIL0E2QG2_3_LC_5_12_7.LUT_INIT=16'b0100010110111010;
    LogicCell40 beamY_RNIL0E2QG2_3_LC_5_12_7 (
            .in0(N__10859),
            .in1(N__11653),
            .in2(N__9938),
            .in3(N__11588),
            .lcout(beamY_RNIL0E2QG2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0 (
            .in0(_gnd_net_),
            .in1(N__14334),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_6_4_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_6_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(N__9868),
            .in2(N__9878),
            .in3(N__9923),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_6_4_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_6_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_6_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_6_4_2 (
            .in0(_gnd_net_),
            .in1(N__11878),
            .in2(N__11204),
            .in3(N__9911),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_6_4_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_6_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_6_4_3 (
            .in0(N__9895),
            .in1(N__9869),
            .in2(N__11903),
            .in3(N__9902),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_6_4_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_6_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_6_4_4 (
            .in0(_gnd_net_),
            .in1(N__11891),
            .in2(_gnd_net_),
            .in3(N__9899),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_4_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_6_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13678),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_6_4_6.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_6_4_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_6_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_6_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11877),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_6_4_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_6_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_6_4_7 (
            .in0(N__14335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_6_5_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_6_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14476),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_5_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_5_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10489),
            .in3(N__10343),
            .lcout(charx_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_5_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_5_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10519),
            .in3(N__10340),
            .lcout(charx_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_5_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(N__14236),
            .in2(N__10737),
            .in3(N__10337),
            .lcout(chessboardpixel_un152_pixel_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_5_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_5_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_6_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10773),
            .in3(N__10334),
            .lcout(charx_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_5_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_5_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_6_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10687),
            .in3(N__10331),
            .lcout(charx_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_5_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_6_5_6 (
            .in0(_gnd_net_),
            .in1(N__14237),
            .in2(N__10565),
            .in3(N__10328),
            .lcout(charx_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_5_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_5_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_6_5_7 (
            .in0(_gnd_net_),
            .in1(N__11162),
            .in2(_gnd_net_),
            .in3(N__10325),
            .lcout(charx_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_6_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_6_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_6_6_0 (
            .in0(_gnd_net_),
            .in1(N__14266),
            .in2(N__10635),
            .in3(N__10412),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_6_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_6_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_6_6_1 (
            .in0(_gnd_net_),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__10409),
            .lcout(CO3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_6_6_2.C_ON=1'b0;
    defparam beamX_1_LC_6_6_2.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_6_6_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 beamX_1_LC_6_6_2 (
            .in0(N__14475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10488),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13146),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_1_LC_6_6_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_1_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_1_LC_6_6_3.LUT_INIT=16'b0101011100010101;
    LogicCell40 un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_1_LC_6_6_3 (
            .in0(N__10406),
            .in1(N__10810),
            .in2(N__16325),
            .in3(N__16135),
            .lcout(un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_6_6_5.C_ON=1'b0;
    defparam beamX_0_LC_6_6_5.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_6_6_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_0_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(N__14474),
            .in2(_gnd_net_),
            .in3(N__11507),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13146),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_5_LC_6_7_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_5_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_5_LC_6_7_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_6_1_5__un4_row_5_LC_6_7_1 (
            .in0(N__10400),
            .in1(N__10379),
            .in2(N__11999),
            .in3(N__12362),
            .lcout(un114_pixel_6_1_5__un4_rowZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un3_beamx_5_LC_6_7_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un3_beamx_5_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un3_beamx_5_LC_6_7_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 un114_pixel_6_1_5__un3_beamx_5_LC_6_7_3 (
            .in0(N__10771),
            .in1(N__10517),
            .in2(N__11140),
            .in3(N__10486),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un3_beamx_7_LC_6_7_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un3_beamx_7_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un3_beamx_7_LC_6_7_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 un114_pixel_6_1_5__un3_beamx_7_LC_6_7_4 (
            .in0(N__10563),
            .in1(N__10735),
            .in2(N__10361),
            .in3(N__14500),
            .lcout(un114_pixel_6_1_5__un3_beamxZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g3_0_1_LC_6_7_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g3_0_1_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g3_0_1_LC_6_7_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 un114_pixel_6_1_5__g3_0_1_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(N__10599),
            .in2(_gnd_net_),
            .in3(N__10633),
            .lcout(un114_pixel_6_1_5__g3_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_LC_6_7_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_LC_6_7_6.LUT_INIT=16'b1000001010010010;
    LogicCell40 un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_LC_6_7_6 (
            .in0(N__10820),
            .in1(N__10814),
            .in2(N__10799),
            .in3(N__16145),
            .lcout(chessboardpixel_un174_pixel_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un13_beamylto7_LC_6_8_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un13_beamylto7_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un13_beamylto7_LC_6_8_0.LUT_INIT=16'b1010101010000000;
    LogicCell40 un114_pixel_6_1_5__un13_beamylto7_LC_6_8_0 (
            .in0(N__11173),
            .in1(N__10689),
            .in2(N__10703),
            .in3(N__10567),
            .lcout(un13_beamylt10_0),
            .ltout(un13_beamylt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un15_beamy_LC_6_8_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un15_beamy_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un15_beamy_LC_6_8_1.LUT_INIT=16'b0011000100000000;
    LogicCell40 un114_pixel_6_1_5__un15_beamy_LC_6_8_1 (
            .in0(N__11191),
            .in1(N__10787),
            .in2(N__10781),
            .in3(N__10444),
            .lcout(un15_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un13_beamylto5_1_LC_6_8_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un13_beamylto5_1_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un13_beamylto5_1_LC_6_8_2.LUT_INIT=16'b1010100010001000;
    LogicCell40 un114_pixel_6_1_5__un13_beamylto5_1_LC_6_8_2 (
            .in0(N__10774),
            .in1(N__10738),
            .in2(N__10454),
            .in3(N__14477),
            .lcout(un18_beamylt5_0),
            .ltout(un18_beamylt5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un15_beamy_1_LC_6_8_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un15_beamy_1_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un15_beamy_1_LC_6_8_3.LUT_INIT=16'b0011011100000000;
    LogicCell40 un114_pixel_6_1_5__un15_beamy_1_LC_6_8_3 (
            .in0(N__10688),
            .in1(N__10529),
            .in2(N__10646),
            .in3(N__10643),
            .lcout(un114_pixel_6_1_5__un15_beamyZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un18_beamylto9_2_LC_6_8_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un18_beamylto9_2_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un18_beamylto9_2_LC_6_8_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_6_1_5__un18_beamylto9_2_LC_6_8_4 (
            .in0(N__11172),
            .in1(N__10636),
            .in2(N__10601),
            .in3(N__10566),
            .lcout(un114_pixel_6_1_5__un18_beamylto9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un13_beamylto2_0_LC_6_8_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un13_beamylto2_0_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un13_beamylto2_0_LC_6_8_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 un114_pixel_6_1_5__un13_beamylto2_0_LC_6_8_5 (
            .in0(N__10523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10490),
            .lcout(un114_pixel_6_1_5__un13_beamylto2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_19_LC_6_8_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_19_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_19_LC_6_8_6.LUT_INIT=16'b0010001000100000;
    LogicCell40 un114_pixel_6_1_5__g0_19_LC_6_8_6 (
            .in0(N__10445),
            .in1(N__10436),
            .in2(N__10430),
            .in3(N__10418),
            .lcout(un114_pixel_6_1_5__g0_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_6_8_7.C_ON=1'b0;
    defparam HSync_1_LC_6_8_7.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_6_8_7.LUT_INIT=16'b1111111111111101;
    LogicCell40 HSync_1_LC_6_8_7 (
            .in0(N__11192),
            .in1(N__11174),
            .in2(N__11141),
            .in3(N__11108),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13144),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_7_LC_6_9_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_7_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_7_LC_6_9_3.LUT_INIT=16'b0000000000101000;
    LogicCell40 un114_pixel_6_1_5__un4_row_7_LC_6_9_3 (
            .in0(N__11069),
            .in1(N__11060),
            .in2(N__11024),
            .in3(N__12434),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_LC_6_9_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_LC_6_9_4.LUT_INIT=16'b1000000000100000;
    LogicCell40 un114_pixel_6_1_5__un4_row_LC_6_9_4 (
            .in0(N__10985),
            .in1(N__10973),
            .in2(N__10967),
            .in3(N__10964),
            .lcout(un4_row),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_LC_6_9_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_LC_6_9_5.LUT_INIT=16'b1000000001000000;
    LogicCell40 un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_LC_6_9_5 (
            .in0(N__10955),
            .in1(N__10928),
            .in2(N__14905),
            .in3(N__10915),
            .lcout(),
            .ltout(chessboardpixel_un200_pixellt10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto10_1_LC_6_9_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto10_1_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__chessboardpixel_un200_pixellto10_1_LC_6_9_6.LUT_INIT=16'b0000001100001001;
    LogicCell40 un114_pixel_6_1_5__chessboardpixel_un200_pixellto10_1_LC_6_9_6 (
            .in0(N__10916),
            .in1(N__10892),
            .in2(N__10880),
            .in3(N__10877),
            .lcout(chessboardpixel_un200_pixel_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_6_10_0.C_ON=1'b0;
    defparam beamY_1_LC_6_10_0.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_6_10_0.LUT_INIT=16'b0100010001101100;
    LogicCell40 beamY_1_LC_6_10_0 (
            .in0(N__11542),
            .in1(N__14855),
            .in2(N__15143),
            .in3(N__11448),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13143),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_1_LC_6_11_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_1_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_1_LC_6_11_0.LUT_INIT=16'b1010010110010110;
    LogicCell40 un114_pixel_6_1_5__g0_1_LC_6_11_0 (
            .in0(N__11603),
            .in1(N__11615),
            .in2(N__11830),
            .in3(N__10865),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_0_LC_6_11_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_0_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_0_LC_6_11_1.LUT_INIT=16'b0111101010011110;
    LogicCell40 un114_pixel_6_1_5__g0_0_0_LC_6_11_1 (
            .in0(N__14847),
            .in1(N__11370),
            .in2(N__10823),
            .in3(N__11216),
            .lcout(un114_pixel_6_1_5__font_un126_pixel_m_4_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g2_LC_6_11_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g2_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g2_LC_6_11_2.LUT_INIT=16'b0000000001001000;
    LogicCell40 un114_pixel_6_1_5__g2_LC_6_11_2 (
            .in0(N__11369),
            .in1(N__11837),
            .in2(N__11829),
            .in3(N__11678),
            .lcout(g2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_12_LC_6_11_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_12_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_12_LC_6_11_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 un114_pixel_6_1_5__g0_12_LC_6_11_4 (
            .in0(N__12536),
            .in1(N__15107),
            .in2(_gnd_net_),
            .in3(N__13248),
            .lcout(N_357_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPG1SS93_2_LC_6_11_5.C_ON=1'b0;
    defparam beamY_RNIPG1SS93_2_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIPG1SS93_2_LC_6_11_5.LUT_INIT=16'b0000011010010000;
    LogicCell40 beamY_RNIPG1SS93_2_LC_6_11_5 (
            .in0(N__11609),
            .in1(N__11602),
            .in2(N__11381),
            .in3(N__11561),
            .lcout(beamY_RNIPG1SS93Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_13_0.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_13_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_6_13_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_i_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16439),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_6_13_2.C_ON=1'b0;
    defparam beamY_0_LC_6_13_2.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_6_13_2.LUT_INIT=16'b0010001001100110;
    LogicCell40 beamY_0_LC_6_13_2 (
            .in0(N__15052),
            .in1(N__11553),
            .in2(_gnd_net_),
            .in3(N__11449),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13148),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_6_LC_6_13_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_6_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_6_LC_6_13_3.LUT_INIT=16'b0100010000100010;
    LogicCell40 un114_pixel_6_1_5__g0_6_LC_6_13_3 (
            .in0(N__11379),
            .in1(N__11225),
            .in2(_gnd_net_),
            .in3(N__11215),
            .lcout(font_un28_pixel_0_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13693),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_7_3_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_7_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__11854),
            .in2(N__11864),
            .in3(N__11195),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_7_3_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_7_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__12629),
            .in2(N__12596),
            .in3(N__11894),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_7_3_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_7_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_7_3_3 (
            .in0(N__11879),
            .in1(N__11855),
            .in2(N__12620),
            .in3(N__11885),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_7_3_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_7_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__12608),
            .in2(_gnd_net_),
            .in3(N__11882),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_7_3_6.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_7_3_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_7_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_1_LC_7_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13614),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_7_3_7.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_7_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12591),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_4_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__14329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_m_2_LC_7_4_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_2_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_2_LC_7_4_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_m_2_LC_7_4_1 (
            .in0(N__12713),
            .in1(N__13945),
            .in2(N__11942),
            .in3(N__11846),
            .lcout(if_generate_plus_mult1_un47_sum_m_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_4_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__11933),
            .in2(N__12293),
            .in3(N__11843),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_4_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__13946),
            .in2(N__12284),
            .in3(N__11840),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_4_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_4_4.LUT_INIT=16'b1000000001111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_4_4 (
            .in0(N__13947),
            .in1(N__13609),
            .in2(N__13685),
            .in3(N__11948),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_5),
            .ltout(column_1_if_generate_plus_mult1_un47_sum1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_571_i_LC_7_4_5.C_ON=1'b0;
    defparam column_1_N_571_i_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam column_1_N_571_i_LC_7_4_5.LUT_INIT=16'b0011001100001111;
    LogicCell40 column_1_N_571_i_LC_7_4_5 (
            .in0(_gnd_net_),
            .in1(N__12766),
            .in2(N__11945),
            .in3(N__13948),
            .lcout(N_571_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_7_4_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_7_4_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_7_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_3_LC_7_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13667),
            .lcout(un5_visiblex_i_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_7_5_0.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_7_5_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_3_LC_7_5_0 (
            .in0(N__13888),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un26_sum_axb_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_7_5_1.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_7_5_1.LUT_INIT=16'b1001100111000011;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_7_5_1 (
            .in0(N__12692),
            .in1(N__11974),
            .in2(N__11927),
            .in3(N__13893),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_7_5_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_7_5_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_m_5_LC_7_5_2 (
            .in0(N__13891),
            .in1(_gnd_net_),
            .in2(N__12748),
            .in3(N__12765),
            .lcout(if_generate_plus_mult1_un47_sum_m_5),
            .ltout(if_generate_plus_mult1_un47_sum_m_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_5_3.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_5_3.LUT_INIT=16'b1100001110100101;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_5_3 (
            .in0(N__11915),
            .in1(N__12701),
            .in2(N__11909),
            .in3(N__13892),
            .lcout(),
            .ltout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_5_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_5_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11906),
            .in3(N__12396),
            .lcout(if_generate_plus_mult1_un54_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_7_5_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_7_5_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_2_LC_7_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13887),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m15_LC_7_5_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m15_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m15_LC_7_5_6.LUT_INIT=16'b0110011010011001;
    LogicCell40 un114_pixel_6_1_5__m15_LC_7_5_6 (
            .in0(N__13889),
            .in1(N__13671),
            .in2(_gnd_net_),
            .in3(N__13591),
            .lcout(N_11_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_7_5_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_7_5_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_7_5_7.LUT_INIT=16'b0101111100110011;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_7_5_7 (
            .in0(N__13592),
            .in1(N__13552),
            .in2(N__13686),
            .in3(N__13890),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_m_1_LC_7_6_1.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_1_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_1_LC_7_6_1.LUT_INIT=16'b0011001100001111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_m_1_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__14330),
            .in2(N__14345),
            .in3(N__13886),
            .lcout(if_generate_plus_mult1_un47_sum_m_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_6_2.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_6_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13666),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_2_LC_7_6_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_2_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_2_LC_7_6_3.LUT_INIT=16'b0000000001110000;
    LogicCell40 un114_pixel_6_1_5__un4_row_2_LC_7_6_3 (
            .in0(N__12275),
            .in1(N__12175),
            .in2(N__12731),
            .in3(N__12113),
            .lcout(un114_pixel_6_1_5__un4_rowZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_7_6_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_7_6_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13918),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un26_sum_s_2_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_7_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__15285),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_7_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__12403),
            .in2(N__11990),
            .in3(N__11981),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_7_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(N__11978),
            .in2(N__11963),
            .in3(N__11951),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_7_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_7_3 (
            .in0(N__12360),
            .in1(N__12416),
            .in2(N__12407),
            .in3(N__12383),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_7_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__12380),
            .in2(_gnd_net_),
            .in3(N__12371),
            .lcout(if_generate_plus_mult1_un54_sum_s_5),
            .ltout(if_generate_plus_mult1_un54_sum_s_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_7_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12368),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__16156),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__12331),
            .in2(N__12302),
            .in3(N__12365),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__12361),
            .in2(N__12344),
            .in3(N__12335),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3 (
            .in0(N__15385),
            .in1(N__12332),
            .in2(N__12323),
            .in3(N__12314),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__12311),
            .in2(_gnd_net_),
            .in3(N__12305),
            .lcout(un5_rowlto3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_562_i_LC_7_8_5.C_ON=1'b0;
    defparam column_1_N_562_i_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam column_1_N_562_i_LC_7_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_N_562_i_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15286),
            .lcout(N_562_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__Pixel_3_sqmuxa_LC_7_9_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__Pixel_3_sqmuxa_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__Pixel_3_sqmuxa_LC_7_9_1.LUT_INIT=16'b0001000001000000;
    LogicCell40 un114_pixel_6_1_5__Pixel_3_sqmuxa_LC_7_9_1 (
            .in0(N__13039),
            .in1(N__12449),
            .in2(N__12892),
            .in3(N__12440),
            .lcout(Pixel_3_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_rowlto3_sbtinv_LC_7_9_5.C_ON=1'b0;
    defparam un5_rowlto3_sbtinv_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam un5_rowlto3_sbtinv_LC_7_9_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_rowlto3_sbtinv_LC_7_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15383),
            .lcout(un5_rowlto3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_9_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_i_LC_7_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16157),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_7_1_LC_7_9_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_7_1_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_7_1_LC_7_9_7.LUT_INIT=16'b0000000001110111;
    LogicCell40 un114_pixel_6_1_5__un4_row_7_1_LC_7_9_7 (
            .in0(N__15685),
            .in1(N__16014),
            .in2(_gnd_net_),
            .in3(N__15384),
            .lcout(un114_pixel_6_1_5__un4_row_7Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI59CM492_LC_7_10_2.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI59CM492_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI59CM492_LC_7_10_2.LUT_INIT=16'b0101010111110011;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI59CM492_LC_7_10_2 (
            .in0(N__12428),
            .in1(N__16017),
            .in2(N__15233),
            .in3(N__13380),
            .lcout(),
            .ltout(N_18_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6M26DQ1_1_LC_7_10_3.C_ON=1'b0;
    defparam beamY_RNI6M26DQ1_1_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI6M26DQ1_1_LC_7_10_3.LUT_INIT=16'b1010111100000101;
    LogicCell40 beamY_RNI6M26DQ1_1_LC_7_10_3 (
            .in0(N__14848),
            .in1(_gnd_net_),
            .in2(N__12422),
            .in3(N__12461),
            .lcout(N_23_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7LRQVE2_0_LC_7_10_4.C_ON=1'b0;
    defparam beamY_RNI7LRQVE2_0_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI7LRQVE2_0_LC_7_10_4.LUT_INIT=16'b0001111101110111;
    LogicCell40 beamY_RNI7LRQVE2_0_LC_7_10_4 (
            .in0(N__13097),
            .in1(N__16016),
            .in2(N__15162),
            .in3(N__13379),
            .lcout(),
            .ltout(N_7_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQVAMG32_1_LC_7_10_5.C_ON=1'b0;
    defparam beamY_RNIQVAMG32_1_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIQVAMG32_1_LC_7_10_5.LUT_INIT=16'b1000110110001101;
    LogicCell40 beamY_RNIQVAMG32_1_LC_7_10_5 (
            .in0(N__14849),
            .in1(N__12479),
            .in2(N__12419),
            .in3(_gnd_net_),
            .lcout(N_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_9_LC_7_10_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_9_LC_7_10_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_9_LC_7_10_6.LUT_INIT=16'b0000010001011111;
    LogicCell40 un114_pixel_6_1_5__g0_9_LC_7_10_6 (
            .in0(N__15862),
            .in1(N__14729),
            .in2(N__14929),
            .in3(N__16018),
            .lcout(),
            .ltout(un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_2_LC_7_10_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_2_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_2_LC_7_10_7.LUT_INIT=16'b1011110100100100;
    LogicCell40 un114_pixel_6_1_5__g0_2_LC_7_10_7 (
            .in0(N__14850),
            .in1(N__12494),
            .in2(N__12482),
            .in3(N__13253),
            .lcout(N_342_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISS6QGK3_0_LC_7_11_0.C_ON=1'b0;
    defparam beamY_RNISS6QGK3_0_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam beamY_RNISS6QGK3_0_LC_7_11_0.LUT_INIT=16'b1001100100001111;
    LogicCell40 beamY_RNISS6QGK3_0_LC_7_11_0 (
            .in0(N__12518),
            .in1(N__15106),
            .in2(N__12503),
            .in3(N__13374),
            .lcout(N_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m24_LC_7_11_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m24_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m24_LC_7_11_1.LUT_INIT=16'b0000000000010001;
    LogicCell40 un114_pixel_6_1_5__m24_LC_7_11_1 (
            .in0(N__15857),
            .in1(N__15665),
            .in2(_gnd_net_),
            .in3(N__16009),
            .lcout(column_0111_0),
            .ltout(column_0111_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI05CI5A3_0_0_LC_7_11_2.C_ON=1'b0;
    defparam beamY_RNI05CI5A3_0_0_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI05CI5A3_0_0_LC_7_11_2.LUT_INIT=16'b0000111111001100;
    LogicCell40 beamY_RNI05CI5A3_0_0_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(N__14382),
            .in2(N__12473),
            .in3(N__15101),
            .lcout(),
            .ltout(beamY_RNI05CI5A3_0Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBABJS01_1_LC_7_11_3.C_ON=1'b0;
    defparam beamY_RNIBABJS01_1_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIBABJS01_1_LC_7_11_3.LUT_INIT=16'b1111110001110100;
    LogicCell40 beamY_RNIBABJS01_1_LC_7_11_3 (
            .in0(N__15102),
            .in1(N__14935),
            .in2(N__12470),
            .in3(N__12566),
            .lcout(),
            .ltout(beamY_RNIBABJS01Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__font_un126_pixel_2_am_LC_7_11_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__font_un126_pixel_2_am_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__font_un126_pixel_2_am_LC_7_11_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 un114_pixel_6_1_5__font_un126_pixel_2_am_LC_7_11_4 (
            .in0(_gnd_net_),
            .in1(N__12644),
            .in2(N__12467),
            .in3(N__13373),
            .lcout(font_un126_pixel_2_am),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2QTJEJ1_0_LC_7_11_5.C_ON=1'b0;
    defparam beamY_RNI2QTJEJ1_0_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI2QTJEJ1_0_LC_7_11_5.LUT_INIT=16'b0000001010010001;
    LogicCell40 beamY_RNI2QTJEJ1_0_LC_7_11_5 (
            .in0(N__15858),
            .in1(N__15666),
            .in2(N__15145),
            .in3(N__16010),
            .lcout(),
            .ltout(N_21_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIAVDE8H3_0_LC_7_11_6.C_ON=1'b0;
    defparam beamY_RNIAVDE8H3_0_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIAVDE8H3_0_LC_7_11_6.LUT_INIT=16'b1111000000110011;
    LogicCell40 beamY_RNIAVDE8H3_0_LC_7_11_6 (
            .in0(_gnd_net_),
            .in1(N__15200),
            .in2(N__12464),
            .in3(N__13372),
            .lcout(N_22_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNINIKJ5A3_1_LC_7_11_7.C_ON=1'b0;
    defparam beamY_RNINIKJ5A3_1_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam beamY_RNINIKJ5A3_1_LC_7_11_7.LUT_INIT=16'b1000111010111110;
    LogicCell40 beamY_RNINIKJ5A3_1_LC_7_11_7 (
            .in0(N__14383),
            .in1(N__14934),
            .in2(N__15144),
            .in3(N__12455),
            .lcout(beamY_RNINIKJ5A3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_3_bm_6_LC_7_12_0.C_ON=1'b0;
    defparam un116_pixel_3_bm_6_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_3_bm_6_LC_7_12_0.LUT_INIT=16'b1100011101000111;
    LogicCell40 un116_pixel_3_bm_6_LC_7_12_0 (
            .in0(N__15662),
            .in1(N__16048),
            .in2(N__15854),
            .in3(N__15481),
            .lcout(),
            .ltout(un116_pixel_3_bmZ0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISJITRQ2_1_LC_7_12_1.C_ON=1'b0;
    defparam beamY_RNISJITRQ2_1_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam beamY_RNISJITRQ2_1_LC_7_12_1.LUT_INIT=16'b1010000001110111;
    LogicCell40 beamY_RNISJITRQ2_1_LC_7_12_1 (
            .in0(N__14936),
            .in1(N__12542),
            .in2(N__12524),
            .in3(N__12509),
            .lcout(),
            .ltout(beamY_RNISJITRQ2Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJDHE4C2_1_LC_7_12_2.C_ON=1'b0;
    defparam beamY_RNIJDHE4C2_1_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIJDHE4C2_1_LC_7_12_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 beamY_RNIJDHE4C2_1_LC_7_12_2 (
            .in0(N__12548),
            .in1(_gnd_net_),
            .in2(N__12521),
            .in3(N__13371),
            .lcout(beamY_RNIJDHE4C2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam m11_LC_7_12_3.C_ON=1'b0;
    defparam m11_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam m11_LC_7_12_3.LUT_INIT=16'b0010110000000000;
    LogicCell40 m11_LC_7_12_3 (
            .in0(N__15479),
            .in1(N__15806),
            .in2(N__16083),
            .in3(N__15663),
            .lcout(N_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un114_pixel_3_i_m2_6_LC_7_12_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un114_pixel_3_i_m2_6_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un114_pixel_3_i_m2_6_LC_7_12_4.LUT_INIT=16'b1001011010011110;
    LogicCell40 un114_pixel_6_1_5__un114_pixel_3_i_m2_6_LC_7_12_4 (
            .in0(N__15660),
            .in1(N__16038),
            .in2(N__15853),
            .in3(N__15477),
            .lcout(un114_pixel_7_1_7__N_11_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m26_LC_7_12_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m26_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m26_LC_7_12_5.LUT_INIT=16'b1010000010000000;
    LogicCell40 un114_pixel_6_1_5__m26_LC_7_12_5 (
            .in0(N__15478),
            .in1(N__15799),
            .in2(N__16082),
            .in3(N__15661),
            .lcout(),
            .ltout(N_248_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9GDVDD3_1_LC_7_12_6.C_ON=1'b0;
    defparam beamY_RNI9GDVDD3_1_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI9GDVDD3_1_LC_7_12_6.LUT_INIT=16'b0010011000110111;
    LogicCell40 beamY_RNI9GDVDD3_1_LC_7_12_6 (
            .in0(N__14873),
            .in1(N__15037),
            .in2(N__12512),
            .in3(N__13247),
            .lcout(un116_pixel_3_ns_1_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam m8_e_LC_7_12_7.C_ON=1'b0;
    defparam m8_e_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam m8_e_LC_7_12_7.LUT_INIT=16'b0010111100000000;
    LogicCell40 m8_e_LC_7_12_7 (
            .in0(N__15480),
            .in1(N__15807),
            .in2(N__16084),
            .in3(N__15664),
            .lcout(N_25_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__column_0001_0_LC_7_13_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__column_0001_0_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__column_0001_0_LC_7_13_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 un114_pixel_6_1_5__column_0001_0_LC_7_13_0 (
            .in0(N__16051),
            .in1(N__15655),
            .in2(N__15856),
            .in3(N__15471),
            .lcout(column_0001_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un114_pixel_3_i_a3_7_LC_7_13_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un114_pixel_3_i_a3_7_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un114_pixel_3_i_a3_7_LC_7_13_1.LUT_INIT=16'b0100010010001000;
    LogicCell40 un114_pixel_6_1_5__un114_pixel_3_i_a3_7_LC_7_13_1 (
            .in0(N__15656),
            .in1(N__15813),
            .in2(_gnd_net_),
            .in3(N__16053),
            .lcout(),
            .ltout(un114_pixel_3_i_a3_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI05CI5A3_0_LC_7_13_2.C_ON=1'b0;
    defparam beamY_RNI05CI5A3_0_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI05CI5A3_0_LC_7_13_2.LUT_INIT=16'b0011111100001100;
    LogicCell40 beamY_RNI05CI5A3_0_LC_7_13_2 (
            .in0(_gnd_net_),
            .in1(N__15036),
            .in2(N__12569),
            .in3(N__12562),
            .lcout(beamY_RNI05CI5A3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2QTJEJ1_0_0_LC_7_13_3.C_ON=1'b0;
    defparam beamY_RNI2QTJEJ1_0_0_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI2QTJEJ1_0_0_LC_7_13_3.LUT_INIT=16'b0000000010010001;
    LogicCell40 beamY_RNI2QTJEJ1_0_0_LC_7_13_3 (
            .in0(N__15653),
            .in1(N__15811),
            .in2(N__15097),
            .in3(N__16052),
            .lcout(),
            .ltout(un116_pixel_3_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDVSK5A3_1_LC_7_13_4.C_ON=1'b0;
    defparam beamY_RNIDVSK5A3_1_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIDVSK5A3_1_LC_7_13_4.LUT_INIT=16'b0001010000110110;
    LogicCell40 beamY_RNIDVSK5A3_1_LC_7_13_4 (
            .in0(N__14908),
            .in1(N__15035),
            .in2(N__12551),
            .in3(N__14380),
            .lcout(beamY_RNIDVSK5A3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m12_LC_7_13_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m12_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m12_LC_7_13_6.LUT_INIT=16'b0100110001000100;
    LogicCell40 un114_pixel_6_1_5__m12_LC_7_13_6 (
            .in0(N__16050),
            .in1(N__15654),
            .in2(N__15855),
            .in3(N__15470),
            .lcout(N_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_15_LC_7_13_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_15_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_15_LC_7_13_7.LUT_INIT=16'b0010000011000000;
    LogicCell40 un114_pixel_6_1_5__g0_15_LC_7_13_7 (
            .in0(N__15469),
            .in1(N__15812),
            .in2(N__15684),
            .in3(N__16049),
            .lcout(un114_pixel_0_1__N_6_mux_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_4_bm_1_LC_7_14_0.C_ON=1'b0;
    defparam un116_pixel_4_bm_1_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_4_bm_1_LC_7_14_0.LUT_INIT=16'b1011011010111110;
    LogicCell40 un116_pixel_4_bm_1_LC_7_14_0 (
            .in0(N__16080),
            .in1(N__15594),
            .in2(N__15864),
            .in3(N__15473),
            .lcout(un116_pixel_4_bmZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_1_am_1_LC_7_14_2.C_ON=1'b0;
    defparam un116_pixel_1_am_1_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam un116_pixel_1_am_1_LC_7_14_2.LUT_INIT=16'b1010011111110111;
    LogicCell40 un116_pixel_1_am_1_LC_7_14_2 (
            .in0(N__16079),
            .in1(N__14723),
            .in2(N__15863),
            .in3(N__15593),
            .lcout(),
            .ltout(un116_pixel_1_amZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUEM1HF2_1_LC_7_14_3.C_ON=1'b0;
    defparam beamY_RNIUEM1HF2_1_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIUEM1HF2_1_LC_7_14_3.LUT_INIT=16'b0010001101100111;
    LogicCell40 beamY_RNIUEM1HF2_1_LC_7_14_3 (
            .in0(N__14906),
            .in1(N__15000),
            .in2(N__12527),
            .in3(N__12635),
            .lcout(un116_pixel_3_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_7_14_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_7_14_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_i_LC_7_14_4 (
            .in0(N__16343),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_4_am_1_LC_7_14_5.C_ON=1'b0;
    defparam un116_pixel_4_am_1_LC_7_14_5.SEQ_MODE=4'b0000;
    defparam un116_pixel_4_am_1_LC_7_14_5.LUT_INIT=16'b1000111100110011;
    LogicCell40 un116_pixel_4_am_1_LC_7_14_5 (
            .in0(N__15474),
            .in1(N__15835),
            .in2(N__15659),
            .in3(N__16081),
            .lcout(),
            .ltout(un116_pixel_4_amZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHIRVUS1_1_LC_7_14_6.C_ON=1'b0;
    defparam beamY_RNIHIRVUS1_1_LC_7_14_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIHIRVUS1_1_LC_7_14_6.LUT_INIT=16'b1010000011011101;
    LogicCell40 beamY_RNIHIRVUS1_1_LC_7_14_6 (
            .in0(N__14907),
            .in1(N__12659),
            .in2(N__12653),
            .in3(N__12650),
            .lcout(beamY_RNIHIRVUS1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_1_bm_1_LC_7_14_7.C_ON=1'b0;
    defparam un116_pixel_1_bm_1_LC_7_14_7.SEQ_MODE=4'b0000;
    defparam un116_pixel_1_bm_1_LC_7_14_7.LUT_INIT=16'b1010110000000011;
    LogicCell40 un116_pixel_1_bm_1_LC_7_14_7 (
            .in0(N__15472),
            .in1(N__15828),
            .in2(N__15658),
            .in3(N__16078),
            .lcout(un116_pixel_1_bmZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_3_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__13613),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_8_3_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_8_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(N__12577),
            .in2(N__12722),
            .in3(N__12623),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_8_3_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_8_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(N__13736),
            .in2(N__13757),
            .in3(N__12611),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_8_3_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_8_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_8_3_3 (
            .in0(N__12595),
            .in1(N__12578),
            .in2(N__13724),
            .in3(N__12602),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_8_3_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_8_3_4.LUT_INIT=16'b0110011010011001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_8_3_4 (
            .in0(N__13756),
            .in1(N__13712),
            .in2(_gnd_net_),
            .in3(N__12599),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_8_3_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_8_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13752),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_8_3_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_8_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13956),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_8_4_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_8_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__14350),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_4_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__12674),
            .in2(N__12776),
            .in3(N__12704),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_4_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__12680),
            .in2(N__12785),
            .in3(N__12695),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_4_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(N__13742),
            .in2(N__12668),
            .in3(N__12686),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_4_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_4_4 (
            .in0(_gnd_net_),
            .in1(N__13955),
            .in2(_gnd_net_),
            .in3(N__12683),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_4_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_4_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_4_5 (
            .in0(N__13953),
            .in1(_gnd_net_),
            .in2(N__13550),
            .in3(_gnd_net_),
            .lcout(if_generate_plus_mult1_un47_sum_0_cry_3_ma),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_4_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_4_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_4_6.LUT_INIT=16'b0011001111111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_4_6 (
            .in0(N__13694),
            .in1(N__13535),
            .in2(_gnd_net_),
            .in3(N__13952),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__N_200_0_i_LC_8_4_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__N_200_0_i_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__N_200_0_i_LC_8_4_7.LUT_INIT=16'b0101111101011111;
    LogicCell40 un114_pixel_6_1_5__N_200_0_i_LC_8_4_7 (
            .in0(N__13954),
            .in1(_gnd_net_),
            .in2(N__13551),
            .in3(_gnd_net_),
            .lcout(N_200_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_8_5_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_8_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_8_5_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_8_5_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_8_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12815),
            .in3(N__12806),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_8_5_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_8_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_8_5_2 (
            .in0(_gnd_net_),
            .in1(N__14184),
            .in2(N__12803),
            .in3(N__12794),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_8_5_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_8_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_8_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13961),
            .in3(N__12791),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_8_5_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_8_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_8_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12788),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_5_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_5_5.LUT_INIT=16'b0110011001100110;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_5_5 (
            .in0(N__13684),
            .in1(N__13507),
            .in2(N__13553),
            .in3(N__13960),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_5_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_8_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_2_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13683),
            .lcout(un5_visiblex_i_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un4_row_0_LC_8_5_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un4_row_0_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un4_row_0_LC_8_5_7.LUT_INIT=16'b1000100011110000;
    LogicCell40 un114_pixel_6_1_5__un4_row_0_LC_8_5_7 (
            .in0(N__13546),
            .in1(N__12767),
            .in2(N__12749),
            .in3(N__13959),
            .lcout(un114_pixel_6_1_5__un4_rowZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_6_1.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_6_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13605),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_8_3.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16446),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_5_bm_6_LC_8_8_4.C_ON=1'b0;
    defparam un116_pixel_5_bm_6_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam un116_pixel_5_bm_6_LC_8_8_4.LUT_INIT=16'b1101111100111100;
    LogicCell40 un116_pixel_5_bm_6_LC_8_8_4 (
            .in0(N__15411),
            .in1(N__15869),
            .in2(N__16086),
            .in3(N__15682),
            .lcout(un116_pixel_5_bmZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_5_am_6_LC_8_8_5.C_ON=1'b0;
    defparam un116_pixel_5_am_6_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam un116_pixel_5_am_6_LC_8_8_5.LUT_INIT=16'b1101011011011110;
    LogicCell40 un116_pixel_5_am_6_LC_8_8_5 (
            .in0(N__15683),
            .in1(N__16070),
            .in2(N__15875),
            .in3(N__15412),
            .lcout(),
            .ltout(un116_pixel_5_amZ0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII25UDD3_0_0_LC_8_8_6.C_ON=1'b0;
    defparam beamY_RNII25UDD3_0_0_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNII25UDD3_0_0_LC_8_8_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNII25UDD3_0_0_LC_8_8_6 (
            .in0(_gnd_net_),
            .in1(N__15166),
            .in2(N__12902),
            .in3(N__12899),
            .lcout(beamY_RNII25UDD3_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_LC_8_9_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_LC_8_9_0.LUT_INIT=16'b1010101010001000;
    LogicCell40 un114_pixel_6_1_5__font_un126_pixel_m_1_LC_8_9_0 (
            .in0(N__12893),
            .in1(N__14545),
            .in2(_gnd_net_),
            .in3(N__13387),
            .lcout(),
            .ltout(un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_0_LC_8_9_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_0_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_0_LC_8_9_1.LUT_INIT=16'b0010000010000000;
    LogicCell40 un114_pixel_6_1_5__g0_0_LC_8_9_1 (
            .in0(N__12872),
            .in1(N__14537),
            .in2(N__12860),
            .in3(N__14582),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g0_2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_LC_8_9_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_LC_8_9_2.LUT_INIT=16'b1100000000000000;
    LogicCell40 un114_pixel_6_1_5__g0_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__12857),
            .in2(N__12845),
            .in3(N__13046),
            .lcout(Pixel_1_r_sn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g1_0_LC_8_9_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g1_0_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g1_0_LC_8_9_3.LUT_INIT=16'b1111101011111010;
    LogicCell40 un114_pixel_6_1_5__g1_0_LC_8_9_3 (
            .in0(N__13388),
            .in1(_gnd_net_),
            .in2(N__14549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(un114_pixel_6_1_5__g1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_16_LC_8_9_4.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_16_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_16_LC_8_9_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_6_1_5__g0_16_LC_8_9_4 (
            .in0(N__12842),
            .in1(N__12830),
            .in2(N__12818),
            .in3(N__13045),
            .lcout(un114_pixel_6_1_5__font_un126_pixel_m_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP6FOQ73_1_LC_8_9_5.C_ON=1'b0;
    defparam beamY_RNIP6FOQ73_1_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIP6FOQ73_1_LC_8_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 beamY_RNIP6FOQ73_1_LC_8_9_5 (
            .in0(N__13028),
            .in1(N__13016),
            .in2(_gnd_net_),
            .in3(N__13010),
            .lcout(),
            .ltout(N_1045_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_i_m2_0_LC_8_9_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_i_m2_0_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_i_m2_0_LC_8_9_6.LUT_INIT=16'b1110010011110000;
    LogicCell40 un114_pixel_6_1_5__g0_i_m2_0_LC_8_9_6 (
            .in0(N__15142),
            .in1(N__13004),
            .in2(N__12998),
            .in3(N__14087),
            .lcout(N_396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_10_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__16339),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_10_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__12964),
            .in2(N__12995),
            .in3(N__12986),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_10_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__15413),
            .in2(N__12983),
            .in3(N__12968),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_10_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_10_3 (
            .in0(N__16003),
            .in1(N__12965),
            .in2(N__12956),
            .in3(N__12944),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_10_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(N__12941),
            .in2(_gnd_net_),
            .in3(N__12932),
            .lcout(un5_rowlto2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_3_LC_8_10_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_3_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_3_LC_8_10_5.LUT_INIT=16'b0000111000001010;
    LogicCell40 un114_pixel_6_1_5__g0_3_LC_8_10_5 (
            .in0(N__12929),
            .in1(N__12923),
            .in2(N__12917),
            .in3(N__13076),
            .lcout(),
            .ltout(Pixel_1_r_rn_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_8_10_6.C_ON=1'b0;
    defparam Pixel_1_LC_8_10_6.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_8_10_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 Pixel_1_LC_8_10_6 (
            .in0(_gnd_net_),
            .in1(N__13193),
            .in2(N__13187),
            .in3(N__13184),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13147),
            .ce(),
            .sr(_gnd_net_));
    defparam m6_1_LC_8_10_7.C_ON=1'b0;
    defparam m6_1_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam m6_1_LC_8_10_7.LUT_INIT=16'b0010100000111100;
    LogicCell40 m6_1_LC_8_10_7 (
            .in0(N__15414),
            .in1(N__15686),
            .in2(N__15873),
            .in3(N__16015),
            .lcout(m6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI1M3Q1V2_0_LC_8_11_0.C_ON=1'b0;
    defparam beamX_RNI1M3Q1V2_0_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam beamX_RNI1M3Q1V2_0_LC_8_11_0.LUT_INIT=16'b0101010111011000;
    LogicCell40 beamX_RNI1M3Q1V2_0_LC_8_11_0 (
            .in0(N__13064),
            .in1(N__13205),
            .in2(N__13325),
            .in3(N__14504),
            .lcout(),
            .ltout(beamX_RNI1M3Q1V2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIB75H7E_0_LC_8_11_1.C_ON=1'b0;
    defparam beamX_RNIB75H7E_0_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam beamX_RNIB75H7E_0_LC_8_11_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 beamX_RNIB75H7E_0_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(N__13091),
            .in2(N__13079),
            .in3(N__13259),
            .lcout(N_1039_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_8_11_2.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_8_11_2.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_8_11_2 (
            .in0(N__14533),
            .in1(N__14412),
            .in2(_gnd_net_),
            .in3(N__14578),
            .lcout(font_un3_pixel_29),
            .ltout(font_un3_pixel_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI440R9C_0_LC_8_11_3.C_ON=1'b0;
    defparam beamX_RNI440R9C_0_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam beamX_RNI440R9C_0_LC_8_11_3.LUT_INIT=16'b0000111101100110;
    LogicCell40 beamX_RNI440R9C_0_LC_8_11_3 (
            .in0(N__14579),
            .in1(N__14534),
            .in2(N__13070),
            .in3(N__14501),
            .lcout(),
            .ltout(G_7_0_m4_2_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNII9SNAB_0_LC_8_11_4.C_ON=1'b0;
    defparam beamX_RNII9SNAB_0_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam beamX_RNII9SNAB_0_LC_8_11_4.LUT_INIT=16'b0111000001111010;
    LogicCell40 beamX_RNII9SNAB_0_LC_8_11_4 (
            .in0(N__14502),
            .in1(N__14738),
            .in2(N__13067),
            .in3(N__14678),
            .lcout(G_7_0_m4_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7OTDJ61_1_LC_8_11_5.C_ON=1'b0;
    defparam beamY_RNI7OTDJ61_1_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI7OTDJ61_1_LC_8_11_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 beamY_RNI7OTDJ61_1_LC_8_11_5 (
            .in0(N__13058),
            .in1(_gnd_net_),
            .in2(N__15209),
            .in3(N__13375),
            .lcout(),
            .ltout(beamY_RNI7OTDJ61Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__font_un126_pixel_6_am_LC_8_11_6.C_ON=1'b0;
    defparam un114_pixel_6_1_5__font_un126_pixel_6_am_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__font_un126_pixel_6_am_LC_8_11_6.LUT_INIT=16'b1111100101100000;
    LogicCell40 un114_pixel_6_1_5__font_un126_pixel_6_am_LC_8_11_6 (
            .in0(N__14535),
            .in1(N__14580),
            .in2(N__13049),
            .in3(N__13274),
            .lcout(),
            .ltout(font_un126_pixel_6_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQ6MATS2_0_LC_8_11_7.C_ON=1'b0;
    defparam beamX_RNIQ6MATS2_0_LC_8_11_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIQ6MATS2_0_LC_8_11_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamX_RNIQ6MATS2_0_LC_8_11_7 (
            .in0(_gnd_net_),
            .in1(N__14503),
            .in2(N__13268),
            .in3(N__13265),
            .lcout(beamX_RNIQ6MATS2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII25UDD3_1_0_LC_8_12_0.C_ON=1'b0;
    defparam beamY_RNII25UDD3_1_0_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam beamY_RNII25UDD3_1_0_LC_8_12_0.LUT_INIT=16'b1101110100010001;
    LogicCell40 beamY_RNII25UDD3_1_0_LC_8_12_0 (
            .in0(N__13249),
            .in1(N__15127),
            .in2(_gnd_net_),
            .in3(N__14381),
            .lcout(beamY_RNII25UDD3_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m36_LC_8_12_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m36_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m36_LC_8_12_1.LUT_INIT=16'b0101010111011101;
    LogicCell40 un114_pixel_6_1_5__m36_LC_8_12_1 (
            .in0(N__15841),
            .in1(N__16054),
            .in2(_gnd_net_),
            .in3(N__15673),
            .lcout(),
            .ltout(N_37_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI05CI5A3_1_0_LC_8_12_2.C_ON=1'b0;
    defparam beamY_RNI05CI5A3_1_0_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI05CI5A3_1_0_LC_8_12_2.LUT_INIT=16'b0000001111001111;
    LogicCell40 beamY_RNI05CI5A3_1_0_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(N__15128),
            .in2(N__13226),
            .in3(N__15176),
            .lcout(),
            .ltout(beamY_RNI05CI5A3_1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJFRDMU2_1_LC_8_12_3.C_ON=1'b0;
    defparam beamY_RNIJFRDMU2_1_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIJFRDMU2_1_LC_8_12_3.LUT_INIT=16'b0000010110111011;
    LogicCell40 beamY_RNIJFRDMU2_1_LC_8_12_3 (
            .in0(N__13377),
            .in1(N__14654),
            .in2(N__13223),
            .in3(N__14937),
            .lcout(),
            .ltout(un116_pixel_7_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFHEQCT1_0_LC_8_12_4.C_ON=1'b0;
    defparam beamY_RNIFHEQCT1_0_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIFHEQCT1_0_LC_8_12_4.LUT_INIT=16'b1010110000001111;
    LogicCell40 beamY_RNIFHEQCT1_0_LC_8_12_4 (
            .in0(N__13220),
            .in1(N__13214),
            .in2(N__13208),
            .in3(N__13378),
            .lcout(beamY_RNIFHEQCT1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIA4V0NM1_0_LC_8_12_5.C_ON=1'b0;
    defparam beamY_RNIA4V0NM1_0_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIA4V0NM1_0_LC_8_12_5.LUT_INIT=16'b1000001001000010;
    LogicCell40 beamY_RNIA4V0NM1_0_LC_8_12_5 (
            .in0(N__15842),
            .in1(N__13280),
            .in2(N__15161),
            .in3(N__15674),
            .lcout(),
            .ltout(beamY_RNIA4V0NM1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUJBUM5_1_LC_8_12_6.C_ON=1'b0;
    defparam beamY_RNIUJBUM5_1_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIUJBUM5_1_LC_8_12_6.LUT_INIT=16'b0011001100011101;
    LogicCell40 beamY_RNIUJBUM5_1_LC_8_12_6 (
            .in0(N__13286),
            .in1(N__14930),
            .in2(N__13196),
            .in3(N__13376),
            .lcout(),
            .ltout(un116_pixel_7_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBHJ7AM_0_LC_8_12_7.C_ON=1'b0;
    defparam beamY_RNIBHJ7AM_0_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBHJ7AM_0_LC_8_12_7.LUT_INIT=16'b1010110000001111;
    LogicCell40 beamY_RNIBHJ7AM_0_LC_8_12_7 (
            .in0(N__14669),
            .in1(N__13400),
            .in2(N__13391),
            .in3(N__13381),
            .lcout(beamY_RNIBHJ7AMZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_8_13_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_8_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_8_13_0 (
            .in0(_gnd_net_),
            .in1(N__16583),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_8_13_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_8_13_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_8_13_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_8_13_1 (
            .in0(_gnd_net_),
            .in1(N__13304),
            .in2(N__13316),
            .in3(N__15582),
            .lcout(G_340),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_8_13_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_8_13_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_8_13_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_8_13_2 (
            .in0(_gnd_net_),
            .in1(N__13478),
            .in2(N__15657),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_8_13_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_8_13_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_8_13_3 (
            .in0(_gnd_net_),
            .in1(N__13298),
            .in2(N__13460),
            .in3(N__15583),
            .lcout(G_341),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_8_13_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_8_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_s_5_LC_8_13_4 (
            .in0(_gnd_net_),
            .in1(N__13448),
            .in2(_gnd_net_),
            .in3(N__13292),
            .lcout(un5_rowlto0),
            .ltout(un5_rowlto0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m39_LC_8_13_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m39_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m39_LC_8_13_5.LUT_INIT=16'b0010100000100000;
    LogicCell40 un114_pixel_6_1_5__m39_LC_8_13_5 (
            .in0(N__15632),
            .in1(N__16035),
            .in2(N__13289),
            .in3(N__15475),
            .lcout(un114_pixel_0_1__N_6_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ720T72_0_LC_8_13_6.C_ON=1'b0;
    defparam beamY_RNIJ720T72_0_LC_8_13_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ720T72_0_LC_8_13_6.LUT_INIT=16'b1101000110110010;
    LogicCell40 beamY_RNIJ720T72_0_LC_8_13_6 (
            .in0(N__16037),
            .in1(N__13427),
            .in2(N__15163),
            .in3(N__15848),
            .lcout(beamY_RNIJ720T72Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHD4CEK_0_LC_8_13_7.C_ON=1'b0;
    defparam beamY_RNIHD4CEK_0_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIHD4CEK_0_LC_8_13_7.LUT_INIT=16'b0011001101110111;
    LogicCell40 beamY_RNIHD4CEK_0_LC_8_13_7 (
            .in0(N__15137),
            .in1(N__16036),
            .in2(_gnd_net_),
            .in3(N__15476),
            .lcout(un116_pixel_5_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_14_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_14_0 (
            .in0(_gnd_net_),
            .in1(N__16454),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_8_14_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_8_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_8_14_1 (
            .in0(_gnd_net_),
            .in1(N__16094),
            .in2(N__13490),
            .in3(N__13472),
            .lcout(if_generate_plus_mult1_un75_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_8_14_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_8_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_8_14_2 (
            .in0(_gnd_net_),
            .in1(N__13469),
            .in2(N__16087),
            .in3(N__13451),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_8_14_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_8_14_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_8_14_3 (
            .in0(N__15587),
            .in1(N__13406),
            .in2(N__13421),
            .in3(N__13442),
            .lcout(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_8_14_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_8_14_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_s_5_LC_8_14_4 (
            .in0(_gnd_net_),
            .in1(N__13439),
            .in2(_gnd_net_),
            .in3(N__13430),
            .lcout(un5_rowlto1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m2_0_LC_8_14_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m2_0_LC_8_14_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m2_0_LC_8_14_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 un114_pixel_6_1_5__m2_0_LC_8_14_5 (
            .in0(N__15588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15467),
            .lcout(N_321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6CDEHM3_0_LC_8_14_6.C_ON=1'b0;
    defparam beamY_RNI6CDEHM3_0_LC_8_14_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI6CDEHM3_0_LC_8_14_6.LUT_INIT=16'b0101000001111111;
    LogicCell40 beamY_RNI6CDEHM3_0_LC_8_14_6 (
            .in0(N__15468),
            .in1(N__15133),
            .in2(N__16088),
            .in3(N__15589),
            .lcout(un116_pixel_2_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_8_14_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_8_14_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_8_14_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_8_14_7 (
            .in0(N__13420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16071),
            .lcout(if_generate_plus_mult1_un75_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_3_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_3_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_3_0 (
            .in0(_gnd_net_),
            .in1(N__14221),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_9_3_1.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_9_3_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_9_3_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_9_3_1 (
            .in0(_gnd_net_),
            .in1(N__13700),
            .in2(_gnd_net_),
            .in3(N__13760),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_4_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_4_0.LUT_INIT=16'b1100110000110011;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_4_0 (
            .in0(_gnd_net_),
            .in1(N__13958),
            .in2(_gnd_net_),
            .in3(N__13542),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_9_4_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_9_4_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_9_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_9_4_1 (
            .in0(_gnd_net_),
            .in1(N__14222),
            .in2(_gnd_net_),
            .in3(N__13727),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_9_4_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_9_4_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_9_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_9_4_2 (
            .in0(_gnd_net_),
            .in1(N__14226),
            .in2(N__14265),
            .in3(N__13715),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_4_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13706),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_4_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13703),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__SUM5_3_a3_LC_9_5_0.C_ON=1'b1;
    defparam un114_pixel_6_1_5__SUM5_3_a3_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__SUM5_3_a3_LC_9_5_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_6_1_5__SUM5_3_a3_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__13682),
            .in2(_gnd_net_),
            .in3(N__13615),
            .lcout(N_520),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_9_5_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_9_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__13828),
            .in2(N__13508),
            .in3(N__13493),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_9_5_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_9_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(N__13982),
            .in2(N__13816),
            .in3(N__13976),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_9_5_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_9_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_9_5_3 (
            .in0(N__13789),
            .in1(N__13829),
            .in2(N__13973),
            .in3(N__13964),
            .lcout(charx_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_9_5_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_9_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_9_5_4 (
            .in0(N__13957),
            .in1(N__13841),
            .in2(N__13817),
            .in3(N__13835),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0),
            .ltout(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_9_5_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_9_5_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_9_5_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13832),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_9_5_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_9_5_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_9_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_9_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13827),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_9_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_9_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(N__14346),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_9_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_9_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_9_6_1 (
            .in0(_gnd_net_),
            .in1(N__13802),
            .in2(N__14074),
            .in3(N__13793),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_9_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_9_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(N__13790),
            .in2(N__13778),
            .in3(N__13769),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_9_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_9_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_9_6_3 (
            .in0(N__14012),
            .in1(N__13766),
            .in2(N__14075),
            .in3(N__14060),
            .lcout(charx_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_9_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_9_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_9_6_4 (
            .in0(_gnd_net_),
            .in1(N__14057),
            .in2(_gnd_net_),
            .in3(N__14051),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_7_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_7_0 (
            .in0(_gnd_net_),
            .in1(N__15287),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_9_7_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_9_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(N__14288),
            .in2(N__13996),
            .in3(N__14048),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_9_7_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_9_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(N__14011),
            .in2(N__14045),
            .in3(N__14036),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_9_7_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_9_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_9_7_3 (
            .in0(N__16243),
            .in1(N__14033),
            .in2(N__13997),
            .in3(N__14027),
            .lcout(charx_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_9_7_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_9_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__14024),
            .in2(_gnd_net_),
            .in3(N__14018),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3),
            .ltout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_9_7_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_9_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14015),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_9_7_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_9_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14010),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_7_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_9_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_9_7_7 (
            .in0(N__14351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_9_9_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_9_9_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16664),
            .in3(N__14282),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__14270),
            .in2(N__16652),
            .in3(N__14096),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16621),
            .in3(N__14093),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14090),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__g0_10_LC_9_9_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__g0_10_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__g0_10_LC_9_9_5.LUT_INIT=16'b0110011000110011;
    LogicCell40 un114_pixel_6_1_5__g0_10_LC_9_9_5 (
            .in0(N__14536),
            .in1(N__14414),
            .in2(_gnd_net_),
            .in3(N__14581),
            .lcout(un114_pixel_6_1_5__g2_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_10_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(N__14531),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_9_10_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_9_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(N__14617),
            .in2(N__16598),
            .in3(N__14078),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPB3_LC_9_10_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPB3_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPB3_LC_9_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPB3_LC_9_10_2 (
            .in0(_gnd_net_),
            .in1(N__14636),
            .in2(N__14599),
            .in3(N__14630),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_10_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(N__14618),
            .in2(N__14627),
            .in3(N__14616),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_9_10_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_9_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_9_10_4 (
            .in0(N__14606),
            .in1(N__16622),
            .in2(N__14600),
            .in3(N__14585),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3),
            .ltout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_LC_9_10_5.C_ON=1'b0;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_LC_9_10_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_LC_9_10_5.LUT_INIT=16'b1011011111101101;
    LogicCell40 un114_pixel_6_1_5__font_un126_pixel_m_1_1_LC_9_10_5 (
            .in0(N__14532),
            .in1(N__14558),
            .in2(N__14552),
            .in3(N__14393),
            .lcout(un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_9_10_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_9_10_6.LUT_INIT=16'b1100110000110011;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(N__16577),
            .in2(_gnd_net_),
            .in3(N__16499),
            .lcout(charx_if_generate_plus_mult1_un1_sum_axb1),
            .ltout(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_1_LC_9_10_7.C_ON=1'b0;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_1_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__font_un126_pixel_m_1_1_1_LC_9_10_7.LUT_INIT=16'b0101011001010110;
    LogicCell40 un114_pixel_6_1_5__font_un126_pixel_m_1_1_1_LC_9_10_7 (
            .in0(N__14498),
            .in1(N__14413),
            .in2(N__14396),
            .in3(_gnd_net_),
            .lcout(un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_4_0_15__m15_LC_9_11_0.C_ON=1'b0;
    defparam un114_pixel_4_0_15__m15_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_4_0_15__m15_LC_9_11_0.LUT_INIT=16'b0110100001100000;
    LogicCell40 un114_pixel_4_0_15__m15_LC_9_11_0 (
            .in0(N__15680),
            .in1(N__16011),
            .in2(N__15874),
            .in3(N__15495),
            .lcout(),
            .ltout(m15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII25UDD3_0_LC_9_11_1.C_ON=1'b0;
    defparam beamY_RNII25UDD3_0_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam beamY_RNII25UDD3_0_LC_9_11_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 beamY_RNII25UDD3_0_LC_9_11_1 (
            .in0(N__15146),
            .in1(_gnd_net_),
            .in2(N__14387),
            .in3(N__14384),
            .lcout(beamY_RNII25UDD3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI4NRC8D1_0_LC_9_11_3.C_ON=1'b0;
    defparam beamY_RNI4NRC8D1_0_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI4NRC8D1_0_LC_9_11_3.LUT_INIT=16'b1101111011010100;
    LogicCell40 beamY_RNI4NRC8D1_0_LC_9_11_3 (
            .in0(N__16012),
            .in1(N__14663),
            .in2(N__15165),
            .in3(N__14724),
            .lcout(),
            .ltout(beamY_RNI4NRC8D1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNID79CMQ_1_LC_9_11_4.C_ON=1'b0;
    defparam beamY_RNID79CMQ_1_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam beamY_RNID79CMQ_1_LC_9_11_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNID79CMQ_1_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(N__14925),
            .in2(N__14687),
            .in3(N__14684),
            .lcout(N_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBKJ0H51_0_LC_9_11_5.C_ON=1'b0;
    defparam beamY_RNIBKJ0H51_0_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIBKJ0H51_0_LC_9_11_5.LUT_INIT=16'b0110001101000011;
    LogicCell40 beamY_RNIBKJ0H51_0_LC_9_11_5 (
            .in0(N__15496),
            .in1(N__15868),
            .in2(N__15164),
            .in3(N__15681),
            .lcout(),
            .ltout(un116_pixel_2_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIH01F2S_0_LC_9_11_6.C_ON=1'b0;
    defparam beamY_RNIH01F2S_0_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIH01F2S_0_LC_9_11_6.LUT_INIT=16'b0001111100010000;
    LogicCell40 beamY_RNIH01F2S_0_LC_9_11_6 (
            .in0(N__14725),
            .in1(N__15153),
            .in2(N__14672),
            .in3(N__16013),
            .lcout(beamY_RNIH01F2SZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_ns_1_5_LC_9_12_0.C_ON=1'b0;
    defparam un116_pixel_2_ns_1_5_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_ns_1_5_LC_9_12_0.LUT_INIT=16'b0111000001110011;
    LogicCell40 un116_pixel_2_ns_1_5_LC_9_12_0 (
            .in0(N__15492),
            .in1(N__15794),
            .in2(N__16085),
            .in3(N__15678),
            .lcout(un116_pixel_2_ns_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__un114_pixel_3_0_3_LC_9_12_1.C_ON=1'b0;
    defparam un114_pixel_6_1_5__un114_pixel_3_0_3_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__un114_pixel_3_0_3_LC_9_12_1.LUT_INIT=16'b0110110111101101;
    LogicCell40 un114_pixel_6_1_5__un114_pixel_3_0_3_LC_9_12_1 (
            .in0(N__15679),
            .in1(N__16066),
            .in2(N__15852),
            .in3(N__15494),
            .lcout(),
            .ltout(N_276_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII25UDD3_3_0_LC_9_12_2.C_ON=1'b0;
    defparam beamY_RNII25UDD3_3_0_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam beamY_RNII25UDD3_3_0_LC_9_12_2.LUT_INIT=16'b0000110000111111;
    LogicCell40 beamY_RNII25UDD3_3_0_LC_9_12_2 (
            .in0(_gnd_net_),
            .in1(N__15109),
            .in2(N__14657),
            .in3(N__14645),
            .lcout(beamY_RNII25UDD3_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m7_LC_9_12_3.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m7_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m7_LC_9_12_3.LUT_INIT=16'b0010100100100001;
    LogicCell40 un114_pixel_6_1_5__m7_LC_9_12_3 (
            .in0(N__15677),
            .in1(N__16061),
            .in2(N__15851),
            .in3(N__15491),
            .lcout(m7),
            .ltout(m7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNII25UDD3_2_0_LC_9_12_4.C_ON=1'b0;
    defparam beamY_RNII25UDD3_2_0_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam beamY_RNII25UDD3_2_0_LC_9_12_4.LUT_INIT=16'b0011000011111100;
    LogicCell40 beamY_RNII25UDD3_2_0_LC_9_12_4 (
            .in0(_gnd_net_),
            .in1(N__15108),
            .in2(N__14639),
            .in3(N__15193),
            .lcout(un116_pixel_3_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_LC_9_12_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_LC_9_12_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 un114_pixel_1_0_3__g0_LC_9_12_5 (
            .in0(N__15798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15493),
            .lcout(N_302_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITQPUS72_0_LC_9_12_6.C_ON=1'b0;
    defparam beamY_RNITQPUS72_0_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam beamY_RNITQPUS72_0_LC_9_12_6.LUT_INIT=16'b1110000010010101;
    LogicCell40 beamY_RNITQPUS72_0_LC_9_12_6 (
            .in0(N__16065),
            .in1(N__15182),
            .in2(N__15160),
            .in3(N__15793),
            .lcout(),
            .ltout(beamY_RNITQPUS72Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6B7UAL1_1_LC_9_12_7.C_ON=1'b0;
    defparam beamY_RNI6B7UAL1_1_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI6B7UAL1_1_LC_9_12_7.LUT_INIT=16'b1010000011110101;
    LogicCell40 beamY_RNI6B7UAL1_1_LC_9_12_7 (
            .in0(N__14924),
            .in1(_gnd_net_),
            .in2(N__15218),
            .in3(N__15215),
            .lcout(beamY_RNI6B7UAL1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m31_LC_9_13_0.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m31_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m31_LC_9_13_0.LUT_INIT=16'b0011100000000011;
    LogicCell40 un114_pixel_6_1_5__m31_LC_9_13_0 (
            .in0(N__15497),
            .in1(N__15624),
            .in2(N__15849),
            .in3(N__16056),
            .lcout(m31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_4_1_0_LC_9_13_1.C_ON=1'b0;
    defparam un116_pixel_4_1_0_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam un116_pixel_4_1_0_LC_9_13_1.LUT_INIT=16'b0000111110101111;
    LogicCell40 un116_pixel_4_1_0_LC_9_13_1 (
            .in0(N__16057),
            .in1(_gnd_net_),
            .in2(N__15675),
            .in3(N__15498),
            .lcout(un116_pixel_4_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_6_1_5__m38_LC_9_13_2.C_ON=1'b0;
    defparam un114_pixel_6_1_5__m38_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_6_1_5__m38_LC_9_13_2.LUT_INIT=16'b0000101000000010;
    LogicCell40 un114_pixel_6_1_5__m38_LC_9_13_2 (
            .in0(N__15500),
            .in1(N__15631),
            .in2(N__15850),
            .in3(N__16060),
            .lcout(m38),
            .ltout(m38_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPG8ISM3_1_LC_9_13_3.C_ON=1'b0;
    defparam beamY_RNIPG8ISM3_1_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIPG8ISM3_1_LC_9_13_3.LUT_INIT=16'b0011101100011001;
    LogicCell40 beamY_RNIPG8ISM3_1_LC_9_13_3 (
            .in0(N__14923),
            .in1(N__15138),
            .in2(N__14942),
            .in3(N__15789),
            .lcout(),
            .ltout(un116_pixel_6_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICKDGA43_1_LC_9_13_4.C_ON=1'b0;
    defparam beamY_RNICKDGA43_1_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam beamY_RNICKDGA43_1_LC_9_13_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 beamY_RNICKDGA43_1_LC_9_13_4 (
            .in0(N__14938),
            .in1(N__14693),
            .in2(N__14741),
            .in3(N__15347),
            .lcout(N_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_bm_1_LC_9_13_5.C_ON=1'b0;
    defparam un116_pixel_2_bm_1_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_bm_1_LC_9_13_5.LUT_INIT=16'b1101110111001100;
    LogicCell40 un116_pixel_2_bm_1_LC_9_13_5 (
            .in0(N__16058),
            .in1(N__14722),
            .in2(_gnd_net_),
            .in3(N__15788),
            .lcout(un116_pixel_2_bmZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_rowlto2_sbtinv_LC_9_13_6.C_ON=1'b0;
    defparam un5_rowlto2_sbtinv_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam un5_rowlto2_sbtinv_LC_9_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_rowlto2_sbtinv_LC_9_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16055),
            .lcout(un5_rowlto2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_am_1_LC_9_13_7.C_ON=1'b0;
    defparam un116_pixel_2_am_1_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_am_1_LC_9_13_7.LUT_INIT=16'b1001010010110100;
    LogicCell40 un116_pixel_2_am_1_LC_9_13_7 (
            .in0(N__16059),
            .in1(N__15787),
            .in2(N__15676),
            .in3(N__15499),
            .lcout(un116_pixel_2_amZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(N__16136),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__15239),
            .in2(N__15341),
            .in3(N__15326),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__15323),
            .in2(N__16253),
            .in3(N__15311),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_11_5_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_11_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_11_5_3 (
            .in0(N__16216),
            .in1(N__16267),
            .in2(N__16229),
            .in3(N__15308),
            .lcout(charx_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_11_5_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_11_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(N__15305),
            .in2(_gnd_net_),
            .in3(N__15293),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7),
            .ltout(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_11_5_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_11_5_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_11_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15290),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_11_5_6.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_11_5_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_11_5_6 (
            .in0(N__15284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_11_5_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_11_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_11_5_7 (
            .in0(_gnd_net_),
            .in1(N__16268),
            .in2(_gnd_net_),
            .in3(N__16249),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_11_6_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_11_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__16326),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_11_6_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_11_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__16100),
            .in2(N__16186),
            .in3(N__16220),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_11_6_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_11_6_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_11_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(N__16217),
            .in2(N__16205),
            .in3(N__16196),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_11_6_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_11_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_11_6_3 (
            .in0(N__16399),
            .in1(N__16193),
            .in2(N__16187),
            .in3(N__16172),
            .lcout(charx_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_11_6_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_11_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(N__16169),
            .in2(_gnd_net_),
            .in3(N__16163),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0),
            .ltout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_11_6_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_11_6_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_11_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16160),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_11_6_7.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_11_6_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_11_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_11_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16155),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_11_7_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_11_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_11_7_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_11_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__16295),
            .in2(N__16369),
            .in3(N__16403),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_11_7_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_11_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__16400),
            .in2(N__16388),
            .in3(N__16379),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_11_7_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_11_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_11_7_3 (
            .in0(N__16708),
            .in1(N__16376),
            .in2(N__16370),
            .in3(N__16355),
            .lcout(charx_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_11_7_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_11_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_11_7_4 (
            .in0(_gnd_net_),
            .in1(N__16352),
            .in2(_gnd_net_),
            .in3(N__16346),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_11_7_7.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_11_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_11_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16327),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_8_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(N__16562),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_11_8_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_11_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(N__16289),
            .in2(N__16690),
            .in3(N__16280),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_11_8_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_11_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__16277),
            .in2(N__16709),
            .in3(N__16271),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_11_8_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_11_8_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_11_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(N__16715),
            .in2(N__16691),
            .in3(N__16704),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_11_8_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_11_8_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_11_8_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_11_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16676),
            .in3(N__16667),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_11_9_0.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_11_9_0.LUT_INIT=16'b1011010000001111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_11_9_0 (
            .in0(N__16579),
            .in1(N__16514),
            .in2(N__16639),
            .in3(N__16486),
            .lcout(charx_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_11_9_1.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_11_9_1.LUT_INIT=16'b1101000000101111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_11_9_1 (
            .in0(N__16515),
            .in1(N__16581),
            .in2(N__16495),
            .in3(N__16635),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_11_9_2.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_11_9_2.LUT_INIT=16'b0100101111110000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_11_9_2 (
            .in0(N__16580),
            .in1(N__16516),
            .in2(N__16640),
            .in3(N__16490),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_11_9_3.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_11_9_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_11_9_3.LUT_INIT=16'b0000111110100101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_11_9_3 (
            .in0(N__16491),
            .in1(_gnd_net_),
            .in2(N__16520),
            .in3(N__16582),
            .lcout(charx_i_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_11_9_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_11_9_4.LUT_INIT=16'b1001100111001100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_11_9_4 (
            .in0(N__16578),
            .in1(N__16513),
            .in2(_gnd_net_),
            .in3(N__16485),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
