-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 16:41:40

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic;
    Clock12MHz : in std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__4026\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1877\ : std_logic;
signal \N__1874\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1856\ : std_logic;
signal \VGAClock.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\ : std_logic;
signal \y_RNIA5P7Z0Z_9\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0\ : std_logic;
signal \Pixel_RNOZ0Z_8\ : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \N_11\ : std_logic;
signal \un12_0_1_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2\ : std_logic;
signal \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5\ : std_logic;
signal un2_y_if_generate_plus_mult1_un47_sum_axb_7 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal \y_RNI94P7Z0Z_8\ : std_logic;
signal un2_y_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \G_7_i_a4_0_0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal un4_y_cry_1 : std_logic;
signal un4_y_cry_2 : std_logic;
signal un4_y_cry_3 : std_logic;
signal un4_y_cry_4 : std_logic;
signal un4_y_cry_5 : std_logic;
signal un4_y_cry_6 : std_logic;
signal un4_y_cry_7 : std_logic;
signal un4_y_cry_8 : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \bfn_4_1_0_\ : std_logic;
signal un16_x_cry_1 : std_logic;
signal un16_x_cry_2 : std_logic;
signal un16_x_cry_3 : std_logic;
signal un16_x_cry_4 : std_logic;
signal un16_x_cry_5 : std_logic;
signal un16_x_cry_6 : std_logic;
signal un16_x_cry_7 : std_logic;
signal un16_x_cry_8 : std_logic;
signal \bfn_4_2_0_\ : std_logic;
signal un8_xlt9_0 : std_logic;
signal \Pixel_0_sqmuxa_0_cascade_\ : std_logic;
signal \Pixel_0_sqmuxa_1\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\ : std_logic;
signal \Pixel_RNOZ0Z_5\ : std_logic;
signal un2_x_27 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\ : std_logic;
signal un13lt10 : std_logic;
signal \un1_ylto9_5_cascade_\ : std_logic;
signal \un4_y_cry_2_THRU_CO\ : std_logic;
signal \yZ0Z_5\ : std_logic;
signal \yZ0Z_6\ : std_logic;
signal \yZ0Z_1\ : std_logic;
signal un1_ylto9_4 : std_logic;
signal \un4_y_cry_1_THRU_CO\ : std_logic;
signal \yZ0Z_4\ : std_logic;
signal \yZ0Z_3\ : std_logic;
signal \yZ0Z_2\ : std_logic;
signal \yZ0Z_9\ : std_logic;
signal \yZ0Z_8\ : std_logic;
signal y_12_5 : std_logic;
signal \y_12_6_cascade_\ : std_logic;
signal \yZ0Z_7\ : std_logic;
signal y_12_8 : std_logic;
signal \y_12_8_cascade_\ : std_logic;
signal \yZ0Z_0\ : std_logic;
signal \un11_x_4_0_cascade_\ : std_logic;
signal \x_RNID8R22Z0Z_9\ : std_logic;
signal \xZ0Z_2\ : std_logic;
signal \xZ0Z_1\ : std_logic;
signal \xZ0Z_3\ : std_logic;
signal \xZ0Z_0\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal un11_x_3_0 : std_logic;
signal \xZ0Z_4\ : std_logic;
signal un4_xlt9 : std_logic;
signal \xZ0Z_9\ : std_logic;
signal \HSync_c\ : std_logic;
signal \xZ0Z_8\ : std_logic;
signal un1_xlto9_0 : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un40_sum_i : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_i : std_logic;
signal un1_y : std_logic;
signal \VSync_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \xZ0Z_5\ : std_logic;
signal un11_x_4 : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_i : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\ : std_logic;
signal \xZ0Z_7\ : std_logic;
signal \xZ0Z_6\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un2_x_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\ : std_logic;
signal un2_x_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\ : std_logic;
signal \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\ : std_logic;
signal un2_x_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \VGAClock.PixelClock_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1001010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \VGAClock.PixelClock\,
            REFERENCECLK => \N__1865\,
            RESETB => \N__3308\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \VGAClock.PixelClock_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4026\,
            DIN => \N__4025\,
            DOUT => \N__4024\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4026\,
            PADOUT => \N__4025\,
            PADIN => \N__4024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3731\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4017\,
            DIN => \N__4016\,
            DOUT => \N__4015\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4017\,
            PADOUT => \N__4016\,
            PADIN => \N__4015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3380\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4008\,
            DIN => \N__4007\,
            DOUT => \N__4006\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4008\,
            PADOUT => \N__4007\,
            PADIN => \N__4006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2132\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3999\,
            DIN => \N__3998\,
            DOUT => \N__3997\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3999\,
            PADOUT => \N__3998\,
            PADIN => \N__3997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__873\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3973\
        );

    \I__872\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3973\
        );

    \I__871\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3969\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__3973\,
            I => \N__3965\
        );

    \I__869\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3962\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__3969\,
            I => \N__3959\
        );

    \I__867\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3956\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__3965\,
            I => \N__3953\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__3962\,
            I => \xZ0Z_7\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__3959\,
            I => \xZ0Z_7\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__3956\,
            I => \xZ0Z_7\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__3953\,
            I => \xZ0Z_7\
        );

    \I__861\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3940\
        );

    \I__860\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3937\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__3940\,
            I => \N__3927\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__3937\,
            I => \N__3927\
        );

    \I__857\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3924\
        );

    \I__856\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3921\
        );

    \I__855\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3916\
        );

    \I__854\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3916\
        );

    \I__853\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3913\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__3927\,
            I => \N__3910\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__3924\,
            I => \xZ0Z_6\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__3921\,
            I => \xZ0Z_6\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__3916\,
            I => \xZ0Z_6\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__3913\,
            I => \xZ0Z_6\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__3910\,
            I => \xZ0Z_6\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__845\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__3893\,
            I => un2_x_if_generate_plus_mult1_un54_sum_i
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__842\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__3884\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\
        );

    \I__840\ : InMux
    port map (
            O => \N__3881\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__839\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3874\
        );

    \I__838\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3871\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__3874\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__3871\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__834\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__3860\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__831\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__3851\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\
        );

    \I__829\ : InMux
    port map (
            O => \N__3848\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__828\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3839\
        );

    \I__827\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3839\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__3839\,
            I => un2_x_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__824\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__3830\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\
        );

    \I__822\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3824\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__3824\,
            I => un2_x_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__820\ : InMux
    port map (
            O => \N__3821\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__819\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3815\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__3815\,
            I => un2_x_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__817\ : InMux
    port map (
            O => \N__3812\,
            I => un2_x_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__816\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3805\
        );

    \I__815\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3802\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__3805\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3802\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__3797\,
            I => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\
        );

    \I__811\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3788\
        );

    \I__810\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3788\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__3788\,
            I => un2_x_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__808\ : InMux
    port map (
            O => \N__3785\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__807\ : InMux
    port map (
            O => \N__3782\,
            I => \N__3778\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__3781\,
            I => \N__3775\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3771\
        );

    \I__804\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3766\
        );

    \I__803\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3766\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__3771\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__3766\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__799\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3755\,
            I => un2_x_if_generate_plus_mult1_un61_sum_i
        );

    \I__797\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3749\,
            I => \N__3745\
        );

    \I__795\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3742\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__3745\,
            I => \N__3739\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3736\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__3739\,
            I => un1_y
        );

    \I__791\ : Odrv4
    port map (
            O => \N__3736\,
            I => un1_y
        );

    \I__790\ : IoInMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__788\ : IoSpan4Mux
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__3722\,
            I => \VSync_c\
        );

    \I__786\ : ClkMux
    port map (
            O => \N__3719\,
            I => \N__3692\
        );

    \I__785\ : ClkMux
    port map (
            O => \N__3718\,
            I => \N__3692\
        );

    \I__784\ : ClkMux
    port map (
            O => \N__3717\,
            I => \N__3692\
        );

    \I__783\ : ClkMux
    port map (
            O => \N__3716\,
            I => \N__3692\
        );

    \I__782\ : ClkMux
    port map (
            O => \N__3715\,
            I => \N__3692\
        );

    \I__781\ : ClkMux
    port map (
            O => \N__3714\,
            I => \N__3692\
        );

    \I__780\ : ClkMux
    port map (
            O => \N__3713\,
            I => \N__3692\
        );

    \I__779\ : ClkMux
    port map (
            O => \N__3712\,
            I => \N__3692\
        );

    \I__778\ : ClkMux
    port map (
            O => \N__3711\,
            I => \N__3692\
        );

    \I__777\ : GlobalMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__776\ : gio2CtrlBuf
    port map (
            O => \N__3689\,
            I => \PixelClock_g\
        );

    \I__775\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3681\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__3685\,
            I => \N__3677\
        );

    \I__773\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3672\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3681\,
            I => \N__3669\
        );

    \I__771\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3666\
        );

    \I__770\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3663\
        );

    \I__769\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3660\
        );

    \I__768\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3657\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3672\,
            I => \N__3652\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__3669\,
            I => \N__3652\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3666\,
            I => \N__3649\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3663\,
            I => \xZ0Z_5\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3660\,
            I => \xZ0Z_5\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3657\,
            I => \xZ0Z_5\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__3652\,
            I => \xZ0Z_5\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3649\,
            I => \xZ0Z_5\
        );

    \I__759\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3635\,
            I => \N__3631\
        );

    \I__757\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3628\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__3631\,
            I => un11_x_4
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3628\,
            I => un11_x_4
        );

    \I__754\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3620\,
            I => un2_x_if_generate_plus_mult1_un47_sum_i
        );

    \I__752\ : InMux
    port map (
            O => \N__3617\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__751\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3610\
        );

    \I__750\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3607\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3610\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3607\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__746\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3596\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\
        );

    \I__744\ : InMux
    port map (
            O => \N__3593\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__3590\,
            I => \N__3586\
        );

    \I__742\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3583\
        );

    \I__741\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3580\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3583\,
            I => un2_x_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3580\,
            I => un2_x_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__737\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3569\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\
        );

    \I__735\ : InMux
    port map (
            O => \N__3566\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__734\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3560\,
            I => un2_x_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__732\ : InMux
    port map (
            O => \N__3557\,
            I => un2_x_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__3554\,
            I => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\
        );

    \I__730\ : InMux
    port map (
            O => \N__3551\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__729\ : InMux
    port map (
            O => \N__3548\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3545\,
            I => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3542\,
            I => \N__3539\
        );

    \I__726\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3533\
        );

    \I__725\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3533\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3533\,
            I => \N__3529\
        );

    \I__723\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__3529\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3526\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__720\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3518\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3518\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\
        );

    \I__718\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3512\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\
        );

    \I__716\ : InMux
    port map (
            O => \N__3509\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__714\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3500\,
            I => \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\
        );

    \I__712\ : InMux
    port map (
            O => \N__3497\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__711\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3491\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3491\,
            I => un2_x_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__709\ : InMux
    port map (
            O => \N__3488\,
            I => un2_x_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__708\ : InMux
    port map (
            O => \N__3485\,
            I => un2_x_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__3482\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\
        );

    \I__706\ : InMux
    port map (
            O => \N__3479\,
            I => \N__3475\
        );

    \I__705\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3472\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3475\,
            I => un11_x_3_0
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3472\,
            I => un11_x_3_0
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__701\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3451\
        );

    \I__700\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3451\
        );

    \I__699\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3451\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3461\,
            I => \N__3448\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__3460\,
            I => \N__3445\
        );

    \I__696\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3442\
        );

    \I__695\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3439\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3451\,
            I => \N__3436\
        );

    \I__693\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3433\
        );

    \I__692\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3430\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3442\,
            I => \xZ0Z_4\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3439\,
            I => \xZ0Z_4\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__3436\,
            I => \xZ0Z_4\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3433\,
            I => \xZ0Z_4\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3430\,
            I => \xZ0Z_4\
        );

    \I__686\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3416\,
            I => un4_xlt9
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3413\,
            I => \N__3408\
        );

    \I__683\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3402\
        );

    \I__682\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3399\
        );

    \I__681\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3396\
        );

    \I__680\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3389\
        );

    \I__679\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3389\
        );

    \I__678\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3389\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3402\,
            I => \xZ0Z_9\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3399\,
            I => \xZ0Z_9\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3396\,
            I => \xZ0Z_9\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3389\,
            I => \xZ0Z_9\
        );

    \I__673\ : IoInMux
    port map (
            O => \N__3380\,
            I => \N__3377\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__671\ : Span4Mux_s0_v
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__670\ : Span4Mux_h
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__3368\,
            I => \HSync_c\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__667\ : InMux
    port map (
            O => \N__3362\,
            I => \N__3355\
        );

    \I__666\ : InMux
    port map (
            O => \N__3361\,
            I => \N__3352\
        );

    \I__665\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3349\
        );

    \I__664\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3346\
        );

    \I__663\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3343\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3340\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3352\,
            I => \xZ0Z_8\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3349\,
            I => \xZ0Z_8\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3346\,
            I => \xZ0Z_8\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3343\,
            I => \xZ0Z_8\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__3340\,
            I => \xZ0Z_8\
        );

    \I__656\ : InMux
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3326\,
            I => un1_xlto9_0
        );

    \I__654\ : InMux
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3320\,
            I => un2_x_if_generate_plus_mult1_un40_sum_i
        );

    \I__652\ : InMux
    port map (
            O => \N__3317\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__651\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3311\,
            I => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\
        );

    \I__649\ : IoInMux
    port map (
            O => \N__3308\,
            I => \N__3302\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3307\,
            I => \N__3299\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__3306\,
            I => \N__3295\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__3305\,
            I => \N__3289\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3302\,
            I => \N__3286\
        );

    \I__644\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3279\
        );

    \I__643\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3279\
        );

    \I__642\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3279\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__3294\,
            I => \N__3276\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \N__3273\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3270\
        );

    \I__638\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3267\
        );

    \I__637\ : Span4Mux_s0_v
    port map (
            O => \N__3286\,
            I => \N__3264\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3279\,
            I => \N__3261\
        );

    \I__635\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3258\
        );

    \I__634\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3253\
        );

    \I__633\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3253\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3267\,
            I => \N__3250\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__3264\,
            I => \N__3241\
        );

    \I__630\ : Span4Mux_s1_h
    port map (
            O => \N__3261\,
            I => \N__3241\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3258\,
            I => \N__3241\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3253\,
            I => \N__3241\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__3250\,
            I => \CONSTANT_ONE_NET\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3241\,
            I => \CONSTANT_ONE_NET\
        );

    \I__625\ : InMux
    port map (
            O => \N__3236\,
            I => un2_x_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__624\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__623\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3224\
        );

    \I__622\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3221\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3230\,
            I => \N__3218\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3227\,
            I => \N__3211\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3224\,
            I => \N__3211\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3208\
        );

    \I__617\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3203\
        );

    \I__616\ : InMux
    port map (
            O => \N__3217\,
            I => \N__3203\
        );

    \I__615\ : InMux
    port map (
            O => \N__3216\,
            I => \N__3200\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__3211\,
            I => \N__3197\
        );

    \I__613\ : Odrv12
    port map (
            O => \N__3208\,
            I => \yZ0Z_3\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3203\,
            I => \yZ0Z_3\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3200\,
            I => \yZ0Z_3\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__3197\,
            I => \yZ0Z_3\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__608\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3179\
        );

    \I__607\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3175\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3183\,
            I => \N__3171\
        );

    \I__605\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3167\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3179\,
            I => \N__3164\
        );

    \I__603\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3161\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3175\,
            I => \N__3158\
        );

    \I__601\ : InMux
    port map (
            O => \N__3174\,
            I => \N__3153\
        );

    \I__600\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3153\
        );

    \I__599\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3150\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3167\,
            I => \N__3143\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__3164\,
            I => \N__3143\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3161\,
            I => \N__3143\
        );

    \I__595\ : Span4Mux_s3_h
    port map (
            O => \N__3158\,
            I => \N__3140\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3153\,
            I => \yZ0Z_2\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3150\,
            I => \yZ0Z_2\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__3143\,
            I => \yZ0Z_2\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__3140\,
            I => \yZ0Z_2\
        );

    \I__590\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3124\
        );

    \I__589\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3129\,
            I => \N__3120\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3124\,
            I => \N__3117\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__3123\,
            I => \N__3113\
        );

    \I__585\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3110\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__3117\,
            I => \N__3107\
        );

    \I__583\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3102\
        );

    \I__582\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3102\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3110\,
            I => \yZ0Z_9\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__3107\,
            I => \yZ0Z_9\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3102\,
            I => \yZ0Z_9\
        );

    \I__578\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3088\
        );

    \I__577\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3088\
        );

    \I__576\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3083\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3088\,
            I => \N__3080\
        );

    \I__574\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3077\
        );

    \I__573\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3074\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3083\,
            I => \yZ0Z_8\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__3080\,
            I => \yZ0Z_8\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3077\,
            I => \yZ0Z_8\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3074\,
            I => \yZ0Z_8\
        );

    \I__568\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3062\,
            I => y_12_5
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3059\,
            I => \y_12_6_cascade_\
        );

    \I__565\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3052\
        );

    \I__564\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3049\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3045\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3049\,
            I => \N__3040\
        );

    \I__561\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3037\
        );

    \I__560\ : Span4Mux_h
    port map (
            O => \N__3045\,
            I => \N__3034\
        );

    \I__559\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3029\
        );

    \I__558\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3029\
        );

    \I__557\ : Odrv4
    port map (
            O => \N__3040\,
            I => \yZ0Z_7\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3037\,
            I => \yZ0Z_7\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__3034\,
            I => \yZ0Z_7\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3029\,
            I => \yZ0Z_7\
        );

    \I__553\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3017\,
            I => \N__3012\
        );

    \I__551\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3007\
        );

    \I__550\ : InMux
    port map (
            O => \N__3015\,
            I => \N__3007\
        );

    \I__549\ : Span4Mux_s3_h
    port map (
            O => \N__3012\,
            I => \N__3004\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3007\,
            I => y_12_8
        );

    \I__547\ : Odrv4
    port map (
            O => \N__3004\,
            I => y_12_8
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__2999\,
            I => \y_12_8_cascade_\
        );

    \I__545\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2992\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__2995\,
            I => \N__2987\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2984\
        );

    \I__542\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2977\
        );

    \I__541\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2977\
        );

    \I__540\ : InMux
    port map (
            O => \N__2987\,
            I => \N__2977\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__2984\,
            I => \yZ0Z_0\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__2977\,
            I => \yZ0Z_0\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__2972\,
            I => \un11_x_4_0_cascade_\
        );

    \I__536\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2959\
        );

    \I__535\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2959\
        );

    \I__534\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2959\
        );

    \I__533\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2950\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2959\,
            I => \N__2947\
        );

    \I__531\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2942\
        );

    \I__530\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2942\
        );

    \I__529\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2933\
        );

    \I__528\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2933\
        );

    \I__527\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2933\
        );

    \I__526\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2933\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2930\
        );

    \I__524\ : Sp12to4
    port map (
            O => \N__2947\,
            I => \N__2922\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__2942\,
            I => \N__2922\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2933\,
            I => \N__2919\
        );

    \I__521\ : Span4Mux_h
    port map (
            O => \N__2930\,
            I => \N__2916\
        );

    \I__520\ : InMux
    port map (
            O => \N__2929\,
            I => \N__2913\
        );

    \I__519\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2910\
        );

    \I__518\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2907\
        );

    \I__517\ : Span12Mux_s4_h
    port map (
            O => \N__2922\,
            I => \N__2904\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__2919\,
            I => \N__2899\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__2916\,
            I => \N__2899\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2913\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2910\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2907\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__511\ : Odrv12
    port map (
            O => \N__2904\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__510\ : Odrv4
    port map (
            O => \N__2899\,
            I => \x_RNID8R22Z0Z_9\
        );

    \I__509\ : InMux
    port map (
            O => \N__2888\,
            I => \N__2884\
        );

    \I__508\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2881\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2884\,
            I => \xZ0Z_2\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2881\,
            I => \xZ0Z_2\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__504\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2868\
        );

    \I__503\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2863\
        );

    \I__502\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2863\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2868\,
            I => \xZ0Z_1\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2863\,
            I => \xZ0Z_1\
        );

    \I__499\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2854\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__2857\,
            I => \N__2850\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2854\,
            I => \N__2847\
        );

    \I__496\ : InMux
    port map (
            O => \N__2853\,
            I => \N__2844\
        );

    \I__495\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2841\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__2847\,
            I => \xZ0Z_3\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2844\,
            I => \xZ0Z_3\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2841\,
            I => \xZ0Z_3\
        );

    \I__491\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2828\
        );

    \I__490\ : InMux
    port map (
            O => \N__2833\,
            I => \N__2821\
        );

    \I__489\ : InMux
    port map (
            O => \N__2832\,
            I => \N__2821\
        );

    \I__488\ : InMux
    port map (
            O => \N__2831\,
            I => \N__2821\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2828\,
            I => \xZ0Z_0\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2821\,
            I => \xZ0Z_0\
        );

    \I__485\ : InMux
    port map (
            O => \N__2816\,
            I => \N__2810\
        );

    \I__484\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2810\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2810\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\
        );

    \I__482\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2804\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\
        );

    \I__480\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__2795\,
            I => un13lt10
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__2792\,
            I => \un1_ylto9_5_cascade_\
        );

    \I__476\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__474\ : Odrv12
    port map (
            O => \N__2783\,
            I => \un4_y_cry_2_THRU_CO\
        );

    \I__473\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2776\
        );

    \I__472\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2770\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2776\,
            I => \N__2767\
        );

    \I__470\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2762\
        );

    \I__469\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2762\
        );

    \I__468\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2759\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2770\,
            I => \N__2756\
        );

    \I__466\ : Span4Mux_h
    port map (
            O => \N__2767\,
            I => \N__2753\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2762\,
            I => \N__2750\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2759\,
            I => \yZ0Z_5\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__2756\,
            I => \yZ0Z_5\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__2753\,
            I => \yZ0Z_5\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__2750\,
            I => \yZ0Z_5\
        );

    \I__460\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2737\
        );

    \I__459\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2731\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2737\,
            I => \N__2728\
        );

    \I__457\ : InMux
    port map (
            O => \N__2736\,
            I => \N__2723\
        );

    \I__456\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2723\
        );

    \I__455\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2720\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2731\,
            I => \N__2717\
        );

    \I__453\ : Span4Mux_h
    port map (
            O => \N__2728\,
            I => \N__2714\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2723\,
            I => \N__2711\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2720\,
            I => \yZ0Z_6\
        );

    \I__450\ : Odrv4
    port map (
            O => \N__2717\,
            I => \yZ0Z_6\
        );

    \I__449\ : Odrv4
    port map (
            O => \N__2714\,
            I => \yZ0Z_6\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2711\,
            I => \yZ0Z_6\
        );

    \I__447\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2698\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__2701\,
            I => \N__2695\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2698\,
            I => \N__2692\
        );

    \I__444\ : InMux
    port map (
            O => \N__2695\,
            I => \N__2688\
        );

    \I__443\ : Span4Mux_s3_h
    port map (
            O => \N__2692\,
            I => \N__2683\
        );

    \I__442\ : InMux
    port map (
            O => \N__2691\,
            I => \N__2680\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2688\,
            I => \N__2677\
        );

    \I__440\ : InMux
    port map (
            O => \N__2687\,
            I => \N__2672\
        );

    \I__439\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2672\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__2683\,
            I => \yZ0Z_1\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2680\,
            I => \yZ0Z_1\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__2677\,
            I => \yZ0Z_1\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2672\,
            I => \yZ0Z_1\
        );

    \I__434\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2660\,
            I => un1_ylto9_4
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__2657\,
            I => \N__2654\
        );

    \I__431\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2651\,
            I => \N__2648\
        );

    \I__429\ : Odrv4
    port map (
            O => \N__2648\,
            I => \un4_y_cry_1_THRU_CO\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__2645\,
            I => \N__2642\
        );

    \I__427\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2636\
        );

    \I__426\ : InMux
    port map (
            O => \N__2641\,
            I => \N__2633\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__2640\,
            I => \N__2630\
        );

    \I__424\ : InMux
    port map (
            O => \N__2639\,
            I => \N__2626\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2623\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2633\,
            I => \N__2620\
        );

    \I__421\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2617\
        );

    \I__420\ : InMux
    port map (
            O => \N__2629\,
            I => \N__2614\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2626\,
            I => \N__2611\
        );

    \I__418\ : Span4Mux_h
    port map (
            O => \N__2623\,
            I => \N__2608\
        );

    \I__417\ : Span4Mux_s1_h
    port map (
            O => \N__2620\,
            I => \N__2603\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2617\,
            I => \N__2603\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2614\,
            I => \yZ0Z_4\
        );

    \I__414\ : Odrv4
    port map (
            O => \N__2611\,
            I => \yZ0Z_4\
        );

    \I__413\ : Odrv4
    port map (
            O => \N__2608\,
            I => \yZ0Z_4\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__2603\,
            I => \yZ0Z_4\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__2594\,
            I => \Pixel_0_sqmuxa_0_cascade_\
        );

    \I__410\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__408\ : Span4Mux_s3_h
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__2582\,
            I => \Pixel_0_sqmuxa_1\
        );

    \I__406\ : InMux
    port map (
            O => \N__2579\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__405\ : InMux
    port map (
            O => \N__2576\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__404\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2567\
        );

    \I__403\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2567\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2567\,
            I => un2_x_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__401\ : InMux
    port map (
            O => \N__2564\,
            I => un2_x_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__2561\,
            I => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\
        );

    \I__399\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2555\,
            I => \Pixel_RNOZ0Z_5\
        );

    \I__397\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__2546\,
            I => un2_x_27
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__393\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2537\,
            I => un2_x_if_generate_plus_mult1_un68_sum_i
        );

    \I__391\ : InMux
    port map (
            O => \N__2534\,
            I => un16_x_cry_1
        );

    \I__390\ : InMux
    port map (
            O => \N__2531\,
            I => un16_x_cry_2
        );

    \I__389\ : InMux
    port map (
            O => \N__2528\,
            I => un16_x_cry_3
        );

    \I__388\ : InMux
    port map (
            O => \N__2525\,
            I => un16_x_cry_4
        );

    \I__387\ : InMux
    port map (
            O => \N__2522\,
            I => un16_x_cry_5
        );

    \I__386\ : InMux
    port map (
            O => \N__2519\,
            I => un16_x_cry_6
        );

    \I__385\ : InMux
    port map (
            O => \N__2516\,
            I => un16_x_cry_7
        );

    \I__384\ : InMux
    port map (
            O => \N__2513\,
            I => \bfn_4_2_0_\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__382\ : InMux
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2504\,
            I => un8_xlt9_0
        );

    \I__380\ : InMux
    port map (
            O => \N__2501\,
            I => un4_y_cry_1
        );

    \I__379\ : InMux
    port map (
            O => \N__2498\,
            I => un4_y_cry_2
        );

    \I__378\ : InMux
    port map (
            O => \N__2495\,
            I => un4_y_cry_3
        );

    \I__377\ : InMux
    port map (
            O => \N__2492\,
            I => un4_y_cry_4
        );

    \I__376\ : InMux
    port map (
            O => \N__2489\,
            I => un4_y_cry_5
        );

    \I__375\ : InMux
    port map (
            O => \N__2486\,
            I => un4_y_cry_6
        );

    \I__374\ : InMux
    port map (
            O => \N__2483\,
            I => un4_y_cry_7
        );

    \I__373\ : InMux
    port map (
            O => \N__2480\,
            I => \bfn_2_7_0_\
        );

    \I__372\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2474\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2474\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0\
        );

    \I__370\ : InMux
    port map (
            O => \N__2471\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__369\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2465\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2465\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__2462\,
            I => \N__2459\
        );

    \I__366\ : InMux
    port map (
            O => \N__2459\,
            I => \N__2456\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2456\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0\
        );

    \I__364\ : InMux
    port map (
            O => \N__2453\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__363\ : InMux
    port map (
            O => \N__2450\,
            I => \N__2447\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2447\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\
        );

    \I__361\ : InMux
    port map (
            O => \N__2444\,
            I => \N__2441\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2441\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0\
        );

    \I__359\ : InMux
    port map (
            O => \N__2438\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__2435\,
            I => \N__2431\
        );

    \I__357\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2422\
        );

    \I__356\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2422\
        );

    \I__355\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2422\
        );

    \I__354\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2419\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2422\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2419\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0\
        );

    \I__351\ : InMux
    port map (
            O => \N__2414\,
            I => \N__2409\
        );

    \I__350\ : InMux
    port map (
            O => \N__2413\,
            I => \N__2406\
        );

    \I__349\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2403\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2409\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2406\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2403\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__2396\,
            I => \N__2393\
        );

    \I__344\ : InMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2390\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5\
        );

    \I__342\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2384\,
            I => un2_y_if_generate_plus_mult1_un47_sum_axb_7
        );

    \I__340\ : InMux
    port map (
            O => \N__2381\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__339\ : InMux
    port map (
            O => \N__2378\,
            I => un2_y_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2375\,
            I => \N__2372\
        );

    \I__337\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2369\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2369\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__335\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2363\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2363\,
            I => \y_RNI94P7Z0Z_8\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__332\ : InMux
    port map (
            O => \N__2357\,
            I => \N__2354\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2354\,
            I => un2_y_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__330\ : InMux
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__328\ : Odrv12
    port map (
            O => \N__2345\,
            I => \G_7_i_a4_0_0\
        );

    \I__327\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2339\,
            I => \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21\
        );

    \I__325\ : InMux
    port map (
            O => \N__2336\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2333\,
            I => \N__2330\
        );

    \I__323\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2327\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81\
        );

    \I__321\ : InMux
    port map (
            O => \N__2324\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__320\ : InMux
    port map (
            O => \N__2321\,
            I => \N__2318\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2318\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1\
        );

    \I__318\ : InMux
    port map (
            O => \N__2315\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__2312\,
            I => \N__2309\
        );

    \I__316\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2306\,
            I => un2_y_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__314\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2300\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2300\,
            I => un2_y_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__312\ : InMux
    port map (
            O => \N__2297\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__311\ : InMux
    port map (
            O => \N__2294\,
            I => un2_y_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__310\ : CascadeMux
    port map (
            O => \N__2291\,
            I => \N__2287\
        );

    \I__309\ : InMux
    port map (
            O => \N__2290\,
            I => \N__2278\
        );

    \I__308\ : InMux
    port map (
            O => \N__2287\,
            I => \N__2278\
        );

    \I__307\ : InMux
    port map (
            O => \N__2286\,
            I => \N__2278\
        );

    \I__306\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2275\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2278\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2275\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__2270\,
            I => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__301\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2261\,
            I => un2_y_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__298\ : InMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2252\,
            I => un2_y_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__296\ : InMux
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2246\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9\
        );

    \I__294\ : InMux
    port map (
            O => \N__2243\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__293\ : InMux
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2237\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2234\,
            I => \N__2229\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2233\,
            I => \N__2225\
        );

    \I__289\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2221\
        );

    \I__288\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2212\
        );

    \I__287\ : InMux
    port map (
            O => \N__2228\,
            I => \N__2212\
        );

    \I__286\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2212\
        );

    \I__285\ : InMux
    port map (
            O => \N__2224\,
            I => \N__2212\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2221\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2212\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__2207\,
            I => \N__2204\
        );

    \I__281\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2201\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\
        );

    \I__279\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2195\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2195\,
            I => un2_y_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__277\ : InMux
    port map (
            O => \N__2192\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__2189\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_\
        );

    \I__275\ : InMux
    port map (
            O => \N__2186\,
            I => \N__2183\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2183\,
            I => un2_y_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__273\ : InMux
    port map (
            O => \N__2180\,
            I => \N__2176\
        );

    \I__272\ : InMux
    port map (
            O => \N__2179\,
            I => \N__2173\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2176\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2173\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0\
        );

    \I__269\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2164\
        );

    \I__268\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2161\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2164\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2161\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0\
        );

    \I__265\ : InMux
    port map (
            O => \N__2156\,
            I => \N__2153\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2153\,
            I => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0\
        );

    \I__263\ : InMux
    port map (
            O => \N__2150\,
            I => \N__2147\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2147\,
            I => \Pixel_RNOZ0Z_8\
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__2144\,
            I => \N_8_cascade_\
        );

    \I__260\ : InMux
    port map (
            O => \N__2141\,
            I => \N__2138\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2138\,
            I => \N_11\
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__2135\,
            I => \un12_0_1_cascade_\
        );

    \I__257\ : IoInMux
    port map (
            O => \N__2132\,
            I => \N__2129\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2129\,
            I => \N__2126\
        );

    \I__255\ : IoSpan4Mux
    port map (
            O => \N__2126\,
            I => \N__2123\
        );

    \I__254\ : Span4Mux_s1_v
    port map (
            O => \N__2123\,
            I => \N__2120\
        );

    \I__253\ : Span4Mux_h
    port map (
            O => \N__2120\,
            I => \N__2117\
        );

    \I__252\ : Odrv4
    port map (
            O => \N__2117\,
            I => \Pixel_c\
        );

    \I__251\ : InMux
    port map (
            O => \N__2114\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__250\ : CascadeMux
    port map (
            O => \N__2111\,
            I => \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_\
        );

    \I__249\ : InMux
    port map (
            O => \N__2108\,
            I => un2_y_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2105\,
            I => \N__2102\
        );

    \I__247\ : InMux
    port map (
            O => \N__2102\,
            I => \N__2099\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2099\,
            I => \un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\
        );

    \I__245\ : InMux
    port map (
            O => \N__2096\,
            I => \N__2093\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2093\,
            I => \y_RNIA5P7Z0Z_9\
        );

    \I__243\ : InMux
    port map (
            O => \N__2090\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2087\,
            I => \N__2084\
        );

    \I__241\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2081\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2081\,
            I => \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6\
        );

    \I__239\ : InMux
    port map (
            O => \N__2078\,
            I => un2_y_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__238\ : InMux
    port map (
            O => \N__2075\,
            I => \N__2072\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2072\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2\
        );

    \I__236\ : InMux
    port map (
            O => \N__2069\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__235\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2063\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2063\,
            I => un2_y_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__233\ : InMux
    port map (
            O => \N__2060\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__232\ : InMux
    port map (
            O => \N__2057\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__231\ : CascadeMux
    port map (
            O => \N__2054\,
            I => \N__2050\
        );

    \I__230\ : InMux
    port map (
            O => \N__2053\,
            I => \N__2041\
        );

    \I__229\ : InMux
    port map (
            O => \N__2050\,
            I => \N__2041\
        );

    \I__228\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2041\
        );

    \I__227\ : InMux
    port map (
            O => \N__2048\,
            I => \N__2038\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2041\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2038\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2\
        );

    \I__224\ : CascadeMux
    port map (
            O => \N__2033\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_\
        );

    \I__223\ : CascadeMux
    port map (
            O => \N__2030\,
            I => \N__2027\
        );

    \I__222\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2024\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2024\,
            I => un2_y_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__2021\,
            I => \N__2018\
        );

    \I__219\ : InMux
    port map (
            O => \N__2018\,
            I => \N__2015\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2015\,
            I => un2_y_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__217\ : InMux
    port map (
            O => \N__2012\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__216\ : InMux
    port map (
            O => \N__2009\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__215\ : InMux
    port map (
            O => \N__2006\,
            I => un2_y_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__214\ : CascadeMux
    port map (
            O => \N__2003\,
            I => \N__2000\
        );

    \I__213\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1997\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1997\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4\
        );

    \I__211\ : InMux
    port map (
            O => \N__1994\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__210\ : InMux
    port map (
            O => \N__1991\,
            I => \N__1988\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1988\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5\
        );

    \I__208\ : InMux
    port map (
            O => \N__1985\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__207\ : InMux
    port map (
            O => \N__1982\,
            I => \N__1979\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1979\,
            I => un2_y_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__205\ : InMux
    port map (
            O => \N__1976\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__204\ : InMux
    port map (
            O => \N__1973\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__203\ : CascadeMux
    port map (
            O => \N__1970\,
            I => \N__1966\
        );

    \I__202\ : InMux
    port map (
            O => \N__1969\,
            I => \N__1957\
        );

    \I__201\ : InMux
    port map (
            O => \N__1966\,
            I => \N__1957\
        );

    \I__200\ : InMux
    port map (
            O => \N__1965\,
            I => \N__1957\
        );

    \I__199\ : InMux
    port map (
            O => \N__1964\,
            I => \N__1954\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1957\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1954\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5\
        );

    \I__196\ : CascadeMux
    port map (
            O => \N__1949\,
            I => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_\
        );

    \I__195\ : CascadeMux
    port map (
            O => \N__1946\,
            I => \N__1943\
        );

    \I__194\ : InMux
    port map (
            O => \N__1943\,
            I => \N__1940\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1940\,
            I => un2_y_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__192\ : InMux
    port map (
            O => \N__1937\,
            I => \N__1934\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1934\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1\
        );

    \I__190\ : InMux
    port map (
            O => \N__1931\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1928\,
            I => \N__1925\
        );

    \I__188\ : InMux
    port map (
            O => \N__1925\,
            I => \N__1922\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1922\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2\
        );

    \I__186\ : InMux
    port map (
            O => \N__1919\,
            I => un2_y_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__185\ : InMux
    port map (
            O => \N__1916\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__184\ : InMux
    port map (
            O => \N__1913\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__183\ : InMux
    port map (
            O => \N__1910\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__182\ : InMux
    port map (
            O => \N__1907\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__181\ : InMux
    port map (
            O => \N__1904\,
            I => un2_y_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__180\ : CascadeMux
    port map (
            O => \N__1901\,
            I => \N__1898\
        );

    \I__179\ : InMux
    port map (
            O => \N__1898\,
            I => \N__1895\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1895\,
            I => un2_y_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__177\ : InMux
    port map (
            O => \N__1892\,
            I => \N__1889\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1889\,
            I => \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083\
        );

    \I__175\ : InMux
    port map (
            O => \N__1886\,
            I => un2_y_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__174\ : IoInMux
    port map (
            O => \N__1883\,
            I => \N__1880\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1880\,
            I => \N__1877\
        );

    \I__172\ : Span4Mux_s1_h
    port map (
            O => \N__1877\,
            I => \N__1874\
        );

    \I__171\ : Span4Mux_h
    port map (
            O => \N__1874\,
            I => \N__1871\
        );

    \I__170\ : Sp12to4
    port map (
            O => \N__1871\,
            I => \N__1868\
        );

    \I__169\ : Odrv12
    port map (
            O => \N__1868\,
            I => \VGAClock.PixelClock\
        );

    \I__168\ : IoInMux
    port map (
            O => \N__1865\,
            I => \N__1862\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1862\,
            I => \N__1859\
        );

    \I__166\ : IoSpan4Mux
    port map (
            O => \N__1859\,
            I => \N__1856\
        );

    \I__165\ : Odrv4
    port map (
            O => \N__1856\,
            I => \Clock12MHz_c\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_4_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_1_0_\
        );

    \IN_MUX_bfv_4_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un16_x_cry_8,
            carryinitout => \bfn_4_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_y_cry_8,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \VGAClock.PLLOUTCORE_derived_clock_RNIE579\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1883\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3232\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJ6_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1965\,
            in2 => \N__1901\,
            in3 => \N__1916\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8E9_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1892\,
            in2 => \N__1970\,
            in3 => \N__1913\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10B_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1969\,
            in2 => \N__2003\,
            in3 => \N__1910\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAIONN_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2232\,
            in1 => \N__1991\,
            in2 => \N__1946\,
            in3 => \N__1907\,
            lcout => un2_y_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUB_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1982\,
            in2 => \_gnd_net_\,
            in3 => \N__1904\,
            lcout => \un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2641\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2640\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILP083_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2049\,
            in2 => \N__2021\,
            in3 => \N__1886\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOP4_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1937\,
            in2 => \N__2054\,
            in3 => \N__1994\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FI5_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2053\,
            in2 => \N__1928\,
            in3 => \N__1985\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGA9KB_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__1964\,
            in1 => \N__2075\,
            in2 => \N__2030\,
            in3 => \N__1976\,
            lcout => un2_y_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2066\,
            in2 => \_gnd_net_\,
            in3 => \N__1973\,
            lcout => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5\,
            ltout => \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_0_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1949\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2774\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFL1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2286\,
            in2 => \N__2258\,
            in3 => \N__1931\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4E2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2342\,
            in2 => \N__2291\,
            in3 => \N__1919\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9K2_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2290\,
            in2 => \N__2333\,
            in3 => \N__2069\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNI3IEJ5_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2048\,
            in1 => \N__2321\,
            in2 => \N__2267\,
            in3 => \N__2060\,
            lcout => un2_y_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2303\,
            in2 => \_gnd_net_\,
            in3 => \N__2057\,
            lcout => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2\,
            ltout => \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_0_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2033\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3086\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2096\,
            in2 => \N__3306\,
            in3 => \N__2012\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3298\,
            in2 => \N__2105\,
            in3 => \N__2009\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75T2_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3307\,
            in3 => \N__2006\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un33_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2375\,
            in3 => \N__2114\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0\,
            ltout => \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2111\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQ5_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__2412\,
            in1 => \N__2413\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3123\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => un2_y_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2108\,
            lcout => \un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIA5P7_9_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3116\,
            lcout => \y_RNIA5P7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCC_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2186\,
            in2 => \N__2233\,
            in3 => \N__2090\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJI_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2228\,
            in2 => \N__2087\,
            in3 => \N__2078\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_8_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2249\,
            in2 => \N__2234\,
            in3 => \N__2243\,
            lcout => \Pixel_RNOZ0Z_8\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2240\,
            in2 => \N__2207\,
            in3 => \N__2224\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MON_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2198\,
            in2 => \_gnd_net_\,
            in3 => \N__2192\,
            lcout => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0\,
            ltout => \un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_7_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2351\,
            in1 => \N__2180\,
            in2 => \N__2189\,
            in3 => \N__2167\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_6_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__2179\,
            in1 => \N__2168\,
            in2 => \N__3188\,
            in3 => \N__2156\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_2_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__2702\,
            in1 => \N__2150\,
            in2 => \N__2144\,
            in3 => \N__2141\,
            lcout => OPEN,
            ltout => \un12_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000100"
        )
    port map (
            in0 => \N__2801\,
            in1 => \N__2591\,
            in2 => \N__2135\,
            in3 => \N__2552\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2735\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIG21_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2430\,
            in2 => \N__2360\,
            in3 => \N__2336\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68K81_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2477\,
            in2 => \N__2435\,
            in3 => \N__2324\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHB1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2434\,
            in2 => \N__2462\,
            in3 => \N__2315\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI678Q2_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2285\,
            in1 => \N__2444\,
            in2 => \N__2312\,
            in3 => \N__2297\,
            lcout => un2_y_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2387\,
            in2 => \_gnd_net_\,
            in3 => \N__2294\,
            lcout => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91\,
            ltout => \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_0_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2270\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3043\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERG_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2366\,
            in2 => \N__3292\,
            in3 => \N__2471\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJ_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2468\,
            in2 => \N__3294\,
            in3 => \N__2453\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KO_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2450\,
            in2 => \N__3293\,
            in3 => \N__2438\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0\,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNIAP1U_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2429\,
            in1 => \N__2414\,
            in2 => \N__2396\,
            in3 => \N__2381\,
            lcout => un2_y_if_generate_plus_mult1_un47_sum_axb_7,
            ltout => OPEN,
            carryin => un2_y_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => un2_y_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2378\,
            lcout => \un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNI94P7_8_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3087\,
            lcout => \y_RNI94P7Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_y_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_11_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2996\,
            in2 => \N__2701\,
            in3 => \N__3178\,
            lcout => \G_7_i_a4_0_0\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => un4_y_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_y_cry_1_THRU_LUT4_0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3182\,
            in2 => \_gnd_net_\,
            in3 => \N__2501\,
            lcout => \un4_y_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => un4_y_cry_1,
            carryout => un4_y_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_y_cry_2_THRU_LUT4_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3231\,
            in2 => \_gnd_net_\,
            in3 => \N__2498\,
            lcout => \un4_y_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => un4_y_cry_2,
            carryout => un4_y_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_4_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2967\,
            in1 => \N__2629\,
            in2 => \_gnd_net_\,
            in3 => \N__2495\,
            lcout => \yZ0Z_4\,
            ltout => OPEN,
            carryin => un4_y_cry_3,
            carryout => un4_y_cry_4,
            clk => \N__3712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_5_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2957\,
            in1 => \N__2773\,
            in2 => \_gnd_net_\,
            in3 => \N__2492\,
            lcout => \yZ0Z_5\,
            ltout => OPEN,
            carryin => un4_y_cry_4,
            carryout => un4_y_cry_5,
            clk => \N__3712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2968\,
            in1 => \N__2734\,
            in2 => \_gnd_net_\,
            in3 => \N__2489\,
            lcout => \yZ0Z_6\,
            ltout => OPEN,
            carryin => un4_y_cry_5,
            carryout => un4_y_cry_6,
            clk => \N__3712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_7_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2958\,
            in1 => \N__3048\,
            in2 => \_gnd_net_\,
            in3 => \N__2486\,
            lcout => \yZ0Z_7\,
            ltout => OPEN,
            carryin => un4_y_cry_6,
            carryout => un4_y_cry_7,
            clk => \N__3712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_8_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2969\,
            in1 => \N__3093\,
            in2 => \_gnd_net_\,
            in3 => \N__2483\,
            lcout => \yZ0Z_8\,
            ltout => OPEN,
            carryin => un4_y_cry_7,
            carryout => un4_y_cry_8,
            clk => \N__3712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_9_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__3020\,
            in1 => \N__2966\,
            in2 => \N__3129\,
            in3 => \N__2480\,
            lcout => \yZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un16_x_cry_1_c_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2834\,
            in2 => \N__2876\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_1_0_\,
            carryout => un16_x_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_2_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2888\,
            in2 => \_gnd_net_\,
            in3 => \N__2534\,
            lcout => \xZ0Z_2\,
            ltout => OPEN,
            carryin => un16_x_cry_1,
            carryout => un16_x_cry_2,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_3_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2853\,
            in2 => \_gnd_net_\,
            in3 => \N__2531\,
            lcout => \xZ0Z_3\,
            ltout => OPEN,
            carryin => un16_x_cry_2,
            carryout => un16_x_cry_3,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_4_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3459\,
            in2 => \_gnd_net_\,
            in3 => \N__2528\,
            lcout => \xZ0Z_4\,
            ltout => OPEN,
            carryin => un16_x_cry_3,
            carryout => un16_x_cry_4,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_5_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2928\,
            in1 => \N__3676\,
            in2 => \_gnd_net_\,
            in3 => \N__2525\,
            lcout => \xZ0Z_5\,
            ltout => OPEN,
            carryin => un16_x_cry_4,
            carryout => un16_x_cry_5,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_6_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3936\,
            in2 => \_gnd_net_\,
            in3 => \N__2522\,
            lcout => \xZ0Z_6\,
            ltout => OPEN,
            carryin => un16_x_cry_5,
            carryout => un16_x_cry_6,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_7_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3972\,
            in2 => \_gnd_net_\,
            in3 => \N__2519\,
            lcout => \xZ0Z_7\,
            ltout => OPEN,
            carryin => un16_x_cry_6,
            carryout => un16_x_cry_7,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_8_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2927\,
            in1 => \N__3361\,
            in2 => \_gnd_net_\,
            in3 => \N__2516\,
            lcout => \xZ0Z_8\,
            ltout => OPEN,
            carryin => un16_x_cry_7,
            carryout => un16_x_cry_8,
            clk => \N__3716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_9_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3412\,
            in1 => \N__2929\,
            in2 => \_gnd_net_\,
            in3 => \N__2513\,
            lcout => \xZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_10_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__3675\,
            in1 => \N__3932\,
            in2 => \N__3460\,
            in3 => \N__3968\,
            lcout => un8_xlt9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_4_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111100"
        )
    port map (
            in0 => \N__3419\,
            in1 => \N__3359\,
            in2 => \N__2510\,
            in3 => \N__3411\,
            lcout => OPEN,
            ltout => \Pixel_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__3748\,
            in1 => \_gnd_net_\,
            in2 => \N__2594\,
            in3 => \_gnd_net_\,
            lcout => \Pixel_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3462\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2572\,
            in2 => \N__2543\,
            in3 => \N__2579\,
            lcout => \un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_5_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3515\,
            in2 => \N__3781\,
            in3 => \N__2576\,
            lcout => \Pixel_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2573\,
            in2 => \N__3506\,
            in3 => \N__3774\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3494\,
            in2 => \_gnd_net_\,
            in3 => \N__2564\,
            lcout => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0\,
            ltout => \un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_1_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111110110000"
        )
    port map (
            in0 => \N__3463\,
            in1 => \N__2815\,
            in2 => \N__2561\,
            in3 => \N__2558\,
            lcout => un2_x_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI5UL6_5_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3684\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_3_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001010001100"
        )
    port map (
            in0 => \N__2858\,
            in1 => \N__2816\,
            in2 => \N__3467\,
            in3 => \N__2807\,
            lcout => un13lt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIQ64V_4_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2780\,
            in1 => \N__2741\,
            in2 => \N__2645\,
            in3 => \N__3056\,
            lcout => OPEN,
            ltout => \un1_ylto9_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIMA162_3_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2663\,
            in1 => \N__3216\,
            in2 => \N__2792\,
            in3 => \N__3170\,
            lcout => un1_y,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_3_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001111000"
        )
    port map (
            in0 => \N__2954\,
            in1 => \N__2789\,
            in2 => \N__3230\,
            in3 => \N__3016\,
            lcout => \yZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__2687\,
            in1 => \N__2955\,
            in2 => \_gnd_net_\,
            in3 => \N__2991\,
            lcout => \yZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIGS3V_0_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2691\,
            in1 => \N__2779\,
            in2 => \N__2995\,
            in3 => \N__2740\,
            lcout => y_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIL6BN_9_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2686\,
            in1 => \N__3094\,
            in2 => \_gnd_net_\,
            in3 => \N__3130\,
            lcout => un1_ylto9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_2_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100100000"
        )
    port map (
            in0 => \N__2953\,
            in1 => \N__3015\,
            in2 => \N__2657\,
            in3 => \N__3174\,
            lcout => \yZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIM24V_9_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2639\,
            in1 => \N__3217\,
            in2 => \N__3183\,
            in3 => \N__3131\,
            lcout => OPEN,
            ltout => \y_12_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_RNIN6QD2_7_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3095\,
            in1 => \N__3065\,
            in2 => \N__3059\,
            in3 => \N__3055\,
            lcout => y_12_8,
            ltout => \y_12_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2990\,
            in2 => \N__2999\,
            in3 => \N__2956\,
            lcout => \yZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2832\,
            lcout => \xZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2872\,
            in2 => \_gnd_net_\,
            in3 => \N__2833\,
            lcout => \xZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3718\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNIRVNQ_9_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3935\,
            in1 => \N__3360\,
            in2 => \N__3413\,
            in3 => \N__3458\,
            lcout => OPEN,
            ltout => \un11_x_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNID8R22_9_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3638\,
            in2 => \N__2972\,
            in3 => \N__3479\,
            lcout => \x_RNID8R22Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI6ANQ_1_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2887\,
            in1 => \N__2871\,
            in2 => \N__2857\,
            in3 => \N__2831\,
            lcout => un11_x_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3405\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => un2_x_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3485\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => \un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3482\,
            in3 => \_gnd_net_\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_9_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3634\,
            in1 => \N__3478\,
            in2 => \N__3461\,
            in3 => \N__3933\,
            lcout => un4_xlt9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI81M6_8_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3358\,
            lcout => un2_x_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI92M6_9_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSyncZ0_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__3407\,
            in1 => \N__3329\,
            in2 => \N__3685\,
            in3 => \N__3934\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_RNO_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3365\,
            in3 => \N__3978\,
            lcout => un1_xlto9_0,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3323\,
            in2 => \_gnd_net_\,
            in3 => \N__3317\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3314\,
            in2 => \N__3305\,
            in3 => \N__3236\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3613\,
            in1 => \N__3521\,
            in2 => \N__3542\,
            in3 => \N__3551\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3548\,
            lcout => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0\,
            ltout => \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3545\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3532\,
            in2 => \_gnd_net_\,
            in3 => \N__3538\,
            lcout => \un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3680\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3793\,
            in2 => \N__3761\,
            in3 => \N__3509\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3809\,
            in2 => \N__3890\,
            in3 => \N__3497\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3782\,
            in1 => \N__3794\,
            in2 => \N__3857\,
            in3 => \N__3488\,
            lcout => un2_x_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3827\,
            in2 => \_gnd_net_\,
            in3 => \N__3785\,
            lcout => \un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI6VL6_6_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3944\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSyncZ0_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3752\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNICUBD_5_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3979\,
            in2 => \_gnd_net_\,
            in3 => \N__3686\,
            lcout => un11_x_4,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3623\,
            in2 => \N__3590\,
            in3 => \N__3617\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3614\,
            in2 => \N__3602\,
            in3 => \N__3593\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3877\,
            in1 => \N__3589\,
            in2 => \N__3575\,
            in3 => \N__3566\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3563\,
            in2 => \_gnd_net_\,
            in3 => \N__3557\,
            lcout => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1\,
            ltout => \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3554\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \x_RNI70M6_7_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3980\,
            lcout => un2_x_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3943\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3844\,
            in2 => \N__3899\,
            in3 => \N__3881\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3878\,
            in2 => \N__3866\,
            in3 => \N__3848\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2\,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3808\,
            in1 => \N__3845\,
            in2 => \N__3836\,
            in3 => \N__3821\,
            lcout => un2_x_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un2_x_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un2_x_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3818\,
            in2 => \_gnd_net_\,
            in3 => \N__3812\,
            lcout => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2\,
            ltout => \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3797\,
            in3 => \_gnd_net_\,
            lcout => un2_x_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
