// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 17:10:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4454;
    wire N__4453;
    wire N__4452;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4436;
    wire N__4435;
    wire N__4434;
    wire N__4427;
    wire N__4426;
    wire N__4425;
    wire N__4418;
    wire N__4417;
    wire N__4416;
    wire N__4409;
    wire N__4408;
    wire N__4407;
    wire N__4390;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4335;
    wire N__4334;
    wire N__4333;
    wire N__4326;
    wire N__4323;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4263;
    wire N__4262;
    wire N__4259;
    wire N__4258;
    wire N__4255;
    wire N__4254;
    wire N__4251;
    wire N__4242;
    wire N__4237;
    wire N__4234;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4131;
    wire N__4128;
    wire N__4127;
    wire N__4126;
    wire N__4125;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4014;
    wire N__4013;
    wire N__4010;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3988;
    wire N__3985;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3954;
    wire N__3953;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3928;
    wire N__3927;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3912;
    wire N__3911;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3883;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3861;
    wire N__3860;
    wire N__3857;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3845;
    wire N__3842;
    wire N__3835;
    wire N__3832;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3817;
    wire N__3814;
    wire N__3813;
    wire N__3812;
    wire N__3811;
    wire N__3810;
    wire N__3809;
    wire N__3808;
    wire N__3807;
    wire N__3806;
    wire N__3805;
    wire N__3804;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3793;
    wire N__3790;
    wire N__3789;
    wire N__3788;
    wire N__3781;
    wire N__3778;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3747;
    wire N__3746;
    wire N__3743;
    wire N__3734;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3697;
    wire N__3688;
    wire N__3687;
    wire N__3686;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3658;
    wire N__3657;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3642;
    wire N__3639;
    wire N__3638;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3609;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3532;
    wire N__3531;
    wire N__3530;
    wire N__3529;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3525;
    wire N__3508;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3495;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3476;
    wire N__3473;
    wire N__3466;
    wire N__3465;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3448;
    wire N__3447;
    wire N__3446;
    wire N__3445;
    wire N__3442;
    wire N__3437;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3403;
    wire N__3402;
    wire N__3399;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3376;
    wire N__3375;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3367;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3343;
    wire N__3340;
    wire N__3331;
    wire N__3328;
    wire N__3327;
    wire N__3326;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3314;
    wire N__3311;
    wire N__3304;
    wire N__3301;
    wire N__3300;
    wire N__3299;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3287;
    wire N__3284;
    wire N__3277;
    wire N__3274;
    wire N__3273;
    wire N__3272;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3192;
    wire N__3191;
    wire N__3188;
    wire N__3187;
    wire N__3184;
    wire N__3183;
    wire N__3180;
    wire N__3171;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3156;
    wire N__3155;
    wire N__3152;
    wire N__3151;
    wire N__3150;
    wire N__3147;
    wire N__3140;
    wire N__3137;
    wire N__3130;
    wire N__3129;
    wire N__3128;
    wire N__3127;
    wire N__3126;
    wire N__3123;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3109;
    wire N__3106;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3093;
    wire N__3092;
    wire N__3089;
    wire N__3084;
    wire N__3079;
    wire N__3076;
    wire N__3067;
    wire N__3066;
    wire N__3065;
    wire N__3064;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3052;
    wire N__3049;
    wire N__3040;
    wire N__3037;
    wire N__3036;
    wire N__3035;
    wire N__3034;
    wire N__3033;
    wire N__3032;
    wire N__3029;
    wire N__3024;
    wire N__3019;
    wire N__3016;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2977;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2919;
    wire N__2918;
    wire N__2915;
    wire N__2910;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2887;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2824;
    wire N__2823;
    wire N__2822;
    wire N__2821;
    wire N__2820;
    wire N__2819;
    wire N__2816;
    wire N__2811;
    wire N__2808;
    wire N__2803;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2773;
    wire N__2770;
    wire N__2763;
    wire N__2758;
    wire N__2755;
    wire N__2754;
    wire N__2753;
    wire N__2750;
    wire N__2745;
    wire N__2740;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2721;
    wire N__2718;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2688;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2668;
    wire N__2665;
    wire N__2662;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2580;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2572;
    wire N__2569;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2527;
    wire N__2524;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2506;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2473;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2431;
    wire N__2428;
    wire N__2427;
    wire N__2422;
    wire N__2419;
    wire N__2418;
    wire N__2415;
    wire N__2410;
    wire N__2407;
    wire N__2406;
    wire N__2403;
    wire N__2402;
    wire N__2399;
    wire N__2394;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2382;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2374;
    wire N__2371;
    wire N__2366;
    wire N__2359;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2343;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2313;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2299;
    wire N__2296;
    wire N__2293;
    wire N__2290;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2262;
    wire N__2259;
    wire N__2256;
    wire N__2253;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2239;
    wire N__2236;
    wire N__2233;
    wire N__2230;
    wire N__2227;
    wire N__2224;
    wire N__2221;
    wire N__2218;
    wire N__2215;
    wire N__2212;
    wire N__2209;
    wire N__2206;
    wire N__2203;
    wire N__2200;
    wire N__2197;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2187;
    wire N__2184;
    wire N__2181;
    wire N__2176;
    wire N__2173;
    wire N__2170;
    wire N__2167;
    wire N__2164;
    wire N__2161;
    wire N__2158;
    wire N__2155;
    wire N__2152;
    wire N__2149;
    wire N__2146;
    wire N__2143;
    wire N__2140;
    wire N__2137;
    wire N__2134;
    wire N__2133;
    wire N__2130;
    wire N__2129;
    wire N__2126;
    wire N__2121;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2104;
    wire N__2103;
    wire N__2098;
    wire N__2095;
    wire N__2092;
    wire N__2089;
    wire N__2086;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2071;
    wire N__2068;
    wire \VGAClock.PixelClock ;
    wire Clock12MHz_c;
    wire VCCG0;
    wire GNDG0;
    wire bfn_7_3_0_;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_4;
    wire Pixel_1_RNOZ0Z_6;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_i;
    wire bfn_7_4_0_;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_i;
    wire bfn_7_5_0_;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_;
    wire un13_beamx_6_cascade_;
    wire un13_beamx_5;
    wire un1_beamylto9_4;
    wire un1_beamylto9_5_cascade_;
    wire un1_beamy_cascade_;
    wire VSync_c;
    wire un11_beamx_3_cascade_;
    wire un11_beamx_6;
    wire un11_beamx_6_cascade_;
    wire bfn_8_2_0_;
    wire un1_beamX_if_generate_plus_mult1_un68_sum;
    wire un5_visiblex_cry_4;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire un5_visiblex_cry_8;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_;
    wire un5_visiblex_i;
    wire bfn_8_3_0_;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un54_sum;
    wire un5_visiblex_i_24;
    wire un1_beamX_if_generate_plus_mult1_un61_sum;
    wire bfn_8_4_0_;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_i;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un61_sum_i_8;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0;
    wire un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631;
    wire bfn_8_5_0_;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_6;
    wire bfn_8_6_0_;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_axb_6;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_i_0;
    wire un5_visibley_cry_7_c_RNI1L4CZ0Z_0;
    wire un5_visibley_cry_8_c_RNI3O5CZ0Z_0;
    wire bfn_8_7_0_;
    wire un4_beamy_cry_1;
    wire un4_beamy_cry_2;
    wire un4_beamy_cry_3;
    wire un4_beamy_cry_4;
    wire un4_beamy_cry_5;
    wire un4_beamy_cry_6;
    wire un4_beamy_cry_7;
    wire un4_beamy_cry_8;
    wire bfn_8_8_0_;
    wire beamXZ0Z_0;
    wire beamXZ0Z_1;
    wire bfn_9_1_0_;
    wire beamXZ0Z_2;
    wire un16_beamx_cry_1;
    wire beamXZ0Z_3;
    wire un16_beamx_cry_2;
    wire un16_beamx_cry_3;
    wire un16_beamx_cry_4;
    wire un16_beamx_cry_5;
    wire un16_beamx_cry_6;
    wire un16_beamx_cry_7;
    wire un16_beamx_cry_8;
    wire bfn_9_2_0_;
    wire un1_beamy;
    wire un4_beamxlt9;
    wire Pixel_0_sqmuxa_0_cascade_;
    wire un11_beamx_1;
    wire beamXZ0Z_4;
    wire un8_beamxlt9_0;
    wire beamXZ0Z_9;
    wire beamXZ0Z_7;
    wire beamXZ0Z_6;
    wire beamXZ0Z_8;
    wire un1_beamxlto9_0_cascade_;
    wire beamXZ0Z_5;
    wire HSync_c;
    wire un5_visiblex_cry_7_c_RNIVZ0Z952;
    wire bfn_9_3_0_;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_c5_i;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_beamX_if_generate_plus_mult1_un40_sum_c5;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_0;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_;
    wire un1_beamX_if_generate_plus_mult1_un47_sum_i_8;
    wire bfn_9_4_0_;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un47_sum_i_0;
    wire un13_beamx;
    wire beamX_RNIVEM1Z0Z_4;
    wire beamYZ0Z_0;
    wire bfn_9_7_0_;
    wire beamYZ0Z_1;
    wire un5_visibley_cry_0;
    wire beamYZ0Z_2;
    wire un5_visibley_cry_1;
    wire beamYZ0Z_3;
    wire un5_visibley_cry_2;
    wire beamYZ0Z_4;
    wire un5_visibley_cry_3;
    wire beamYZ0Z_5;
    wire un1_visibley_if_generate_plus_mult1_un54_sum;
    wire un5_visibley_cry_4;
    wire beamYZ0Z_6;
    wire un1_visibley_if_generate_plus_mult1_un47_sum;
    wire un5_visibley_cry_5;
    wire beamYZ0Z_7;
    wire un1_visibley_if_generate_plus_mult1_un40_sum;
    wire un5_visibley_cry_6;
    wire un5_visibley_cry_7;
    wire CONSTANT_ONE_NET;
    wire beamYZ0Z_8;
    wire un5_visibley_cry_7_c_RNI1L4CZ0;
    wire bfn_9_8_0_;
    wire beamYZ0Z_9;
    wire un5_visibley_cry_8;
    wire un1_visibley_if_generate_plus_mult1_un33_sum_axb_3;
    wire N_8_cascade_;
    wire un1_beamX_27;
    wire Pixel_0_sqmuxa_1;
    wire un13_0_1_cascade_;
    wire un12lt10;
    wire Pixel_c;
    wire PixelClock_g;
    wire bfn_11_3_0_;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_3;
    wire Pixel_1_RNOZ0Z_9;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0;
    wire N_11;
    wire un1_visibley_if_generate_plus_mult1_un75_sum;
    wire un5_visibley_cry_0_c_RNIJVSBZ0;
    wire G_7_i_a4_0_0;
    wire bfn_11_4_0_;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_i_0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_i_0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum;
    wire bfn_12_4_0_;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_i_7;
    wire un1_visibley_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0;
    wire un1_visibley_if_generate_plus_mult1_un61_sum;
    wire un1_visibley_if_generate_plus_mult1_un61_sum_i_0;
    wire _gnd_net_;

    defparam \VGAClock.PixelClock_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \VGAClock.PixelClock_inst .TEST_MODE=1'b0;
    defparam \VGAClock.PixelClock_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \VGAClock.PixelClock_inst .PLLOUT_SELECT="GENCLK";
    defparam \VGAClock.PixelClock_inst .FILTER_RANGE=3'b001;
    defparam \VGAClock.PixelClock_inst .FEEDBACK_PATH="SIMPLE";
    defparam \VGAClock.PixelClock_inst .FDA_RELATIVE=4'b0000;
    defparam \VGAClock.PixelClock_inst .FDA_FEEDBACK=4'b0000;
    defparam \VGAClock.PixelClock_inst .ENABLE_ICEGATE=1'b0;
    defparam \VGAClock.PixelClock_inst .DIVR=4'b0000;
    defparam \VGAClock.PixelClock_inst .DIVQ=3'b100;
    defparam \VGAClock.PixelClock_inst .DIVF=7'b1001010;
    defparam \VGAClock.PixelClock_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \VGAClock.PixelClock_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\VGAClock.PixelClock ),
            .REFERENCECLK(N__2077),
            .RESETB(N__3789),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__4463),
            .DIN(N__4462),
            .DOUT(N__4461),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__4463),
            .PADOUT(N__4462),
            .PADIN(N__4461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__4454),
            .DIN(N__4453),
            .DOUT(N__4452),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__4454),
            .PADOUT(N__4453),
            .PADIN(N__4452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2262),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__4445),
            .DIN(N__4444),
            .DOUT(N__4443),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__4445),
            .PADOUT(N__4444),
            .PADIN(N__4443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__4436),
            .DIN(N__4435),
            .DOUT(N__4434),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__4436),
            .PADOUT(N__4435),
            .PADIN(N__4434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3555),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__4427),
            .DIN(N__4426),
            .DOUT(N__4425),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__4427),
            .PADOUT(N__4426),
            .PADIN(N__4425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__4418),
            .DIN(N__4417),
            .DOUT(N__4416),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__4418),
            .PADOUT(N__4417),
            .PADIN(N__4416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__4409),
            .DIN(N__4408),
            .DOUT(N__4407),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__4409),
            .PADOUT(N__4408),
            .PADIN(N__4407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3007),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__957 (
            .O(N__4390),
            .I(N__4386));
    InMux I__956 (
            .O(N__4389),
            .I(N__4383));
    LocalMux I__955 (
            .O(N__4386),
            .I(N__4380));
    LocalMux I__954 (
            .O(N__4383),
            .I(N__4377));
    Span4Mux_v I__953 (
            .O(N__4380),
            .I(N__4374));
    Span4Mux_s2_h I__952 (
            .O(N__4377),
            .I(N__4371));
    Odrv4 I__951 (
            .O(N__4374),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum));
    Odrv4 I__950 (
            .O(N__4371),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum));
    CascadeMux I__949 (
            .O(N__4366),
            .I(N__4363));
    InMux I__948 (
            .O(N__4363),
            .I(N__4360));
    LocalMux I__947 (
            .O(N__4360),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49));
    InMux I__946 (
            .O(N__4357),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__945 (
            .O(N__4354),
            .I(N__4351));
    LocalMux I__944 (
            .O(N__4351),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4));
    InMux I__943 (
            .O(N__4348),
            .I(N__4345));
    LocalMux I__942 (
            .O(N__4345),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0));
    InMux I__941 (
            .O(N__4342),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__940 (
            .O(N__4339),
            .I(N__4335));
    InMux I__939 (
            .O(N__4338),
            .I(N__4326));
    InMux I__938 (
            .O(N__4335),
            .I(N__4326));
    InMux I__937 (
            .O(N__4334),
            .I(N__4326));
    InMux I__936 (
            .O(N__4333),
            .I(N__4323));
    LocalMux I__935 (
            .O(N__4326),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8));
    LocalMux I__934 (
            .O(N__4323),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8));
    CascadeMux I__933 (
            .O(N__4318),
            .I(N__4315));
    InMux I__932 (
            .O(N__4315),
            .I(N__4312));
    LocalMux I__931 (
            .O(N__4312),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6));
    InMux I__930 (
            .O(N__4309),
            .I(N__4306));
    LocalMux I__929 (
            .O(N__4306),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0));
    InMux I__928 (
            .O(N__4303),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__927 (
            .O(N__4300),
            .I(N__4297));
    LocalMux I__926 (
            .O(N__4297),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7));
    CascadeMux I__925 (
            .O(N__4294),
            .I(N__4291));
    InMux I__924 (
            .O(N__4291),
            .I(N__4288));
    LocalMux I__923 (
            .O(N__4288),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_i_7));
    CascadeMux I__922 (
            .O(N__4285),
            .I(N__4282));
    InMux I__921 (
            .O(N__4282),
            .I(N__4279));
    LocalMux I__920 (
            .O(N__4279),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__919 (
            .O(N__4276),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__918 (
            .O(N__4273),
            .I(N__4270));
    LocalMux I__917 (
            .O(N__4270),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__916 (
            .O(N__4267),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__915 (
            .O(N__4264),
            .I(N__4259));
    CascadeMux I__914 (
            .O(N__4263),
            .I(N__4255));
    InMux I__913 (
            .O(N__4262),
            .I(N__4251));
    InMux I__912 (
            .O(N__4259),
            .I(N__4242));
    InMux I__911 (
            .O(N__4258),
            .I(N__4242));
    InMux I__910 (
            .O(N__4255),
            .I(N__4242));
    InMux I__909 (
            .O(N__4254),
            .I(N__4242));
    LocalMux I__908 (
            .O(N__4251),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0));
    LocalMux I__907 (
            .O(N__4242),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0));
    InMux I__906 (
            .O(N__4237),
            .I(N__4234));
    LocalMux I__905 (
            .O(N__4234),
            .I(N__4230));
    InMux I__904 (
            .O(N__4233),
            .I(N__4227));
    Span4Mux_v I__903 (
            .O(N__4230),
            .I(N__4224));
    LocalMux I__902 (
            .O(N__4227),
            .I(N__4221));
    Sp12to4 I__901 (
            .O(N__4224),
            .I(N__4218));
    Span4Mux_v I__900 (
            .O(N__4221),
            .I(N__4215));
    Odrv12 I__899 (
            .O(N__4218),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum));
    Odrv4 I__898 (
            .O(N__4215),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum));
    CascadeMux I__897 (
            .O(N__4210),
            .I(N__4207));
    InMux I__896 (
            .O(N__4207),
            .I(N__4204));
    LocalMux I__895 (
            .O(N__4204),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_i_0));
    CascadeMux I__894 (
            .O(N__4201),
            .I(N__4198));
    InMux I__893 (
            .O(N__4198),
            .I(N__4195));
    LocalMux I__892 (
            .O(N__4195),
            .I(N__4192));
    Odrv12 I__891 (
            .O(N__4192),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__890 (
            .O(N__4189),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__889 (
            .O(N__4186),
            .I(N__4183));
    LocalMux I__888 (
            .O(N__4183),
            .I(N__4180));
    Odrv4 I__887 (
            .O(N__4180),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1));
    InMux I__886 (
            .O(N__4177),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__885 (
            .O(N__4174),
            .I(N__4171));
    InMux I__884 (
            .O(N__4171),
            .I(N__4168));
    LocalMux I__883 (
            .O(N__4168),
            .I(N__4165));
    Odrv4 I__882 (
            .O(N__4165),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2));
    InMux I__881 (
            .O(N__4162),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__880 (
            .O(N__4159),
            .I(N__4156));
    LocalMux I__879 (
            .O(N__4156),
            .I(N__4153));
    Odrv4 I__878 (
            .O(N__4153),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3));
    InMux I__877 (
            .O(N__4150),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__876 (
            .O(N__4147),
            .I(N__4144));
    LocalMux I__875 (
            .O(N__4144),
            .I(N__4141));
    Odrv4 I__874 (
            .O(N__4141),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__873 (
            .O(N__4138),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__872 (
            .O(N__4135),
            .I(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_));
    CascadeMux I__871 (
            .O(N__4132),
            .I(N__4128));
    InMux I__870 (
            .O(N__4131),
            .I(N__4116));
    InMux I__869 (
            .O(N__4128),
            .I(N__4116));
    InMux I__868 (
            .O(N__4127),
            .I(N__4116));
    InMux I__867 (
            .O(N__4126),
            .I(N__4116));
    InMux I__866 (
            .O(N__4125),
            .I(N__4113));
    LocalMux I__865 (
            .O(N__4116),
            .I(N__4110));
    LocalMux I__864 (
            .O(N__4113),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4));
    Odrv4 I__863 (
            .O(N__4110),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4));
    CascadeMux I__862 (
            .O(N__4105),
            .I(N__4102));
    InMux I__861 (
            .O(N__4102),
            .I(N__4099));
    LocalMux I__860 (
            .O(N__4099),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__859 (
            .O(N__4096),
            .I(N__4093));
    LocalMux I__858 (
            .O(N__4093),
            .I(N__4090));
    Odrv4 I__857 (
            .O(N__4090),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__856 (
            .O(N__4087),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__855 (
            .O(N__4084),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__854 (
            .O(N__4081),
            .I(N__4078));
    LocalMux I__853 (
            .O(N__4078),
            .I(Pixel_1_RNOZ0Z_9));
    InMux I__852 (
            .O(N__4075),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__851 (
            .O(N__4072),
            .I(N__4069));
    InMux I__850 (
            .O(N__4069),
            .I(N__4066));
    LocalMux I__849 (
            .O(N__4066),
            .I(un1_visibley_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__848 (
            .O(N__4063),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__847 (
            .O(N__4060),
            .I(N__4057));
    LocalMux I__846 (
            .O(N__4057),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11));
    InMux I__845 (
            .O(N__4054),
            .I(N__4050));
    InMux I__844 (
            .O(N__4053),
            .I(N__4047));
    LocalMux I__843 (
            .O(N__4050),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0));
    LocalMux I__842 (
            .O(N__4047),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0));
    CascadeMux I__841 (
            .O(N__4042),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_));
    InMux I__840 (
            .O(N__4039),
            .I(N__4035));
    InMux I__839 (
            .O(N__4038),
            .I(N__4032));
    LocalMux I__838 (
            .O(N__4035),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0));
    LocalMux I__837 (
            .O(N__4032),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0));
    InMux I__836 (
            .O(N__4027),
            .I(N__4024));
    LocalMux I__835 (
            .O(N__4024),
            .I(N_11));
    CascadeMux I__834 (
            .O(N__4021),
            .I(N__4018));
    InMux I__833 (
            .O(N__4018),
            .I(N__4015));
    LocalMux I__832 (
            .O(N__4015),
            .I(N__4010));
    InMux I__831 (
            .O(N__4014),
            .I(N__4005));
    InMux I__830 (
            .O(N__4013),
            .I(N__4005));
    Span4Mux_s2_h I__829 (
            .O(N__4010),
            .I(N__4002));
    LocalMux I__828 (
            .O(N__4005),
            .I(N__3999));
    Span4Mux_v I__827 (
            .O(N__4002),
            .I(N__3996));
    Span4Mux_s2_h I__826 (
            .O(N__3999),
            .I(N__3993));
    Odrv4 I__825 (
            .O(N__3996),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum));
    Odrv4 I__824 (
            .O(N__3993),
            .I(un1_visibley_if_generate_plus_mult1_un75_sum));
    InMux I__823 (
            .O(N__3988),
            .I(N__3985));
    LocalMux I__822 (
            .O(N__3985),
            .I(N__3981));
    InMux I__821 (
            .O(N__3984),
            .I(N__3978));
    Span4Mux_s2_v I__820 (
            .O(N__3981),
            .I(N__3975));
    LocalMux I__819 (
            .O(N__3978),
            .I(N__3972));
    Span4Mux_v I__818 (
            .O(N__3975),
            .I(N__3969));
    Span4Mux_s2_h I__817 (
            .O(N__3972),
            .I(N__3966));
    Odrv4 I__816 (
            .O(N__3969),
            .I(un5_visibley_cry_0_c_RNIJVSBZ0));
    Odrv4 I__815 (
            .O(N__3966),
            .I(un5_visibley_cry_0_c_RNIJVSBZ0));
    InMux I__814 (
            .O(N__3961),
            .I(N__3958));
    LocalMux I__813 (
            .O(N__3958),
            .I(G_7_i_a4_0_0));
    CascadeMux I__812 (
            .O(N__3955),
            .I(N__3949));
    InMux I__811 (
            .O(N__3954),
            .I(N__3946));
    InMux I__810 (
            .O(N__3953),
            .I(N__3943));
    InMux I__809 (
            .O(N__3952),
            .I(N__3940));
    InMux I__808 (
            .O(N__3949),
            .I(N__3937));
    LocalMux I__807 (
            .O(N__3946),
            .I(beamYZ0Z_5));
    LocalMux I__806 (
            .O(N__3943),
            .I(beamYZ0Z_5));
    LocalMux I__805 (
            .O(N__3940),
            .I(beamYZ0Z_5));
    LocalMux I__804 (
            .O(N__3937),
            .I(beamYZ0Z_5));
    InMux I__803 (
            .O(N__3928),
            .I(N__3922));
    InMux I__802 (
            .O(N__3927),
            .I(N__3922));
    LocalMux I__801 (
            .O(N__3922),
            .I(N__3919));
    Odrv4 I__800 (
            .O(N__3919),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum));
    InMux I__799 (
            .O(N__3916),
            .I(un5_visibley_cry_4));
    CascadeMux I__798 (
            .O(N__3913),
            .I(N__3907));
    CascadeMux I__797 (
            .O(N__3912),
            .I(N__3904));
    InMux I__796 (
            .O(N__3911),
            .I(N__3901));
    InMux I__795 (
            .O(N__3910),
            .I(N__3898));
    InMux I__794 (
            .O(N__3907),
            .I(N__3895));
    InMux I__793 (
            .O(N__3904),
            .I(N__3892));
    LocalMux I__792 (
            .O(N__3901),
            .I(beamYZ0Z_6));
    LocalMux I__791 (
            .O(N__3898),
            .I(beamYZ0Z_6));
    LocalMux I__790 (
            .O(N__3895),
            .I(beamYZ0Z_6));
    LocalMux I__789 (
            .O(N__3892),
            .I(beamYZ0Z_6));
    CascadeMux I__788 (
            .O(N__3883),
            .I(N__3879));
    InMux I__787 (
            .O(N__3882),
            .I(N__3876));
    InMux I__786 (
            .O(N__3879),
            .I(N__3873));
    LocalMux I__785 (
            .O(N__3876),
            .I(N__3868));
    LocalMux I__784 (
            .O(N__3873),
            .I(N__3868));
    Odrv4 I__783 (
            .O(N__3868),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum));
    InMux I__782 (
            .O(N__3865),
            .I(un5_visibley_cry_5));
    CascadeMux I__781 (
            .O(N__3862),
            .I(N__3857));
    CascadeMux I__780 (
            .O(N__3861),
            .I(N__3853));
    InMux I__779 (
            .O(N__3860),
            .I(N__3850));
    InMux I__778 (
            .O(N__3857),
            .I(N__3845));
    InMux I__777 (
            .O(N__3856),
            .I(N__3845));
    InMux I__776 (
            .O(N__3853),
            .I(N__3842));
    LocalMux I__775 (
            .O(N__3850),
            .I(beamYZ0Z_7));
    LocalMux I__774 (
            .O(N__3845),
            .I(beamYZ0Z_7));
    LocalMux I__773 (
            .O(N__3842),
            .I(beamYZ0Z_7));
    InMux I__772 (
            .O(N__3835),
            .I(N__3832));
    LocalMux I__771 (
            .O(N__3832),
            .I(N__3828));
    InMux I__770 (
            .O(N__3831),
            .I(N__3825));
    Span4Mux_h I__769 (
            .O(N__3828),
            .I(N__3822));
    LocalMux I__768 (
            .O(N__3825),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum));
    Odrv4 I__767 (
            .O(N__3822),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum));
    InMux I__766 (
            .O(N__3817),
            .I(un5_visibley_cry_6));
    CascadeMux I__765 (
            .O(N__3814),
            .I(N__3800));
    CascadeMux I__764 (
            .O(N__3813),
            .I(N__3797));
    CascadeMux I__763 (
            .O(N__3812),
            .I(N__3794));
    CascadeMux I__762 (
            .O(N__3811),
            .I(N__3790));
    InMux I__761 (
            .O(N__3810),
            .I(N__3781));
    InMux I__760 (
            .O(N__3809),
            .I(N__3781));
    InMux I__759 (
            .O(N__3808),
            .I(N__3781));
    InMux I__758 (
            .O(N__3807),
            .I(N__3778));
    InMux I__757 (
            .O(N__3806),
            .I(N__3773));
    InMux I__756 (
            .O(N__3805),
            .I(N__3773));
    InMux I__755 (
            .O(N__3804),
            .I(N__3770));
    InMux I__754 (
            .O(N__3803),
            .I(N__3767));
    InMux I__753 (
            .O(N__3800),
            .I(N__3764));
    InMux I__752 (
            .O(N__3797),
            .I(N__3757));
    InMux I__751 (
            .O(N__3794),
            .I(N__3757));
    InMux I__750 (
            .O(N__3793),
            .I(N__3757));
    InMux I__749 (
            .O(N__3790),
            .I(N__3754));
    IoInMux I__748 (
            .O(N__3789),
            .I(N__3751));
    CascadeMux I__747 (
            .O(N__3788),
            .I(N__3748));
    LocalMux I__746 (
            .O(N__3781),
            .I(N__3743));
    LocalMux I__745 (
            .O(N__3778),
            .I(N__3734));
    LocalMux I__744 (
            .O(N__3773),
            .I(N__3734));
    LocalMux I__743 (
            .O(N__3770),
            .I(N__3734));
    LocalMux I__742 (
            .O(N__3767),
            .I(N__3734));
    LocalMux I__741 (
            .O(N__3764),
            .I(N__3727));
    LocalMux I__740 (
            .O(N__3757),
            .I(N__3727));
    LocalMux I__739 (
            .O(N__3754),
            .I(N__3727));
    LocalMux I__738 (
            .O(N__3751),
            .I(N__3724));
    InMux I__737 (
            .O(N__3748),
            .I(N__3721));
    CascadeMux I__736 (
            .O(N__3747),
            .I(N__3718));
    CascadeMux I__735 (
            .O(N__3746),
            .I(N__3715));
    Span4Mux_v I__734 (
            .O(N__3743),
            .I(N__3708));
    Span4Mux_v I__733 (
            .O(N__3734),
            .I(N__3708));
    Span4Mux_s3_v I__732 (
            .O(N__3727),
            .I(N__3708));
    IoSpan4Mux I__731 (
            .O(N__3724),
            .I(N__3705));
    LocalMux I__730 (
            .O(N__3721),
            .I(N__3702));
    InMux I__729 (
            .O(N__3718),
            .I(N__3697));
    InMux I__728 (
            .O(N__3715),
            .I(N__3697));
    Odrv4 I__727 (
            .O(N__3708),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__726 (
            .O(N__3705),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__725 (
            .O(N__3702),
            .I(CONSTANT_ONE_NET));
    LocalMux I__724 (
            .O(N__3697),
            .I(CONSTANT_ONE_NET));
    InMux I__723 (
            .O(N__3688),
            .I(N__3682));
    CascadeMux I__722 (
            .O(N__3687),
            .I(N__3679));
    InMux I__721 (
            .O(N__3686),
            .I(N__3676));
    InMux I__720 (
            .O(N__3685),
            .I(N__3673));
    LocalMux I__719 (
            .O(N__3682),
            .I(N__3670));
    InMux I__718 (
            .O(N__3679),
            .I(N__3667));
    LocalMux I__717 (
            .O(N__3676),
            .I(beamYZ0Z_8));
    LocalMux I__716 (
            .O(N__3673),
            .I(beamYZ0Z_8));
    Odrv4 I__715 (
            .O(N__3670),
            .I(beamYZ0Z_8));
    LocalMux I__714 (
            .O(N__3667),
            .I(beamYZ0Z_8));
    InMux I__713 (
            .O(N__3658),
            .I(N__3652));
    InMux I__712 (
            .O(N__3657),
            .I(N__3652));
    LocalMux I__711 (
            .O(N__3652),
            .I(N__3649));
    Odrv4 I__710 (
            .O(N__3649),
            .I(un5_visibley_cry_7_c_RNI1L4CZ0));
    InMux I__709 (
            .O(N__3646),
            .I(bfn_9_8_0_));
    InMux I__708 (
            .O(N__3643),
            .I(N__3639));
    InMux I__707 (
            .O(N__3642),
            .I(N__3634));
    LocalMux I__706 (
            .O(N__3639),
            .I(N__3631));
    InMux I__705 (
            .O(N__3638),
            .I(N__3628));
    InMux I__704 (
            .O(N__3637),
            .I(N__3625));
    LocalMux I__703 (
            .O(N__3634),
            .I(beamYZ0Z_9));
    Odrv4 I__702 (
            .O(N__3631),
            .I(beamYZ0Z_9));
    LocalMux I__701 (
            .O(N__3628),
            .I(beamYZ0Z_9));
    LocalMux I__700 (
            .O(N__3625),
            .I(beamYZ0Z_9));
    InMux I__699 (
            .O(N__3616),
            .I(un5_visibley_cry_8));
    CascadeMux I__698 (
            .O(N__3613),
            .I(N__3610));
    InMux I__697 (
            .O(N__3610),
            .I(N__3604));
    InMux I__696 (
            .O(N__3609),
            .I(N__3604));
    LocalMux I__695 (
            .O(N__3604),
            .I(N__3601));
    Odrv4 I__694 (
            .O(N__3601),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_axb_3));
    CascadeMux I__693 (
            .O(N__3598),
            .I(N_8_cascade_));
    InMux I__692 (
            .O(N__3595),
            .I(N__3592));
    LocalMux I__691 (
            .O(N__3592),
            .I(N__3589));
    Odrv12 I__690 (
            .O(N__3589),
            .I(un1_beamX_27));
    InMux I__689 (
            .O(N__3586),
            .I(N__3583));
    LocalMux I__688 (
            .O(N__3583),
            .I(N__3580));
    Odrv4 I__687 (
            .O(N__3580),
            .I(Pixel_0_sqmuxa_1));
    CascadeMux I__686 (
            .O(N__3577),
            .I(un13_0_1_cascade_));
    InMux I__685 (
            .O(N__3574),
            .I(N__3571));
    LocalMux I__684 (
            .O(N__3571),
            .I(N__3568));
    Span4Mux_s2_v I__683 (
            .O(N__3568),
            .I(N__3565));
    Odrv4 I__682 (
            .O(N__3565),
            .I(un12lt10));
    IoInMux I__681 (
            .O(N__3562),
            .I(N__3559));
    LocalMux I__680 (
            .O(N__3559),
            .I(N__3556));
    Span4Mux_s3_v I__679 (
            .O(N__3556),
            .I(N__3552));
    IoInMux I__678 (
            .O(N__3555),
            .I(N__3549));
    Span4Mux_v I__677 (
            .O(N__3552),
            .I(N__3546));
    LocalMux I__676 (
            .O(N__3549),
            .I(N__3543));
    Span4Mux_v I__675 (
            .O(N__3546),
            .I(N__3540));
    Span4Mux_s1_v I__674 (
            .O(N__3543),
            .I(N__3537));
    Odrv4 I__673 (
            .O(N__3540),
            .I(Pixel_c));
    Odrv4 I__672 (
            .O(N__3537),
            .I(Pixel_c));
    ClkMux I__671 (
            .O(N__3532),
            .I(N__3508));
    ClkMux I__670 (
            .O(N__3531),
            .I(N__3508));
    ClkMux I__669 (
            .O(N__3530),
            .I(N__3508));
    ClkMux I__668 (
            .O(N__3529),
            .I(N__3508));
    ClkMux I__667 (
            .O(N__3528),
            .I(N__3508));
    ClkMux I__666 (
            .O(N__3527),
            .I(N__3508));
    ClkMux I__665 (
            .O(N__3526),
            .I(N__3508));
    ClkMux I__664 (
            .O(N__3525),
            .I(N__3508));
    GlobalMux I__663 (
            .O(N__3508),
            .I(N__3505));
    gio2CtrlBuf I__662 (
            .O(N__3505),
            .I(PixelClock_g));
    InMux I__661 (
            .O(N__3502),
            .I(N__3499));
    LocalMux I__660 (
            .O(N__3499),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__659 (
            .O(N__3496),
            .I(N__3490));
    InMux I__658 (
            .O(N__3495),
            .I(N__3487));
    InMux I__657 (
            .O(N__3494),
            .I(N__3484));
    InMux I__656 (
            .O(N__3493),
            .I(N__3481));
    LocalMux I__655 (
            .O(N__3490),
            .I(N__3476));
    LocalMux I__654 (
            .O(N__3487),
            .I(N__3476));
    LocalMux I__653 (
            .O(N__3484),
            .I(N__3473));
    LocalMux I__652 (
            .O(N__3481),
            .I(un13_beamx));
    Odrv4 I__651 (
            .O(N__3476),
            .I(un13_beamx));
    Odrv4 I__650 (
            .O(N__3473),
            .I(un13_beamx));
    CEMux I__649 (
            .O(N__3466),
            .I(N__3461));
    CEMux I__648 (
            .O(N__3465),
            .I(N__3458));
    CEMux I__647 (
            .O(N__3464),
            .I(N__3455));
    LocalMux I__646 (
            .O(N__3461),
            .I(N__3452));
    LocalMux I__645 (
            .O(N__3458),
            .I(N__3449));
    LocalMux I__644 (
            .O(N__3455),
            .I(N__3442));
    Span4Mux_v I__643 (
            .O(N__3452),
            .I(N__3437));
    Span4Mux_v I__642 (
            .O(N__3449),
            .I(N__3437));
    InMux I__641 (
            .O(N__3448),
            .I(N__3432));
    InMux I__640 (
            .O(N__3447),
            .I(N__3432));
    InMux I__639 (
            .O(N__3446),
            .I(N__3429));
    InMux I__638 (
            .O(N__3445),
            .I(N__3426));
    Span4Mux_v I__637 (
            .O(N__3442),
            .I(N__3423));
    Span4Mux_v I__636 (
            .O(N__3437),
            .I(N__3420));
    LocalMux I__635 (
            .O(N__3432),
            .I(beamX_RNIVEM1Z0Z_4));
    LocalMux I__634 (
            .O(N__3429),
            .I(beamX_RNIVEM1Z0Z_4));
    LocalMux I__633 (
            .O(N__3426),
            .I(beamX_RNIVEM1Z0Z_4));
    Odrv4 I__632 (
            .O(N__3423),
            .I(beamX_RNIVEM1Z0Z_4));
    Odrv4 I__631 (
            .O(N__3420),
            .I(beamX_RNIVEM1Z0Z_4));
    InMux I__630 (
            .O(N__3409),
            .I(N__3403));
    CascadeMux I__629 (
            .O(N__3408),
            .I(N__3399));
    InMux I__628 (
            .O(N__3407),
            .I(N__3394));
    InMux I__627 (
            .O(N__3406),
            .I(N__3394));
    LocalMux I__626 (
            .O(N__3403),
            .I(N__3391));
    InMux I__625 (
            .O(N__3402),
            .I(N__3388));
    InMux I__624 (
            .O(N__3399),
            .I(N__3385));
    LocalMux I__623 (
            .O(N__3394),
            .I(beamYZ0Z_0));
    Odrv4 I__622 (
            .O(N__3391),
            .I(beamYZ0Z_0));
    LocalMux I__621 (
            .O(N__3388),
            .I(beamYZ0Z_0));
    LocalMux I__620 (
            .O(N__3385),
            .I(beamYZ0Z_0));
    CascadeMux I__619 (
            .O(N__3376),
            .I(N__3371));
    InMux I__618 (
            .O(N__3375),
            .I(N__3368));
    CascadeMux I__617 (
            .O(N__3374),
            .I(N__3363));
    InMux I__616 (
            .O(N__3371),
            .I(N__3360));
    LocalMux I__615 (
            .O(N__3368),
            .I(N__3357));
    CascadeMux I__614 (
            .O(N__3367),
            .I(N__3354));
    InMux I__613 (
            .O(N__3366),
            .I(N__3351));
    InMux I__612 (
            .O(N__3363),
            .I(N__3348));
    LocalMux I__611 (
            .O(N__3360),
            .I(N__3343));
    Span4Mux_v I__610 (
            .O(N__3357),
            .I(N__3343));
    InMux I__609 (
            .O(N__3354),
            .I(N__3340));
    LocalMux I__608 (
            .O(N__3351),
            .I(beamYZ0Z_1));
    LocalMux I__607 (
            .O(N__3348),
            .I(beamYZ0Z_1));
    Odrv4 I__606 (
            .O(N__3343),
            .I(beamYZ0Z_1));
    LocalMux I__605 (
            .O(N__3340),
            .I(beamYZ0Z_1));
    InMux I__604 (
            .O(N__3331),
            .I(un5_visibley_cry_0));
    CascadeMux I__603 (
            .O(N__3328),
            .I(N__3322));
    InMux I__602 (
            .O(N__3327),
            .I(N__3319));
    InMux I__601 (
            .O(N__3326),
            .I(N__3314));
    InMux I__600 (
            .O(N__3325),
            .I(N__3314));
    InMux I__599 (
            .O(N__3322),
            .I(N__3311));
    LocalMux I__598 (
            .O(N__3319),
            .I(beamYZ0Z_2));
    LocalMux I__597 (
            .O(N__3314),
            .I(beamYZ0Z_2));
    LocalMux I__596 (
            .O(N__3311),
            .I(beamYZ0Z_2));
    InMux I__595 (
            .O(N__3304),
            .I(un5_visibley_cry_1));
    CascadeMux I__594 (
            .O(N__3301),
            .I(N__3295));
    InMux I__593 (
            .O(N__3300),
            .I(N__3292));
    InMux I__592 (
            .O(N__3299),
            .I(N__3287));
    InMux I__591 (
            .O(N__3298),
            .I(N__3287));
    InMux I__590 (
            .O(N__3295),
            .I(N__3284));
    LocalMux I__589 (
            .O(N__3292),
            .I(beamYZ0Z_3));
    LocalMux I__588 (
            .O(N__3287),
            .I(beamYZ0Z_3));
    LocalMux I__587 (
            .O(N__3284),
            .I(beamYZ0Z_3));
    InMux I__586 (
            .O(N__3277),
            .I(un5_visibley_cry_2));
    CascadeMux I__585 (
            .O(N__3274),
            .I(N__3268));
    InMux I__584 (
            .O(N__3273),
            .I(N__3265));
    InMux I__583 (
            .O(N__3272),
            .I(N__3262));
    InMux I__582 (
            .O(N__3271),
            .I(N__3259));
    InMux I__581 (
            .O(N__3268),
            .I(N__3256));
    LocalMux I__580 (
            .O(N__3265),
            .I(beamYZ0Z_4));
    LocalMux I__579 (
            .O(N__3262),
            .I(beamYZ0Z_4));
    LocalMux I__578 (
            .O(N__3259),
            .I(beamYZ0Z_4));
    LocalMux I__577 (
            .O(N__3256),
            .I(beamYZ0Z_4));
    InMux I__576 (
            .O(N__3247),
            .I(un5_visibley_cry_3));
    CascadeMux I__575 (
            .O(N__3244),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_));
    InMux I__574 (
            .O(N__3241),
            .I(N__3238));
    LocalMux I__573 (
            .O(N__3238),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__572 (
            .O(N__3235),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__571 (
            .O(N__3232),
            .I(N__3229));
    InMux I__570 (
            .O(N__3229),
            .I(N__3226));
    LocalMux I__569 (
            .O(N__3226),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1));
    InMux I__568 (
            .O(N__3223),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__567 (
            .O(N__3220),
            .I(N__3217));
    LocalMux I__566 (
            .O(N__3217),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1));
    InMux I__565 (
            .O(N__3214),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__564 (
            .O(N__3211),
            .I(N__3208));
    LocalMux I__563 (
            .O(N__3208),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1));
    InMux I__562 (
            .O(N__3205),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__561 (
            .O(N__3202),
            .I(N__3199));
    LocalMux I__560 (
            .O(N__3199),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__559 (
            .O(N__3196),
            .I(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__558 (
            .O(N__3193),
            .I(N__3188));
    CascadeMux I__557 (
            .O(N__3192),
            .I(N__3184));
    InMux I__556 (
            .O(N__3191),
            .I(N__3180));
    InMux I__555 (
            .O(N__3188),
            .I(N__3171));
    InMux I__554 (
            .O(N__3187),
            .I(N__3171));
    InMux I__553 (
            .O(N__3184),
            .I(N__3171));
    InMux I__552 (
            .O(N__3183),
            .I(N__3171));
    LocalMux I__551 (
            .O(N__3180),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1));
    LocalMux I__550 (
            .O(N__3171),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1));
    CascadeMux I__549 (
            .O(N__3166),
            .I(N__3163));
    InMux I__548 (
            .O(N__3163),
            .I(N__3160));
    LocalMux I__547 (
            .O(N__3160),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__546 (
            .O(N__3157),
            .I(N__3152));
    InMux I__545 (
            .O(N__3156),
            .I(N__3147));
    InMux I__544 (
            .O(N__3155),
            .I(N__3140));
    InMux I__543 (
            .O(N__3152),
            .I(N__3140));
    InMux I__542 (
            .O(N__3151),
            .I(N__3140));
    InMux I__541 (
            .O(N__3150),
            .I(N__3137));
    LocalMux I__540 (
            .O(N__3147),
            .I(beamXZ0Z_9));
    LocalMux I__539 (
            .O(N__3140),
            .I(beamXZ0Z_9));
    LocalMux I__538 (
            .O(N__3137),
            .I(beamXZ0Z_9));
    CascadeMux I__537 (
            .O(N__3130),
            .I(N__3123));
    InMux I__536 (
            .O(N__3129),
            .I(N__3119));
    InMux I__535 (
            .O(N__3128),
            .I(N__3116));
    InMux I__534 (
            .O(N__3127),
            .I(N__3109));
    InMux I__533 (
            .O(N__3126),
            .I(N__3109));
    InMux I__532 (
            .O(N__3123),
            .I(N__3109));
    InMux I__531 (
            .O(N__3122),
            .I(N__3106));
    LocalMux I__530 (
            .O(N__3119),
            .I(beamXZ0Z_7));
    LocalMux I__529 (
            .O(N__3116),
            .I(beamXZ0Z_7));
    LocalMux I__528 (
            .O(N__3109),
            .I(beamXZ0Z_7));
    LocalMux I__527 (
            .O(N__3106),
            .I(beamXZ0Z_7));
    InMux I__526 (
            .O(N__3097),
            .I(N__3089));
    InMux I__525 (
            .O(N__3096),
            .I(N__3084));
    InMux I__524 (
            .O(N__3095),
            .I(N__3084));
    InMux I__523 (
            .O(N__3094),
            .I(N__3079));
    InMux I__522 (
            .O(N__3093),
            .I(N__3079));
    InMux I__521 (
            .O(N__3092),
            .I(N__3076));
    LocalMux I__520 (
            .O(N__3089),
            .I(beamXZ0Z_6));
    LocalMux I__519 (
            .O(N__3084),
            .I(beamXZ0Z_6));
    LocalMux I__518 (
            .O(N__3079),
            .I(beamXZ0Z_6));
    LocalMux I__517 (
            .O(N__3076),
            .I(beamXZ0Z_6));
    InMux I__516 (
            .O(N__3067),
            .I(N__3060));
    InMux I__515 (
            .O(N__3066),
            .I(N__3057));
    InMux I__514 (
            .O(N__3065),
            .I(N__3052));
    InMux I__513 (
            .O(N__3064),
            .I(N__3052));
    InMux I__512 (
            .O(N__3063),
            .I(N__3049));
    LocalMux I__511 (
            .O(N__3060),
            .I(beamXZ0Z_8));
    LocalMux I__510 (
            .O(N__3057),
            .I(beamXZ0Z_8));
    LocalMux I__509 (
            .O(N__3052),
            .I(beamXZ0Z_8));
    LocalMux I__508 (
            .O(N__3049),
            .I(beamXZ0Z_8));
    CascadeMux I__507 (
            .O(N__3040),
            .I(un1_beamxlto9_0_cascade_));
    InMux I__506 (
            .O(N__3037),
            .I(N__3029));
    InMux I__505 (
            .O(N__3036),
            .I(N__3024));
    InMux I__504 (
            .O(N__3035),
            .I(N__3024));
    InMux I__503 (
            .O(N__3034),
            .I(N__3019));
    InMux I__502 (
            .O(N__3033),
            .I(N__3019));
    InMux I__501 (
            .O(N__3032),
            .I(N__3016));
    LocalMux I__500 (
            .O(N__3029),
            .I(beamXZ0Z_5));
    LocalMux I__499 (
            .O(N__3024),
            .I(beamXZ0Z_5));
    LocalMux I__498 (
            .O(N__3019),
            .I(beamXZ0Z_5));
    LocalMux I__497 (
            .O(N__3016),
            .I(beamXZ0Z_5));
    IoInMux I__496 (
            .O(N__3007),
            .I(N__3004));
    LocalMux I__495 (
            .O(N__3004),
            .I(N__3001));
    Span4Mux_s2_v I__494 (
            .O(N__3001),
            .I(N__2998));
    Span4Mux_v I__493 (
            .O(N__2998),
            .I(N__2995));
    Span4Mux_v I__492 (
            .O(N__2995),
            .I(N__2991));
    IoInMux I__491 (
            .O(N__2994),
            .I(N__2988));
    Span4Mux_v I__490 (
            .O(N__2991),
            .I(N__2985));
    LocalMux I__489 (
            .O(N__2988),
            .I(N__2982));
    Odrv4 I__488 (
            .O(N__2985),
            .I(HSync_c));
    Odrv4 I__487 (
            .O(N__2982),
            .I(HSync_c));
    InMux I__486 (
            .O(N__2977),
            .I(N__2973));
    InMux I__485 (
            .O(N__2976),
            .I(N__2970));
    LocalMux I__484 (
            .O(N__2973),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__483 (
            .O(N__2970),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    InMux I__482 (
            .O(N__2965),
            .I(N__2962));
    LocalMux I__481 (
            .O(N__2962),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_c5_i));
    CascadeMux I__480 (
            .O(N__2959),
            .I(N__2956));
    InMux I__479 (
            .O(N__2956),
            .I(N__2953));
    LocalMux I__478 (
            .O(N__2953),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365));
    InMux I__477 (
            .O(N__2950),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__476 (
            .O(N__2947),
            .I(N__2944));
    InMux I__475 (
            .O(N__2944),
            .I(N__2941));
    LocalMux I__474 (
            .O(N__2941),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575));
    InMux I__473 (
            .O(N__2938),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5));
    CascadeMux I__472 (
            .O(N__2935),
            .I(N__2932));
    InMux I__471 (
            .O(N__2932),
            .I(N__2929));
    LocalMux I__470 (
            .O(N__2929),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO));
    InMux I__469 (
            .O(N__2926),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__468 (
            .O(N__2923),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__467 (
            .O(N__2920),
            .I(N__2915));
    InMux I__466 (
            .O(N__2919),
            .I(N__2910));
    InMux I__465 (
            .O(N__2918),
            .I(N__2910));
    LocalMux I__464 (
            .O(N__2915),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_c5));
    LocalMux I__463 (
            .O(N__2910),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_c5));
    InMux I__462 (
            .O(N__2905),
            .I(N__2902));
    LocalMux I__461 (
            .O(N__2902),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_0));
    InMux I__460 (
            .O(N__2899),
            .I(N__2895));
    InMux I__459 (
            .O(N__2898),
            .I(N__2892));
    LocalMux I__458 (
            .O(N__2895),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    LocalMux I__457 (
            .O(N__2892),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    InMux I__456 (
            .O(N__2887),
            .I(N__2883));
    InMux I__455 (
            .O(N__2886),
            .I(N__2880));
    LocalMux I__454 (
            .O(N__2883),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23));
    LocalMux I__453 (
            .O(N__2880),
            .I(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23));
    InMux I__452 (
            .O(N__2875),
            .I(un16_beamx_cry_4));
    InMux I__451 (
            .O(N__2872),
            .I(un16_beamx_cry_5));
    InMux I__450 (
            .O(N__2869),
            .I(un16_beamx_cry_6));
    InMux I__449 (
            .O(N__2866),
            .I(un16_beamx_cry_7));
    InMux I__448 (
            .O(N__2863),
            .I(bfn_9_2_0_));
    InMux I__447 (
            .O(N__2860),
            .I(N__2857));
    LocalMux I__446 (
            .O(N__2857),
            .I(N__2854));
    Span4Mux_s2_v I__445 (
            .O(N__2854),
            .I(N__2851));
    Span4Mux_v I__444 (
            .O(N__2851),
            .I(N__2848));
    Odrv4 I__443 (
            .O(N__2848),
            .I(un1_beamy));
    InMux I__442 (
            .O(N__2845),
            .I(N__2842));
    LocalMux I__441 (
            .O(N__2842),
            .I(un4_beamxlt9));
    CascadeMux I__440 (
            .O(N__2839),
            .I(Pixel_0_sqmuxa_0_cascade_));
    InMux I__439 (
            .O(N__2836),
            .I(N__2832));
    InMux I__438 (
            .O(N__2835),
            .I(N__2829));
    LocalMux I__437 (
            .O(N__2832),
            .I(un11_beamx_1));
    LocalMux I__436 (
            .O(N__2829),
            .I(un11_beamx_1));
    InMux I__435 (
            .O(N__2824),
            .I(N__2816));
    InMux I__434 (
            .O(N__2823),
            .I(N__2811));
    InMux I__433 (
            .O(N__2822),
            .I(N__2811));
    InMux I__432 (
            .O(N__2821),
            .I(N__2808));
    InMux I__431 (
            .O(N__2820),
            .I(N__2803));
    InMux I__430 (
            .O(N__2819),
            .I(N__2803));
    LocalMux I__429 (
            .O(N__2816),
            .I(beamXZ0Z_4));
    LocalMux I__428 (
            .O(N__2811),
            .I(beamXZ0Z_4));
    LocalMux I__427 (
            .O(N__2808),
            .I(beamXZ0Z_4));
    LocalMux I__426 (
            .O(N__2803),
            .I(beamXZ0Z_4));
    InMux I__425 (
            .O(N__2794),
            .I(N__2791));
    LocalMux I__424 (
            .O(N__2791),
            .I(un8_beamxlt9_0));
    InMux I__423 (
            .O(N__2788),
            .I(un4_beamy_cry_5));
    InMux I__422 (
            .O(N__2785),
            .I(un4_beamy_cry_6));
    InMux I__421 (
            .O(N__2782),
            .I(un4_beamy_cry_7));
    InMux I__420 (
            .O(N__2779),
            .I(bfn_8_8_0_));
    InMux I__419 (
            .O(N__2776),
            .I(N__2770));
    InMux I__418 (
            .O(N__2775),
            .I(N__2763));
    InMux I__417 (
            .O(N__2774),
            .I(N__2763));
    InMux I__416 (
            .O(N__2773),
            .I(N__2763));
    LocalMux I__415 (
            .O(N__2770),
            .I(beamXZ0Z_0));
    LocalMux I__414 (
            .O(N__2763),
            .I(beamXZ0Z_0));
    CascadeMux I__413 (
            .O(N__2758),
            .I(N__2755));
    InMux I__412 (
            .O(N__2755),
            .I(N__2750));
    InMux I__411 (
            .O(N__2754),
            .I(N__2745));
    InMux I__410 (
            .O(N__2753),
            .I(N__2745));
    LocalMux I__409 (
            .O(N__2750),
            .I(beamXZ0Z_1));
    LocalMux I__408 (
            .O(N__2745),
            .I(beamXZ0Z_1));
    InMux I__407 (
            .O(N__2740),
            .I(N__2736));
    InMux I__406 (
            .O(N__2739),
            .I(N__2733));
    LocalMux I__405 (
            .O(N__2736),
            .I(beamXZ0Z_2));
    LocalMux I__404 (
            .O(N__2733),
            .I(beamXZ0Z_2));
    InMux I__403 (
            .O(N__2728),
            .I(un16_beamx_cry_1));
    InMux I__402 (
            .O(N__2725),
            .I(N__2722));
    LocalMux I__401 (
            .O(N__2722),
            .I(N__2718));
    CascadeMux I__400 (
            .O(N__2721),
            .I(N__2714));
    Span4Mux_v I__399 (
            .O(N__2718),
            .I(N__2711));
    InMux I__398 (
            .O(N__2717),
            .I(N__2708));
    InMux I__397 (
            .O(N__2714),
            .I(N__2705));
    Odrv4 I__396 (
            .O(N__2711),
            .I(beamXZ0Z_3));
    LocalMux I__395 (
            .O(N__2708),
            .I(beamXZ0Z_3));
    LocalMux I__394 (
            .O(N__2705),
            .I(beamXZ0Z_3));
    InMux I__393 (
            .O(N__2698),
            .I(un16_beamx_cry_2));
    InMux I__392 (
            .O(N__2695),
            .I(un16_beamx_cry_3));
    CascadeMux I__391 (
            .O(N__2692),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    CascadeMux I__390 (
            .O(N__2689),
            .I(N__2684));
    InMux I__389 (
            .O(N__2688),
            .I(N__2681));
    InMux I__388 (
            .O(N__2687),
            .I(N__2678));
    InMux I__387 (
            .O(N__2684),
            .I(N__2675));
    LocalMux I__386 (
            .O(N__2681),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__385 (
            .O(N__2678),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__384 (
            .O(N__2675),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_axb_6));
    InMux I__383 (
            .O(N__2668),
            .I(N__2665));
    LocalMux I__382 (
            .O(N__2665),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__381 (
            .O(N__2662),
            .I(N__2659));
    LocalMux I__380 (
            .O(N__2659),
            .I(un5_visibley_cry_7_c_RNI1L4CZ0Z_0));
    CascadeMux I__379 (
            .O(N__2656),
            .I(N__2653));
    InMux I__378 (
            .O(N__2653),
            .I(N__2650));
    LocalMux I__377 (
            .O(N__2650),
            .I(un5_visibley_cry_8_c_RNI3O5CZ0Z_0));
    InMux I__376 (
            .O(N__2647),
            .I(un4_beamy_cry_1));
    InMux I__375 (
            .O(N__2644),
            .I(un4_beamy_cry_2));
    InMux I__374 (
            .O(N__2641),
            .I(un4_beamy_cry_3));
    InMux I__373 (
            .O(N__2638),
            .I(un4_beamy_cry_4));
    InMux I__372 (
            .O(N__2635),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__371 (
            .O(N__2632),
            .I(N__2629));
    InMux I__370 (
            .O(N__2629),
            .I(N__2626));
    LocalMux I__369 (
            .O(N__2626),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0));
    InMux I__368 (
            .O(N__2623),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__367 (
            .O(N__2620),
            .I(N__2617));
    LocalMux I__366 (
            .O(N__2617),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0));
    InMux I__365 (
            .O(N__2614),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__364 (
            .O(N__2611),
            .I(N__2607));
    InMux I__363 (
            .O(N__2610),
            .I(N__2604));
    LocalMux I__362 (
            .O(N__2607),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0));
    LocalMux I__361 (
            .O(N__2604),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0));
    CascadeMux I__360 (
            .O(N__2599),
            .I(N__2596));
    InMux I__359 (
            .O(N__2596),
            .I(N__2593));
    LocalMux I__358 (
            .O(N__2593),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1));
    InMux I__357 (
            .O(N__2590),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__356 (
            .O(N__2587),
            .I(N__2584));
    LocalMux I__355 (
            .O(N__2584),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    CascadeMux I__354 (
            .O(N__2581),
            .I(N__2576));
    CascadeMux I__353 (
            .O(N__2580),
            .I(N__2573));
    CascadeMux I__352 (
            .O(N__2579),
            .I(N__2569));
    InMux I__351 (
            .O(N__2576),
            .I(N__2560));
    InMux I__350 (
            .O(N__2573),
            .I(N__2560));
    InMux I__349 (
            .O(N__2572),
            .I(N__2560));
    InMux I__348 (
            .O(N__2569),
            .I(N__2560));
    LocalMux I__347 (
            .O(N__2560),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0));
    InMux I__346 (
            .O(N__2557),
            .I(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__345 (
            .O(N__2554),
            .I(N__2551));
    LocalMux I__344 (
            .O(N__2551),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0));
    InMux I__343 (
            .O(N__2548),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__342 (
            .O(N__2545),
            .I(N__2542));
    LocalMux I__341 (
            .O(N__2542),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0));
    InMux I__340 (
            .O(N__2539),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__339 (
            .O(N__2536),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__338 (
            .O(N__2533),
            .I(N__2530));
    LocalMux I__337 (
            .O(N__2530),
            .I(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__336 (
            .O(N__2527),
            .I(N__2524));
    LocalMux I__335 (
            .O(N__2524),
            .I(N__2520));
    InMux I__334 (
            .O(N__2523),
            .I(N__2517));
    Span4Mux_v I__333 (
            .O(N__2520),
            .I(N__2514));
    LocalMux I__332 (
            .O(N__2517),
            .I(N__2511));
    Odrv4 I__331 (
            .O(N__2514),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum));
    Odrv4 I__330 (
            .O(N__2511),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum));
    InMux I__329 (
            .O(N__2506),
            .I(N__2503));
    LocalMux I__328 (
            .O(N__2503),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__327 (
            .O(N__2500),
            .I(N__2497));
    InMux I__326 (
            .O(N__2497),
            .I(N__2494));
    LocalMux I__325 (
            .O(N__2494),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__324 (
            .O(N__2491),
            .I(N__2488));
    InMux I__323 (
            .O(N__2488),
            .I(N__2485));
    LocalMux I__322 (
            .O(N__2485),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731));
    InMux I__321 (
            .O(N__2482),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__320 (
            .O(N__2479),
            .I(N__2476));
    LocalMux I__319 (
            .O(N__2476),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0));
    CascadeMux I__318 (
            .O(N__2473),
            .I(N__2470));
    InMux I__317 (
            .O(N__2470),
            .I(N__2467));
    LocalMux I__316 (
            .O(N__2467),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1));
    InMux I__315 (
            .O(N__2464),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__314 (
            .O(N__2461),
            .I(N__2458));
    LocalMux I__313 (
            .O(N__2458),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__312 (
            .O(N__2455),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__311 (
            .O(N__2452),
            .I(N__2449));
    LocalMux I__310 (
            .O(N__2449),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__309 (
            .O(N__2446),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__308 (
            .O(N__2443),
            .I(N__2439));
    InMux I__307 (
            .O(N__2442),
            .I(N__2436));
    LocalMux I__306 (
            .O(N__2439),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1));
    LocalMux I__305 (
            .O(N__2436),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1));
    CascadeMux I__304 (
            .O(N__2431),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_));
    InMux I__303 (
            .O(N__2428),
            .I(N__2422));
    InMux I__302 (
            .O(N__2427),
            .I(N__2422));
    LocalMux I__301 (
            .O(N__2422),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__300 (
            .O(N__2419),
            .I(N__2415));
    InMux I__299 (
            .O(N__2418),
            .I(N__2410));
    InMux I__298 (
            .O(N__2415),
            .I(N__2410));
    LocalMux I__297 (
            .O(N__2410),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0));
    CascadeMux I__296 (
            .O(N__2407),
            .I(N__2403));
    InMux I__295 (
            .O(N__2406),
            .I(N__2399));
    InMux I__294 (
            .O(N__2403),
            .I(N__2394));
    InMux I__293 (
            .O(N__2402),
            .I(N__2394));
    LocalMux I__292 (
            .O(N__2399),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0));
    LocalMux I__291 (
            .O(N__2394),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0));
    InMux I__290 (
            .O(N__2389),
            .I(N__2386));
    LocalMux I__289 (
            .O(N__2386),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631));
    CascadeMux I__288 (
            .O(N__2383),
            .I(N__2379));
    InMux I__287 (
            .O(N__2382),
            .I(N__2374));
    InMux I__286 (
            .O(N__2379),
            .I(N__2371));
    InMux I__285 (
            .O(N__2378),
            .I(N__2366));
    InMux I__284 (
            .O(N__2377),
            .I(N__2366));
    LocalMux I__283 (
            .O(N__2374),
            .I(un5_visiblex_i));
    LocalMux I__282 (
            .O(N__2371),
            .I(un5_visiblex_i));
    LocalMux I__281 (
            .O(N__2366),
            .I(un5_visiblex_i));
    InMux I__280 (
            .O(N__2359),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__279 (
            .O(N__2356),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__278 (
            .O(N__2353),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__277 (
            .O(N__2350),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__276 (
            .O(N__2347),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_));
    InMux I__275 (
            .O(N__2344),
            .I(N__2338));
    InMux I__274 (
            .O(N__2343),
            .I(N__2338));
    LocalMux I__273 (
            .O(N__2338),
            .I(un1_beamX_if_generate_plus_mult1_un54_sum));
    CascadeMux I__272 (
            .O(N__2335),
            .I(N__2332));
    InMux I__271 (
            .O(N__2332),
            .I(N__2329));
    LocalMux I__270 (
            .O(N__2329),
            .I(un5_visiblex_i_24));
    CascadeMux I__269 (
            .O(N__2326),
            .I(N__2323));
    InMux I__268 (
            .O(N__2323),
            .I(N__2319));
    InMux I__267 (
            .O(N__2322),
            .I(N__2316));
    LocalMux I__266 (
            .O(N__2319),
            .I(N__2313));
    LocalMux I__265 (
            .O(N__2316),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum));
    Odrv4 I__264 (
            .O(N__2313),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum));
    InMux I__263 (
            .O(N__2308),
            .I(un5_visiblex_cry_4));
    InMux I__262 (
            .O(N__2305),
            .I(un5_visiblex_cry_5));
    InMux I__261 (
            .O(N__2302),
            .I(un5_visiblex_cry_6));
    InMux I__260 (
            .O(N__2299),
            .I(un5_visiblex_cry_7));
    InMux I__259 (
            .O(N__2296),
            .I(un5_visiblex_cry_8));
    CascadeMux I__258 (
            .O(N__2293),
            .I(un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_));
    CascadeMux I__257 (
            .O(N__2290),
            .I(un13_beamx_6_cascade_));
    InMux I__256 (
            .O(N__2287),
            .I(N__2284));
    LocalMux I__255 (
            .O(N__2284),
            .I(un13_beamx_5));
    InMux I__254 (
            .O(N__2281),
            .I(N__2278));
    LocalMux I__253 (
            .O(N__2278),
            .I(un1_beamylto9_4));
    CascadeMux I__252 (
            .O(N__2275),
            .I(un1_beamylto9_5_cascade_));
    CascadeMux I__251 (
            .O(N__2272),
            .I(un1_beamy_cascade_));
    IoInMux I__250 (
            .O(N__2269),
            .I(N__2266));
    LocalMux I__249 (
            .O(N__2266),
            .I(N__2263));
    Span4Mux_s2_v I__248 (
            .O(N__2263),
            .I(N__2259));
    IoInMux I__247 (
            .O(N__2262),
            .I(N__2256));
    Span4Mux_h I__246 (
            .O(N__2259),
            .I(N__2253));
    LocalMux I__245 (
            .O(N__2256),
            .I(N__2250));
    Span4Mux_v I__244 (
            .O(N__2253),
            .I(N__2247));
    Span4Mux_s2_v I__243 (
            .O(N__2250),
            .I(N__2244));
    Odrv4 I__242 (
            .O(N__2247),
            .I(VSync_c));
    Odrv4 I__241 (
            .O(N__2244),
            .I(VSync_c));
    CascadeMux I__240 (
            .O(N__2239),
            .I(un11_beamx_3_cascade_));
    InMux I__239 (
            .O(N__2236),
            .I(N__2233));
    LocalMux I__238 (
            .O(N__2233),
            .I(un11_beamx_6));
    CascadeMux I__237 (
            .O(N__2230),
            .I(un11_beamx_6_cascade_));
    CascadeMux I__236 (
            .O(N__2227),
            .I(N__2224));
    InMux I__235 (
            .O(N__2224),
            .I(N__2221));
    LocalMux I__234 (
            .O(N__2221),
            .I(un1_beamX_if_generate_plus_mult1_un61_sum_i));
    InMux I__233 (
            .O(N__2218),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__232 (
            .O(N__2215),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__231 (
            .O(N__2212),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__230 (
            .O(N__2209),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__229 (
            .O(N__2206),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__228 (
            .O(N__2203),
            .I(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_));
    InMux I__227 (
            .O(N__2200),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__226 (
            .O(N__2197),
            .I(N__2194));
    LocalMux I__225 (
            .O(N__2194),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57));
    CascadeMux I__224 (
            .O(N__2191),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_));
    InMux I__223 (
            .O(N__2188),
            .I(N__2184));
    InMux I__222 (
            .O(N__2187),
            .I(N__2181));
    LocalMux I__221 (
            .O(N__2184),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0));
    LocalMux I__220 (
            .O(N__2181),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0));
    CascadeMux I__219 (
            .O(N__2176),
            .I(N__2173));
    InMux I__218 (
            .O(N__2173),
            .I(N__2170));
    LocalMux I__217 (
            .O(N__2170),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_i));
    InMux I__216 (
            .O(N__2167),
            .I(N__2164));
    LocalMux I__215 (
            .O(N__2164),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1));
    InMux I__214 (
            .O(N__2161),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__213 (
            .O(N__2158),
            .I(N__2155));
    InMux I__212 (
            .O(N__2155),
            .I(N__2152));
    LocalMux I__211 (
            .O(N__2152),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2));
    InMux I__210 (
            .O(N__2149),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__209 (
            .O(N__2146),
            .I(N__2143));
    LocalMux I__208 (
            .O(N__2143),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__207 (
            .O(N__2140),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__206 (
            .O(N__2137),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__205 (
            .O(N__2134),
            .I(N__2130));
    InMux I__204 (
            .O(N__2133),
            .I(N__2126));
    InMux I__203 (
            .O(N__2130),
            .I(N__2121));
    InMux I__202 (
            .O(N__2129),
            .I(N__2121));
    LocalMux I__201 (
            .O(N__2126),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3));
    LocalMux I__200 (
            .O(N__2121),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3));
    InMux I__199 (
            .O(N__2116),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__198 (
            .O(N__2113),
            .I(N__2110));
    LocalMux I__197 (
            .O(N__2110),
            .I(Pixel_1_RNOZ0Z_6));
    InMux I__196 (
            .O(N__2107),
            .I(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__195 (
            .O(N__2104),
            .I(N__2098));
    InMux I__194 (
            .O(N__2103),
            .I(N__2098));
    LocalMux I__193 (
            .O(N__2098),
            .I(un1_beamX_if_generate_plus_mult1_un68_sum_i_8));
    IoInMux I__192 (
            .O(N__2095),
            .I(N__2092));
    LocalMux I__191 (
            .O(N__2092),
            .I(N__2089));
    Span4Mux_s1_h I__190 (
            .O(N__2089),
            .I(N__2086));
    Span4Mux_h I__189 (
            .O(N__2086),
            .I(N__2083));
    Sp12to4 I__188 (
            .O(N__2083),
            .I(N__2080));
    Odrv12 I__187 (
            .O(N__2080),
            .I(\VGAClock.PixelClock ));
    IoInMux I__186 (
            .O(N__2077),
            .I(N__2074));
    LocalMux I__185 (
            .O(N__2074),
            .I(N__2071));
    IoSpan4Mux I__184 (
            .O(N__2071),
            .I(N__2068));
    Odrv4 I__183 (
            .O(N__2068),
            .I(Clock12MHz_c));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(un5_visibley_cry_7),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(un4_beamy_cry_8),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(un16_beamx_cry_8),
            .carryinitout(bfn_9_2_0_));
    ICE_GB \VGAClock.PLLOUTCORE_derived_clock_RNIE579  (
            .USERSIGNALTOGLOBALBUFFER(N__2095),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_4_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_4_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_1_LC_7_2_5.C_ON=1'b0;
    defparam Pixel_1_RNO_1_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_1_LC_7_2_5.LUT_INIT=16'b0011100111001100;
    LogicCell40 Pixel_1_RNO_1_LC_7_2_5 (
            .in0(N__2187),
            .in1(N__2113),
            .in2(N__2383),
            .in3(N__2197),
            .lcout(un1_beamX_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_3_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__2377),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_7_3_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_7_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__2103),
            .in2(N__2176),
            .in3(N__2116),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_6_LC_7_3_2.C_ON=1'b1;
    defparam Pixel_1_RNO_6_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_6_LC_7_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_6_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__2167),
            .in2(N__2134),
            .in3(N__2107),
            .lcout(Pixel_1_RNOZ0Z_6),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_3_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_3_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(N__2104),
            .in2(N__2158),
            .in3(N__2129),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCR57_LC_7_3_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCR57_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCR57_LC_7_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCR57_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__2146),
            .in2(_gnd_net_),
            .in3(N__2200),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57),
            .ltout(un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNIJCRZ0Z57_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_2_LC_7_3_5.C_ON=1'b0;
    defparam Pixel_1_RNO_2_LC_7_3_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_2_LC_7_3_5.LUT_INIT=16'b1010110101000000;
    LogicCell40 Pixel_1_RNO_2_LC_7_3_5 (
            .in0(N__2378),
            .in1(N__2725),
            .in2(N__2191),
            .in3(N__2188),
            .lcout(un12lt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_3_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_7_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2322),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_4_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2326),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRM1_LC_7_4_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRM1_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRM1_LC_7_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRM1_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__2427),
            .in2(N__2227),
            .in3(N__2161),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNI1QRMZ0Z1),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1O2_LC_7_4_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1O2_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1O2_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1O2_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__2443),
            .in2(N__2491),
            .in3(N__2149),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI3F1OZ0Z2),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIG1IT6_LC_7_4_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIG1IT6_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIG1IT6_LC_7_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIG1IT6_LC_7_4_3 (
            .in0(N__2133),
            .in1(N__2428),
            .in2(N__2473),
            .in3(N__2140),
            .lcout(un1_beamX_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3P3_LC_7_4_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3P3_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3P3_LC_7_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3P3_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(N__2461),
            .in2(_gnd_net_),
            .in3(N__2137),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIAG3PZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_7_4_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_7_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_7_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2527),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0 (
            .in0(_gnd_net_),
            .in1(N__3835),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6O_LC_7_5_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6O_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6O_LC_7_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6O_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(N__2662),
            .in2(N__3746),
            .in3(N__2218),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNIHN6OZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3U_LC_7_5_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3U_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3U_LC_7_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3U_LC_7_5_2 (
            .in0(_gnd_net_),
            .in1(N__2554),
            .in2(N__3788),
            .in3(N__2215),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNI6M3UZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5U_LC_7_5_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5U_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5U_LC_7_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5U_LC_7_5_3 (
            .in0(_gnd_net_),
            .in1(N__2545),
            .in2(N__3747),
            .in3(N__2212),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8Q5UZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2689),
            .in3(N__2209),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883I_LC_7_5_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883I_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883I_LC_7_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883I_LC_7_5_5 (
            .in0(_gnd_net_),
            .in1(N__2533),
            .in2(_gnd_net_),
            .in3(N__2206),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0),
            .ltout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNI883IZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29G1_LC_7_5_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29G1_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29G1_LC_7_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29G1_LC_7_5_6 (
            .in0(N__2611),
            .in1(_gnd_net_),
            .in2(N__2203),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG29GZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIB625_9_LC_7_6_0.C_ON=1'b0;
    defparam beamY_RNIB625_9_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIB625_9_LC_7_6_0.LUT_INIT=16'b0000000100000000;
    LogicCell40 beamY_RNIB625_9_LC_7_6_0 (
            .in0(N__3953),
            .in1(N__3272),
            .in2(N__3376),
            .in3(N__3643),
            .lcout(),
            .ltout(un13_beamx_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_0_LC_7_6_1.C_ON=1'b0;
    defparam beamY_RNI9DLC_0_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_0_LC_7_6_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamY_RNI9DLC_0_LC_7_6_1 (
            .in0(N__2287),
            .in1(N__3409),
            .in2(N__2290),
            .in3(N__3685),
            .lcout(un13_beamx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIA525_2_LC_7_7_1.C_ON=1'b0;
    defparam beamY_RNIA525_2_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIA525_2_LC_7_7_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamY_RNIA525_2_LC_7_7_1 (
            .in0(N__3326),
            .in1(N__3910),
            .in2(N__3862),
            .in3(N__3299),
            .lcout(un13_beamx_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJNP3_2_LC_7_7_2.C_ON=1'b0;
    defparam beamY_RNIJNP3_2_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIJNP3_2_LC_7_7_2.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_RNIJNP3_2_LC_7_7_2 (
            .in0(N__3688),
            .in1(N__3856),
            .in2(_gnd_net_),
            .in3(N__3325),
            .lcout(un1_beamylto9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_1_LC_7_7_3.C_ON=1'b0;
    defparam beamY_RNI6125_1_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_1_LC_7_7_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamY_RNI6125_1_LC_7_7_3 (
            .in0(N__3271),
            .in1(N__3298),
            .in2(N__3913),
            .in3(N__3375),
            .lcout(),
            .ltout(un1_beamylto9_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0DB_9_LC_7_7_4.C_ON=1'b0;
    defparam beamY_RNIJ0DB_9_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0DB_9_LC_7_7_4.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamY_RNIJ0DB_9_LC_7_7_4 (
            .in0(N__2281),
            .in1(N__3638),
            .in2(N__2275),
            .in3(N__3952),
            .lcout(un1_beamy),
            .ltout(un1_beamy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_7_7_5.C_ON=1'b0;
    defparam VSync_1_LC_7_7_5.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_7_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 VSync_1_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2272),
            .in3(_gnd_net_),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3525),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIG3M_5_LC_8_1_0.C_ON=1'b0;
    defparam beamX_RNIG3M_5_LC_8_1_0.SEQ_MODE=4'b0000;
    defparam beamX_RNIG3M_5_LC_8_1_0.LUT_INIT=16'b0000000010001000;
    LogicCell40 beamX_RNIG3M_5_LC_8_1_0 (
            .in0(N__3036),
            .in1(N__2835),
            .in2(_gnd_net_),
            .in3(N__3096),
            .lcout(),
            .ltout(un11_beamx_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_4_LC_8_1_1.C_ON=1'b0;
    defparam beamX_RNIVEM1_4_LC_8_1_1.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_4_LC_8_1_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNIVEM1_4_LC_8_1_1 (
            .in0(N__2236),
            .in1(N__3128),
            .in2(N__2239),
            .in3(N__2823),
            .lcout(beamX_RNIVEM1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_8_1_2.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_8_1_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_8_1_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNIQCL_1_LC_8_1_2 (
            .in0(N__2739),
            .in1(N__2753),
            .in2(N__2721),
            .in3(N__2773),
            .lcout(un11_beamx_6),
            .ltout(un11_beamx_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_5_LC_8_1_3.C_ON=1'b0;
    defparam Pixel_1_RNO_5_LC_8_1_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_5_LC_8_1_3.LUT_INIT=16'b0001000100010101;
    LogicCell40 Pixel_1_RNO_5_LC_8_1_3 (
            .in0(N__3095),
            .in1(N__3035),
            .in2(N__2230),
            .in3(N__2822),
            .lcout(un4_beamxlt9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_8_1_5.C_ON=1'b0;
    defparam beamX_0_LC_8_1_5.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_8_1_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 beamX_0_LC_8_1_5 (
            .in0(N__2774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3529),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_8_1_6.C_ON=1'b0;
    defparam beamX_1_LC_8_1_6.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_8_1_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_8_1_6 (
            .in0(_gnd_net_),
            .in1(N__2754),
            .in2(_gnd_net_),
            .in3(N__2775),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3529),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_LC_8_2_0.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_LC_8_2_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_LC_8_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_4_c_LC_8_2_0 (
            .in0(_gnd_net_),
            .in1(N__2819),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_8_2_1 (
            .in0(_gnd_net_),
            .in1(N__3032),
            .in2(N__3814),
            .in3(N__2308),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_8_2_2 (
            .in0(_gnd_net_),
            .in1(N__3092),
            .in2(N__3812),
            .in3(N__2305),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_2_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_8_2_3 (
            .in0(_gnd_net_),
            .in1(N__3122),
            .in2(_gnd_net_),
            .in3(N__2302),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_2_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_8_2_4 (
            .in0(_gnd_net_),
            .in1(N__3063),
            .in2(N__3813),
            .in3(N__2299),
            .lcout(un5_visiblex_cry_7_c_RNIVZ0Z952),
            .ltout(),
            .carryin(un5_visiblex_cry_7),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5 (
            .in0(_gnd_net_),
            .in1(N__3150),
            .in2(_gnd_net_),
            .in3(N__2296),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_c5),
            .ltout(un1_beamX_if_generate_plus_mult1_un40_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_2_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_2_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_2_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_8_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2293),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un40_sum_c5_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_2_7.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_2_7.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_2_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_2_7 (
            .in0(N__2820),
            .in1(N__3793),
            .in2(_gnd_net_),
            .in3(N__2382),
            .lcout(un5_visiblex_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_3_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__2343),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_3_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(N__2899),
            .in2(N__2335),
            .in3(N__2359),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_3_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(N__2886),
            .in2(N__2959),
            .in3(N__2356),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6C831_LC_8_3_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6C831_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6C831_LC_8_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI6C831_LC_8_3_3 (
            .in0(N__2406),
            .in1(N__3241),
            .in2(N__2947),
            .in3(N__2353),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_LC_8_3_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_LC_8_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_LC_8_3_4 (
            .in0(N__2887),
            .in1(N__2920),
            .in2(N__2935),
            .in3(N__2350),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0),
            .ltout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LHZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_0_LC_8_3_5.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_0_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_0_LC_8_3_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNI48LH_0_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2347),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_3_6.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_8_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2344),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_3_7.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_8_3_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_8_3_7 (
            .in0(N__2977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_4_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__2523),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISM731_LC_8_4_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISM731_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISM731_LC_8_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISM731_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__2506),
            .in2(N__2500),
            .in3(N__2482),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNISMZ0Z731),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJF1_LC_8_4_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJF1_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJF1_LC_8_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJF1_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__2479),
            .in2(N__2407),
            .in3(N__2464),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNIUMJFZ0Z1),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5E1N3_LC_8_4_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5E1N3_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5E1N3_LC_8_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNI5E1N3_LC_8_4_3 (
            .in0(N__2442),
            .in1(N__2389),
            .in2(N__2419),
            .in3(N__2455),
            .lcout(un1_beamX_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_LC_8_4_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_LC_8_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_LC_8_4_4 (
            .in0(_gnd_net_),
            .in1(N__2452),
            .in2(_gnd_net_),
            .in3(N__2446),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1),
            .ltout(un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPIZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_0_LC_8_4_5.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_0_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_0_LC_8_4_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI4QPI1_0_LC_8_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2431),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI48631_LC_8_4_7.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI48631_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI48631_LC_8_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI48631_LC_8_4_7 (
            .in0(N__2418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2402),
            .lcout(un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNIZ0Z48631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_5_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453A1_LC_8_5_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453A1_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453A1_LC_8_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453A1_LC_8_5_1 (
            .in0(_gnd_net_),
            .in1(N__2668),
            .in2(N__2579),
            .in3(N__2635),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNI453AZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTO1_LC_8_5_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTO1_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTO1_LC_8_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTO1_LC_8_5_2 (
            .in0(_gnd_net_),
            .in1(N__2572),
            .in2(N__2632),
            .in3(N__2623),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNIHOTOZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRU1_LC_8_5_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRU1_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRU1_LC_8_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRU1_LC_8_5_3 (
            .in0(_gnd_net_),
            .in1(N__2620),
            .in2(N__2580),
            .in3(N__2614),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7PRUZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNI894A4_LC_8_5_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNI894A4_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNI894A4_LC_8_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNI894A4_LC_8_5_4 (
            .in0(N__3191),
            .in1(N__2610),
            .in2(N__2599),
            .in3(N__2590),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_LC_8_5_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_LC_8_5_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_LC_8_5_5 (
            .in0(N__2587),
            .in1(N__2687),
            .in2(N__2581),
            .in3(N__2557),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVCZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_6_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__3657),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_8_6_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_8_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__3803),
            .in2(N__2656),
            .in3(N__2548),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_8_6_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_8_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(N__3804),
            .in2(N__3613),
            .in3(N__2539),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_6_3.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_8_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2536),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_6_4.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_6_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2692),
            .in3(N__2688),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_6_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3831),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_8_6_6.C_ON=1'b0;
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_8_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visibley_cry_7_c_RNI1L4C_0_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3658),
            .lcout(un5_visibley_cry_7_c_RNI1L4CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_8_6_7.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_8_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_0_LC_8_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3609),
            .lcout(un5_visibley_cry_8_c_RNI3O5CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_beamy_cry_1_c_LC_8_7_0.C_ON=1'b1;
    defparam un4_beamy_cry_1_c_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un4_beamy_cry_1_c_LC_8_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_beamy_cry_1_c_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(N__3402),
            .in2(N__3374),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(un4_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_8_7_1.C_ON=1'b1;
    defparam beamY_2_LC_8_7_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_8_7_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_2_LC_8_7_1 (
            .in0(N__3493),
            .in1(N__3327),
            .in2(_gnd_net_),
            .in3(N__2647),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(un4_beamy_cry_1),
            .carryout(un4_beamy_cry_2),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_3_LC_8_7_2.C_ON=1'b1;
    defparam beamY_3_LC_8_7_2.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_8_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_3_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__3300),
            .in2(_gnd_net_),
            .in3(N__2644),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(un4_beamy_cry_2),
            .carryout(un4_beamy_cry_3),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_4_LC_8_7_3.C_ON=1'b1;
    defparam beamY_4_LC_8_7_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_8_7_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_4_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(N__3273),
            .in2(_gnd_net_),
            .in3(N__2641),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un4_beamy_cry_3),
            .carryout(un4_beamy_cry_4),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_5_LC_8_7_4.C_ON=1'b1;
    defparam beamY_5_LC_8_7_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_8_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_8_7_4 (
            .in0(_gnd_net_),
            .in1(N__3954),
            .in2(_gnd_net_),
            .in3(N__2638),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un4_beamy_cry_4),
            .carryout(un4_beamy_cry_5),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_6_LC_8_7_5.C_ON=1'b1;
    defparam beamY_6_LC_8_7_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_8_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(N__3911),
            .in2(_gnd_net_),
            .in3(N__2788),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un4_beamy_cry_5),
            .carryout(un4_beamy_cry_6),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_7_LC_8_7_6.C_ON=1'b1;
    defparam beamY_7_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_8_7_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_7_LC_8_7_6 (
            .in0(N__3496),
            .in1(N__3860),
            .in2(_gnd_net_),
            .in3(N__2785),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(un4_beamy_cry_6),
            .carryout(un4_beamy_cry_7),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_8_LC_8_7_7.C_ON=1'b1;
    defparam beamY_8_LC_8_7_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_8_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_8_7_7 (
            .in0(_gnd_net_),
            .in1(N__3686),
            .in2(_gnd_net_),
            .in3(N__2782),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un4_beamy_cry_7),
            .carryout(un4_beamy_cry_8),
            .clk(N__3527),
            .ce(N__3466),
            .sr(_gnd_net_));
    defparam beamY_9_LC_8_8_0.C_ON=1'b0;
    defparam beamY_9_LC_8_8_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_8_8_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_8_8_0 (
            .in0(N__3642),
            .in1(N__3495),
            .in2(_gnd_net_),
            .in3(N__2779),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3526),
            .ce(N__3465),
            .sr(_gnd_net_));
    defparam un16_beamx_cry_1_c_LC_9_1_0.C_ON=1'b1;
    defparam un16_beamx_cry_1_c_LC_9_1_0.SEQ_MODE=4'b0000;
    defparam un16_beamx_cry_1_c_LC_9_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un16_beamx_cry_1_c_LC_9_1_0 (
            .in0(_gnd_net_),
            .in1(N__2776),
            .in2(N__2758),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(un16_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_9_1_1.C_ON=1'b1;
    defparam beamX_2_LC_9_1_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_9_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_9_1_1 (
            .in0(_gnd_net_),
            .in1(N__2740),
            .in2(_gnd_net_),
            .in3(N__2728),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un16_beamx_cry_1),
            .carryout(un16_beamx_cry_2),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_9_1_2.C_ON=1'b1;
    defparam beamX_3_LC_9_1_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_9_1_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(N__2717),
            .in2(_gnd_net_),
            .in3(N__2698),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un16_beamx_cry_2),
            .carryout(un16_beamx_cry_3),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_9_1_3.C_ON=1'b1;
    defparam beamX_4_LC_9_1_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_9_1_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_4_LC_9_1_3 (
            .in0(_gnd_net_),
            .in1(N__2824),
            .in2(_gnd_net_),
            .in3(N__2695),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un16_beamx_cry_3),
            .carryout(un16_beamx_cry_4),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_9_1_4.C_ON=1'b1;
    defparam beamX_5_LC_9_1_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_9_1_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_9_1_4 (
            .in0(_gnd_net_),
            .in1(N__3037),
            .in2(_gnd_net_),
            .in3(N__2875),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un16_beamx_cry_4),
            .carryout(un16_beamx_cry_5),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_9_1_5.C_ON=1'b1;
    defparam beamX_6_LC_9_1_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_9_1_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_6_LC_9_1_5 (
            .in0(N__3447),
            .in1(N__3097),
            .in2(_gnd_net_),
            .in3(N__2872),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un16_beamx_cry_5),
            .carryout(un16_beamx_cry_6),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_9_1_6.C_ON=1'b1;
    defparam beamX_7_LC_9_1_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_9_1_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_7_LC_9_1_6 (
            .in0(N__3445),
            .in1(N__3129),
            .in2(_gnd_net_),
            .in3(N__2869),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un16_beamx_cry_6),
            .carryout(un16_beamx_cry_7),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_9_1_7.C_ON=1'b1;
    defparam beamX_8_LC_9_1_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_9_1_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_8_LC_9_1_7 (
            .in0(N__3448),
            .in1(N__3066),
            .in2(_gnd_net_),
            .in3(N__2866),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un16_beamx_cry_7),
            .carryout(un16_beamx_cry_8),
            .clk(N__3531),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_9_2_0.C_ON=1'b0;
    defparam beamX_9_LC_9_2_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_9_2_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_9_LC_9_2_0 (
            .in0(N__3156),
            .in1(N__3446),
            .in2(_gnd_net_),
            .in3(N__2863),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3530),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_4_LC_9_2_1.C_ON=1'b0;
    defparam Pixel_1_RNO_4_LC_9_2_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_4_LC_9_2_1.LUT_INIT=16'b0000000011111110;
    LogicCell40 Pixel_1_RNO_4_LC_9_2_1 (
            .in0(N__3065),
            .in1(N__2794),
            .in2(N__3157),
            .in3(N__2860),
            .lcout(),
            .ltout(Pixel_0_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_0_LC_9_2_2.C_ON=1'b0;
    defparam Pixel_1_RNO_0_LC_9_2_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_0_LC_9_2_2.LUT_INIT=16'b1011000011110000;
    LogicCell40 Pixel_1_RNO_0_LC_9_2_2 (
            .in0(N__2845),
            .in1(N__2836),
            .in2(N__2839),
            .in3(N__3126),
            .lcout(Pixel_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_9_2_4.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_9_2_4.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_9_2_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamX_RNIR4B_9_LC_9_2_4 (
            .in0(_gnd_net_),
            .in1(N__3151),
            .in2(_gnd_net_),
            .in3(N__3064),
            .lcout(un11_beamx_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_10_LC_9_2_5.C_ON=1'b0;
    defparam Pixel_1_RNO_10_LC_9_2_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_10_LC_9_2_5.LUT_INIT=16'b1111000011100000;
    LogicCell40 Pixel_1_RNO_10_LC_9_2_5 (
            .in0(N__3093),
            .in1(N__3033),
            .in2(N__3130),
            .in3(N__2821),
            .lcout(un8_beamxlt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_RNO_0_LC_9_2_6.C_ON=1'b0;
    defparam HSync_1_RNO_0_LC_9_2_6.SEQ_MODE=4'b0000;
    defparam HSync_1_RNO_0_LC_9_2_6.LUT_INIT=16'b0000000000110011;
    LogicCell40 HSync_1_RNO_0_LC_9_2_6 (
            .in0(_gnd_net_),
            .in1(N__3155),
            .in2(_gnd_net_),
            .in3(N__3127),
            .lcout(),
            .ltout(un1_beamxlto9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_9_2_7.C_ON=1'b0;
    defparam HSync_1_LC_9_2_7.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_9_2_7.LUT_INIT=16'b1110111111001111;
    LogicCell40 HSync_1_LC_9_2_7 (
            .in0(N__3094),
            .in1(N__3067),
            .in2(N__3040),
            .in3(N__3034),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3530),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_3_0.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_9_3_0 (
            .in0(_gnd_net_),
            .in1(N__2976),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_9_3_1.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_9_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_9_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_9_3_1 (
            .in0(_gnd_net_),
            .in1(N__2965),
            .in2(_gnd_net_),
            .in3(N__2950),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNI1575_LC_9_3_2.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNI1575_LC_9_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNI1575_LC_9_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNI1575_LC_9_3_2 (
            .in0(_gnd_net_),
            .in1(N__2905),
            .in2(N__3811),
            .in3(N__2938),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIZ0Z1575),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_9_3_3.C_ON=1'b1;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_9_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_9_3_3 (
            .in0(_gnd_net_),
            .in1(N__2919),
            .in2(_gnd_net_),
            .in3(N__2926),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_beamX_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_9_3_4.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_9_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_9_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2923),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_3_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_3_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_9_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2918),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_9_3_6.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_9_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_9_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_9_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2898),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23),
            .ltout(un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_9_3_7.C_ON=1'b0;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_9_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_9_3_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_9_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3244),
            .in3(_gnd_net_),
            .lcout(un1_beamX_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_4_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_4_0 (
            .in0(_gnd_net_),
            .in1(N__3927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQ1_LC_9_4_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQ1_LC_9_4_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQ1_LC_9_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQ1_LC_9_4_1 (
            .in0(_gnd_net_),
            .in1(N__3502),
            .in2(N__3192),
            .in3(N__3235),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNIN2AQZ0Z1),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTR2_LC_9_4_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTR2_LC_9_4_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTR2_LC_9_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTR2_LC_9_4_2 (
            .in0(_gnd_net_),
            .in1(N__3187),
            .in2(N__3232),
            .in3(N__3223),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNIGMTRZ0Z2),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPA3_LC_9_4_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPA3_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPA3_LC_9_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPA3_LC_9_4_3 (
            .in0(_gnd_net_),
            .in1(N__3220),
            .in2(N__3193),
            .in3(N__3214),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIUBPAZ0Z3),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMVQV7_LC_9_4_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMVQV7_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMVQV7_LC_9_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMVQV7_LC_9_4_4 (
            .in0(N__4125),
            .in1(N__3211),
            .in2(N__3166),
            .in3(N__3205),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_LC_9_4_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_LC_9_4_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_LC_9_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_LC_9_4_5 (
            .in0(_gnd_net_),
            .in1(N__3202),
            .in2(_gnd_net_),
            .in3(N__3196),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2FZ0Z4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_0_LC_9_4_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_0_LC_9_4_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_0_LC_9_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMFVC1_0_LC_9_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3183),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_4_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_4_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_4_7 (
            .in0(N__3928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_0.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3882),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_9_6_0.C_ON=1'b0;
    defparam beamY_0_LC_9_6_0.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_9_6_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_0_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(N__3494),
            .in2(_gnd_net_),
            .in3(N__3406),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3528),
            .ce(N__3464),
            .sr(_gnd_net_));
    defparam beamY_1_LC_9_6_5.C_ON=1'b0;
    defparam beamY_1_LC_9_6_5.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_9_6_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 beamY_1_LC_9_6_5 (
            .in0(N__3407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3366),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3528),
            .ce(N__3464),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_0_c_LC_9_7_0.C_ON=1'b1;
    defparam un5_visibley_cry_0_c_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_0_c_LC_9_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visibley_cry_0_c_LC_9_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3408),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(un5_visibley_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_9_7_1.C_ON=1'b1;
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_0_c_RNIJVSB_LC_9_7_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_0_c_RNIJVSB_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3367),
            .in3(N__3331),
            .lcout(un5_visibley_cry_0_c_RNIJVSBZ0),
            .ltout(),
            .carryin(un5_visibley_cry_0),
            .carryout(un5_visibley_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_9_7_2.C_ON=1'b1;
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_1_c_RNIL2UB_LC_9_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_1_c_RNIL2UB_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(N__3808),
            .in2(N__3328),
            .in3(N__3304),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visibley_cry_1),
            .carryout(un5_visibley_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_9_7_3.C_ON=1'b1;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_9_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_2_c_RNIN5VB_LC_9_7_3 (
            .in0(_gnd_net_),
            .in1(N__3805),
            .in2(N__3301),
            .in3(N__3277),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visibley_cry_2),
            .carryout(un5_visibley_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_3_c_RNIP80C_LC_9_7_4.C_ON=1'b1;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_9_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_3_c_RNIP80C_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__3809),
            .in2(N__3274),
            .in3(N__3247),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visibley_cry_3),
            .carryout(un5_visibley_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_9_7_5.C_ON=1'b1;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_9_7_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_4_c_RNIRB1C_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3955),
            .in3(N__3916),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visibley_cry_4),
            .carryout(un5_visibley_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_5_c_RNITE2C_LC_9_7_6.C_ON=1'b1;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_9_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_5_c_RNITE2C_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(N__3810),
            .in2(N__3912),
            .in3(N__3865),
            .lcout(un1_visibley_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visibley_cry_5),
            .carryout(un5_visibley_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_9_7_7.C_ON=1'b1;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_9_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_6_c_RNIVH3C_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(N__3806),
            .in2(N__3861),
            .in3(N__3817),
            .lcout(un1_visibley_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visibley_cry_6),
            .carryout(un5_visibley_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_9_8_0.C_ON=1'b1;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_9_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_7_c_RNI1L4C_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__3807),
            .in2(N__3687),
            .in3(N__3646),
            .lcout(un5_visibley_cry_7_c_RNI1L4CZ0),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(un5_visibley_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_9_8_1.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_9_8_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__3637),
            .in2(_gnd_net_),
            .in3(N__3616),
            .lcout(un1_visibley_if_generate_plus_mult1_un33_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_7_LC_11_2_3.C_ON=1'b0;
    defparam Pixel_1_RNO_7_LC_11_2_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_7_LC_11_2_3.LUT_INIT=16'b1110111111111111;
    LogicCell40 Pixel_1_RNO_7_LC_11_2_3 (
            .in0(N__4053),
            .in1(N__4038),
            .in2(N__4021),
            .in3(N__4060),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_3_LC_11_2_4.C_ON=1'b0;
    defparam Pixel_1_RNO_3_LC_11_2_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_3_LC_11_2_4.LUT_INIT=16'b0000000000110100;
    LogicCell40 Pixel_1_RNO_3_LC_11_2_4 (
            .in0(N__3988),
            .in1(N__4081),
            .in2(N__3598),
            .in3(N__4027),
            .lcout(),
            .ltout(un13_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_11_2_5.C_ON=1'b0;
    defparam Pixel_1_LC_11_2_5.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_11_2_5.LUT_INIT=16'b1100000010000100;
    LogicCell40 Pixel_1_LC_11_2_5 (
            .in0(N__3595),
            .in1(N__3586),
            .in2(N__3577),
            .in3(N__3574),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3532),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_3_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_3_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_3_0 (
            .in0(_gnd_net_),
            .in1(N__4013),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCH_LC_11_3_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCH_LC_11_3_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCH_LC_11_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCH_LC_11_3_1 (
            .in0(_gnd_net_),
            .in1(N__4096),
            .in2(N__4263),
            .in3(N__4087),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNI7TSCHZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6Q_LC_11_3_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6Q_LC_11_3_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6Q_LC_11_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6Q_LC_11_3_2 (
            .in0(_gnd_net_),
            .in1(N__4258),
            .in2(N__4366),
            .in3(N__4084),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNI8VC6QZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_9_LC_11_3_3.C_ON=1'b1;
    defparam Pixel_1_RNO_9_LC_11_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_9_LC_11_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_9_LC_11_3_3 (
            .in0(_gnd_net_),
            .in1(N__4348),
            .in2(N__4264),
            .in3(N__4075),
            .lcout(Pixel_1_RNOZ0Z_9),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_3_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_3_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_3_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_3_4 (
            .in0(_gnd_net_),
            .in1(N__4309),
            .in2(N__4072),
            .in3(N__4254),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDG11_LC_11_3_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDG11_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDG11_LC_11_3_5.LUT_INIT=16'b0000111111110000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDG11_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4285),
            .in3(N__4063),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11),
            .ltout(un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNICMDGZ0Z11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_8_LC_11_3_6.C_ON=1'b0;
    defparam Pixel_1_RNO_8_LC_11_3_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_8_LC_11_3_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_8_LC_11_3_6 (
            .in0(N__3961),
            .in1(N__4054),
            .in2(N__4042),
            .in3(N__4039),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_11_LC_11_3_7.C_ON=1'b0;
    defparam Pixel_1_RNO_11_LC_11_3_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_11_LC_11_3_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 Pixel_1_RNO_11_LC_11_3_7 (
            .in0(N__4014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3984),
            .lcout(G_7_i_a4_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_4_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_4_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_4_0 (
            .in0(_gnd_net_),
            .in1(N__4233),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGS4_LC_11_4_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGS4_LC_11_4_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGS4_LC_11_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGS4_LC_11_4_1 (
            .in0(_gnd_net_),
            .in1(N__4127),
            .in2(N__4201),
            .in3(N__4189),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNIUNGSZ0Z4),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEK6_LC_11_4_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEK6_LC_11_4_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEK6_LC_11_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEK6_LC_11_4_2 (
            .in0(_gnd_net_),
            .in1(N__4186),
            .in2(N__4132),
            .in3(N__4177),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNICUEKZ0Z6),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3M7_LC_11_4_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3M7_LC_11_4_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3M7_LC_11_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3M7_LC_11_4_3 (
            .in0(_gnd_net_),
            .in1(N__4131),
            .in2(N__4174),
            .in3(N__4162),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI6K3MZ0Z7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNI2S0GG_LC_11_4_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNI2S0GG_LC_11_4_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNI2S0GG_LC_11_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNI2S0GG_LC_11_4_4 (
            .in0(N__4333),
            .in1(N__4159),
            .in2(N__4105),
            .in3(N__4150),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_LC_11_4_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_LC_11_4_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_LC_11_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_LC_11_4_5 (
            .in0(_gnd_net_),
            .in1(N__4147),
            .in2(_gnd_net_),
            .in3(N__4138),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8),
            .ltout(un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0BZ0Z8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_0_LC_11_4_6.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_0_LC_11_4_6.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_0_LC_11_4_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDG0B8_0_LC_11_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4135),
            .in3(_gnd_net_),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_0_LC_11_4_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_0_LC_11_4_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_0_LC_11_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI1H2F4_0_LC_11_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4126),
            .lcout(un1_visibley_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_5_4.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_5_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4390),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(N__4389),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMR49_LC_12_4_1.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMR49_LC_12_4_1.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMR49_LC_12_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMR49_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__4334),
            .in2(N__4210),
            .in3(N__4357),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNIFMRZ0Z49),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LD_LC_12_4_2.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LD_LC_12_4_2.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LD_LC_12_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LD_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(N__4354),
            .in2(N__4339),
            .in3(N__4342),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI674LDZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DF_LC_12_4_3.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DF_LC_12_4_3.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DF_LC_12_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DF_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(N__4338),
            .in2(N__4318),
            .in3(N__4303),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNILF3DFZ0),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIG8GC11_LC_12_4_4.C_ON=1'b1;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIG8GC11_LC_12_4_4.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIG8GC11_LC_12_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIG8GC11_LC_12_4_4 (
            .in0(N__4262),
            .in1(N__4300),
            .in2(N__4294),
            .in3(N__4276),
            .lcout(un1_visibley_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_visibley_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTG_LC_12_4_5.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTG_LC_12_4_5.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTG_LC_12_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTG_LC_12_4_5 (
            .in0(_gnd_net_),
            .in1(N__4273),
            .in2(_gnd_net_),
            .in3(N__4267),
            .lcout(un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNI01NTGZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_7.C_ON=1'b0;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_7.SEQ_MODE=4'b0000;
    defparam un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4237),
            .lcout(un1_visibley_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
