// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 16:41:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSync,
    Pixel,
    HSync,
    Clock12MHz);

    output VSync;
    output Pixel;
    output HSync;
    input Clock12MHz;

    wire N__4026;
    wire N__4025;
    wire N__4024;
    wire N__4017;
    wire N__4016;
    wire N__4015;
    wire N__4008;
    wire N__4007;
    wire N__4006;
    wire N__3999;
    wire N__3998;
    wire N__3997;
    wire N__3980;
    wire N__3979;
    wire N__3978;
    wire N__3973;
    wire N__3972;
    wire N__3969;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3944;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3936;
    wire N__3935;
    wire N__3934;
    wire N__3933;
    wire N__3932;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3844;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3797;
    wire N__3794;
    wire N__3793;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3774;
    wire N__3771;
    wire N__3766;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3718;
    wire N__3717;
    wire N__3716;
    wire N__3715;
    wire N__3714;
    wire N__3713;
    wire N__3712;
    wire N__3711;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3685;
    wire N__3684;
    wire N__3681;
    wire N__3680;
    wire N__3677;
    wire N__3676;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3652;
    wire N__3649;
    wire N__3638;
    wire N__3635;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3538;
    wire N__3533;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3467;
    wire N__3464;
    wire N__3463;
    wire N__3462;
    wire N__3461;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3412;
    wire N__3411;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3389;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3361;
    wire N__3360;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3307;
    wire N__3306;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3298;
    wire N__3295;
    wire N__3294;
    wire N__3293;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3253;
    wire N__3250;
    wire N__3241;
    wire N__3236;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3217;
    wire N__3216;
    wire N__3211;
    wire N__3208;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3188;
    wire N__3185;
    wire N__3184;
    wire N__3183;
    wire N__3182;
    wire N__3179;
    wire N__3178;
    wire N__3175;
    wire N__3174;
    wire N__3171;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3153;
    wire N__3150;
    wire N__3143;
    wire N__3140;
    wire N__3131;
    wire N__3130;
    wire N__3129;
    wire N__3124;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3102;
    wire N__3095;
    wire N__3094;
    wire N__3093;
    wire N__3088;
    wire N__3087;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3048;
    wire N__3045;
    wire N__3044;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3029;
    wire N__3020;
    wire N__3017;
    wire N__3016;
    wire N__3015;
    wire N__3012;
    wire N__3007;
    wire N__3004;
    wire N__2999;
    wire N__2996;
    wire N__2995;
    wire N__2992;
    wire N__2991;
    wire N__2990;
    wire N__2987;
    wire N__2984;
    wire N__2977;
    wire N__2972;
    wire N__2969;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2959;
    wire N__2958;
    wire N__2957;
    wire N__2956;
    wire N__2955;
    wire N__2954;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2942;
    wire N__2933;
    wire N__2930;
    wire N__2929;
    wire N__2928;
    wire N__2927;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2899;
    wire N__2888;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2876;
    wire N__2873;
    wire N__2872;
    wire N__2871;
    wire N__2868;
    wire N__2863;
    wire N__2858;
    wire N__2857;
    wire N__2854;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2834;
    wire N__2833;
    wire N__2832;
    wire N__2831;
    wire N__2828;
    wire N__2821;
    wire N__2816;
    wire N__2815;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2779;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2741;
    wire N__2740;
    wire N__2737;
    wire N__2736;
    wire N__2735;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2702;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2691;
    wire N__2688;
    wire N__2687;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2672;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2641;
    wire N__2640;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2603;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2572;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2434;
    wire N__2431;
    wire N__2430;
    wire N__2429;
    wire N__2422;
    wire N__2419;
    wire N__2414;
    wire N__2413;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2290;
    wire N__2287;
    wire N__2286;
    wire N__2285;
    wire N__2278;
    wire N__2275;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2233;
    wire N__2232;
    wire N__2229;
    wire N__2228;
    wire N__2225;
    wire N__2224;
    wire N__2221;
    wire N__2212;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2179;
    wire N__2176;
    wire N__2173;
    wire N__2168;
    wire N__2167;
    wire N__2164;
    wire N__2161;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2111;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2096;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2066;
    wire N__2063;
    wire N__2060;
    wire N__2057;
    wire N__2054;
    wire N__2053;
    wire N__2050;
    wire N__2049;
    wire N__2048;
    wire N__2041;
    wire N__2038;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2015;
    wire N__2012;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2000;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1979;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1969;
    wire N__1966;
    wire N__1965;
    wire N__1964;
    wire N__1957;
    wire N__1954;
    wire N__1949;
    wire N__1946;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1922;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1907;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1877;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1865;
    wire N__1862;
    wire N__1859;
    wire N__1856;
    wire \VGAClock.PixelClock ;
    wire Clock12MHz_c;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_2_0_;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un61_sum_i_0;
    wire bfn_1_3_0_;
    wire un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5;
    wire un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_;
    wire un2_y_if_generate_plus_mult1_un61_sum_i_7;
    wire bfn_1_4_0_;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un61_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2;
    wire un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_;
    wire un2_y_if_generate_plus_mult1_un54_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_i_0;
    wire bfn_1_5_0_;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_;
    wire bfn_1_6_0_;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO;
    wire y_RNIA5P7Z0Z_9;
    wire bfn_2_2_0_;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0;
    wire un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un75_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_;
    wire un2_y_if_generate_plus_mult1_un68_sum_i_0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0;
    wire un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0;
    wire Pixel_RNOZ0Z_8;
    wire N_8_cascade_;
    wire N_11;
    wire un12_0_1_cascade_;
    wire Pixel_c;
    wire bfn_2_4_0_;
    wire un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un40_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un54_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91;
    wire un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_;
    wire un2_y_if_generate_plus_mult1_un47_sum_i_7;
    wire un2_y_if_generate_plus_mult1_un47_sum_i_0;
    wire bfn_2_5_0_;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_2;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_3;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_4;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2;
    wire un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5;
    wire un2_y_if_generate_plus_mult1_un47_sum_axb_7;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_5;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_6;
    wire un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire y_RNI94P7Z0Z_8;
    wire un2_y_if_generate_plus_mult1_un40_sum_i_0;
    wire G_7_i_a4_0_0;
    wire bfn_2_6_0_;
    wire un4_y_cry_1;
    wire un4_y_cry_2;
    wire un4_y_cry_3;
    wire un4_y_cry_4;
    wire un4_y_cry_5;
    wire un4_y_cry_6;
    wire un4_y_cry_7;
    wire un4_y_cry_8;
    wire bfn_2_7_0_;
    wire bfn_4_1_0_;
    wire un16_x_cry_1;
    wire un16_x_cry_2;
    wire un16_x_cry_3;
    wire un16_x_cry_4;
    wire un16_x_cry_5;
    wire un16_x_cry_6;
    wire un16_x_cry_7;
    wire un16_x_cry_8;
    wire bfn_4_2_0_;
    wire un8_xlt9_0;
    wire Pixel_0_sqmuxa_0_cascade_;
    wire Pixel_0_sqmuxa_1;
    wire bfn_4_3_0_;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un68_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_;
    wire Pixel_RNOZ0Z_5;
    wire un2_x_27;
    wire un2_x_if_generate_plus_mult1_un68_sum_i;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747;
    wire un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0;
    wire un13lt10;
    wire un1_ylto9_5_cascade_;
    wire un4_y_cry_2_THRU_CO;
    wire yZ0Z_5;
    wire yZ0Z_6;
    wire yZ0Z_1;
    wire un1_ylto9_4;
    wire un4_y_cry_1_THRU_CO;
    wire yZ0Z_4;
    wire yZ0Z_3;
    wire yZ0Z_2;
    wire yZ0Z_9;
    wire yZ0Z_8;
    wire y_12_5;
    wire y_12_6_cascade_;
    wire yZ0Z_7;
    wire y_12_8;
    wire y_12_8_cascade_;
    wire yZ0Z_0;
    wire un11_x_4_0_cascade_;
    wire x_RNID8R22Z0Z_9;
    wire xZ0Z_2;
    wire xZ0Z_1;
    wire xZ0Z_3;
    wire xZ0Z_0;
    wire bfn_5_2_0_;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_;
    wire un11_x_3_0;
    wire xZ0Z_4;
    wire un4_xlt9;
    wire xZ0Z_9;
    wire HSync_c;
    wire xZ0Z_8;
    wire un1_xlto9_0;
    wire bfn_5_3_0_;
    wire un2_x_if_generate_plus_mult1_un40_sum_i;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8;
    wire CONSTANT_ONE_NET;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0;
    wire bfn_5_4_0_;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un75_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5;
    wire un2_x_if_generate_plus_mult1_un61_sum_i;
    wire un1_y;
    wire VSync_c;
    wire PixelClock_g;
    wire xZ0Z_5;
    wire un11_x_4;
    wire bfn_6_3_0_;
    wire un2_x_if_generate_plus_mult1_un47_sum_i;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un47_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un54_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_;
    wire xZ0Z_7;
    wire xZ0Z_6;
    wire bfn_6_4_0_;
    wire un2_x_if_generate_plus_mult1_un54_sum_i;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_4;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_5;
    wire un2_x_if_generate_plus_mult1_un54_sum_i_8;
    wire un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0;
    wire un2_x_if_generate_plus_mult1_un68_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_6;
    wire un2_x_if_generate_plus_mult1_un61_sum_axb_8;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2;
    wire un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_;
    wire un2_x_if_generate_plus_mult1_un61_sum_i_8;
    wire _gnd_net_;

    defparam \VGAClock.PixelClock_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \VGAClock.PixelClock_inst .TEST_MODE=1'b0;
    defparam \VGAClock.PixelClock_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \VGAClock.PixelClock_inst .PLLOUT_SELECT="GENCLK";
    defparam \VGAClock.PixelClock_inst .FILTER_RANGE=3'b001;
    defparam \VGAClock.PixelClock_inst .FEEDBACK_PATH="SIMPLE";
    defparam \VGAClock.PixelClock_inst .FDA_RELATIVE=4'b0000;
    defparam \VGAClock.PixelClock_inst .FDA_FEEDBACK=4'b0000;
    defparam \VGAClock.PixelClock_inst .ENABLE_ICEGATE=1'b0;
    defparam \VGAClock.PixelClock_inst .DIVR=4'b0000;
    defparam \VGAClock.PixelClock_inst .DIVQ=3'b100;
    defparam \VGAClock.PixelClock_inst .DIVF=7'b1001010;
    defparam \VGAClock.PixelClock_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \VGAClock.PixelClock_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\VGAClock.PixelClock ),
            .REFERENCECLK(N__1865),
            .RESETB(N__3308),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__4026),
            .DIN(N__4025),
            .DOUT(N__4024),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__4026),
            .PADOUT(N__4025),
            .PADIN(N__4024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3731),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__4017),
            .DIN(N__4016),
            .DOUT(N__4015),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__4017),
            .PADOUT(N__4016),
            .PADIN(N__4015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3380),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__4008),
            .DIN(N__4007),
            .DOUT(N__4006),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__4008),
            .PADOUT(N__4007),
            .PADIN(N__4006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2132),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__3999),
            .DIN(N__3998),
            .DOUT(N__3997),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__3999),
            .PADOUT(N__3998),
            .PADIN(N__3997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__873 (
            .O(N__3980),
            .I(N__3973));
    InMux I__872 (
            .O(N__3979),
            .I(N__3973));
    InMux I__871 (
            .O(N__3978),
            .I(N__3969));
    LocalMux I__870 (
            .O(N__3973),
            .I(N__3965));
    InMux I__869 (
            .O(N__3972),
            .I(N__3962));
    LocalMux I__868 (
            .O(N__3969),
            .I(N__3959));
    InMux I__867 (
            .O(N__3968),
            .I(N__3956));
    Span4Mux_h I__866 (
            .O(N__3965),
            .I(N__3953));
    LocalMux I__865 (
            .O(N__3962),
            .I(xZ0Z_7));
    Odrv4 I__864 (
            .O(N__3959),
            .I(xZ0Z_7));
    LocalMux I__863 (
            .O(N__3956),
            .I(xZ0Z_7));
    Odrv4 I__862 (
            .O(N__3953),
            .I(xZ0Z_7));
    InMux I__861 (
            .O(N__3944),
            .I(N__3940));
    InMux I__860 (
            .O(N__3943),
            .I(N__3937));
    LocalMux I__859 (
            .O(N__3940),
            .I(N__3927));
    LocalMux I__858 (
            .O(N__3937),
            .I(N__3927));
    InMux I__857 (
            .O(N__3936),
            .I(N__3924));
    InMux I__856 (
            .O(N__3935),
            .I(N__3921));
    InMux I__855 (
            .O(N__3934),
            .I(N__3916));
    InMux I__854 (
            .O(N__3933),
            .I(N__3916));
    InMux I__853 (
            .O(N__3932),
            .I(N__3913));
    Span4Mux_h I__852 (
            .O(N__3927),
            .I(N__3910));
    LocalMux I__851 (
            .O(N__3924),
            .I(xZ0Z_6));
    LocalMux I__850 (
            .O(N__3921),
            .I(xZ0Z_6));
    LocalMux I__849 (
            .O(N__3916),
            .I(xZ0Z_6));
    LocalMux I__848 (
            .O(N__3913),
            .I(xZ0Z_6));
    Odrv4 I__847 (
            .O(N__3910),
            .I(xZ0Z_6));
    CascadeMux I__846 (
            .O(N__3899),
            .I(N__3896));
    InMux I__845 (
            .O(N__3896),
            .I(N__3893));
    LocalMux I__844 (
            .O(N__3893),
            .I(un2_x_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__843 (
            .O(N__3890),
            .I(N__3887));
    InMux I__842 (
            .O(N__3887),
            .I(N__3884));
    LocalMux I__841 (
            .O(N__3884),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02));
    InMux I__840 (
            .O(N__3881),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__839 (
            .O(N__3878),
            .I(N__3874));
    InMux I__838 (
            .O(N__3877),
            .I(N__3871));
    LocalMux I__837 (
            .O(N__3874),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1));
    LocalMux I__836 (
            .O(N__3871),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1));
    CascadeMux I__835 (
            .O(N__3866),
            .I(N__3863));
    InMux I__834 (
            .O(N__3863),
            .I(N__3860));
    LocalMux I__833 (
            .O(N__3860),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0));
    CascadeMux I__832 (
            .O(N__3857),
            .I(N__3854));
    InMux I__831 (
            .O(N__3854),
            .I(N__3851));
    LocalMux I__830 (
            .O(N__3851),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2));
    InMux I__829 (
            .O(N__3848),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__828 (
            .O(N__3845),
            .I(N__3839));
    InMux I__827 (
            .O(N__3844),
            .I(N__3839));
    LocalMux I__826 (
            .O(N__3839),
            .I(un2_x_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__825 (
            .O(N__3836),
            .I(N__3833));
    InMux I__824 (
            .O(N__3833),
            .I(N__3830));
    LocalMux I__823 (
            .O(N__3830),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0));
    InMux I__822 (
            .O(N__3827),
            .I(N__3824));
    LocalMux I__821 (
            .O(N__3824),
            .I(un2_x_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__820 (
            .O(N__3821),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__819 (
            .O(N__3818),
            .I(N__3815));
    LocalMux I__818 (
            .O(N__3815),
            .I(un2_x_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__817 (
            .O(N__3812),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__816 (
            .O(N__3809),
            .I(N__3805));
    InMux I__815 (
            .O(N__3808),
            .I(N__3802));
    LocalMux I__814 (
            .O(N__3805),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2));
    LocalMux I__813 (
            .O(N__3802),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2));
    CascadeMux I__812 (
            .O(N__3797),
            .I(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_));
    InMux I__811 (
            .O(N__3794),
            .I(N__3788));
    InMux I__810 (
            .O(N__3793),
            .I(N__3788));
    LocalMux I__809 (
            .O(N__3788),
            .I(un2_x_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__808 (
            .O(N__3785),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__807 (
            .O(N__3782),
            .I(N__3778));
    CascadeMux I__806 (
            .O(N__3781),
            .I(N__3775));
    LocalMux I__805 (
            .O(N__3778),
            .I(N__3771));
    InMux I__804 (
            .O(N__3775),
            .I(N__3766));
    InMux I__803 (
            .O(N__3774),
            .I(N__3766));
    Odrv4 I__802 (
            .O(N__3771),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5));
    LocalMux I__801 (
            .O(N__3766),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5));
    CascadeMux I__800 (
            .O(N__3761),
            .I(N__3758));
    InMux I__799 (
            .O(N__3758),
            .I(N__3755));
    LocalMux I__798 (
            .O(N__3755),
            .I(un2_x_if_generate_plus_mult1_un61_sum_i));
    InMux I__797 (
            .O(N__3752),
            .I(N__3749));
    LocalMux I__796 (
            .O(N__3749),
            .I(N__3745));
    InMux I__795 (
            .O(N__3748),
            .I(N__3742));
    Span4Mux_h I__794 (
            .O(N__3745),
            .I(N__3739));
    LocalMux I__793 (
            .O(N__3742),
            .I(N__3736));
    Odrv4 I__792 (
            .O(N__3739),
            .I(un1_y));
    Odrv4 I__791 (
            .O(N__3736),
            .I(un1_y));
    IoInMux I__790 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__789 (
            .O(N__3728),
            .I(N__3725));
    IoSpan4Mux I__788 (
            .O(N__3725),
            .I(N__3722));
    Odrv4 I__787 (
            .O(N__3722),
            .I(VSync_c));
    ClkMux I__786 (
            .O(N__3719),
            .I(N__3692));
    ClkMux I__785 (
            .O(N__3718),
            .I(N__3692));
    ClkMux I__784 (
            .O(N__3717),
            .I(N__3692));
    ClkMux I__783 (
            .O(N__3716),
            .I(N__3692));
    ClkMux I__782 (
            .O(N__3715),
            .I(N__3692));
    ClkMux I__781 (
            .O(N__3714),
            .I(N__3692));
    ClkMux I__780 (
            .O(N__3713),
            .I(N__3692));
    ClkMux I__779 (
            .O(N__3712),
            .I(N__3692));
    ClkMux I__778 (
            .O(N__3711),
            .I(N__3692));
    GlobalMux I__777 (
            .O(N__3692),
            .I(N__3689));
    gio2CtrlBuf I__776 (
            .O(N__3689),
            .I(PixelClock_g));
    InMux I__775 (
            .O(N__3686),
            .I(N__3681));
    CascadeMux I__774 (
            .O(N__3685),
            .I(N__3677));
    InMux I__773 (
            .O(N__3684),
            .I(N__3672));
    LocalMux I__772 (
            .O(N__3681),
            .I(N__3669));
    InMux I__771 (
            .O(N__3680),
            .I(N__3666));
    InMux I__770 (
            .O(N__3677),
            .I(N__3663));
    InMux I__769 (
            .O(N__3676),
            .I(N__3660));
    InMux I__768 (
            .O(N__3675),
            .I(N__3657));
    LocalMux I__767 (
            .O(N__3672),
            .I(N__3652));
    Span4Mux_h I__766 (
            .O(N__3669),
            .I(N__3652));
    LocalMux I__765 (
            .O(N__3666),
            .I(N__3649));
    LocalMux I__764 (
            .O(N__3663),
            .I(xZ0Z_5));
    LocalMux I__763 (
            .O(N__3660),
            .I(xZ0Z_5));
    LocalMux I__762 (
            .O(N__3657),
            .I(xZ0Z_5));
    Odrv4 I__761 (
            .O(N__3652),
            .I(xZ0Z_5));
    Odrv4 I__760 (
            .O(N__3649),
            .I(xZ0Z_5));
    InMux I__759 (
            .O(N__3638),
            .I(N__3635));
    LocalMux I__758 (
            .O(N__3635),
            .I(N__3631));
    InMux I__757 (
            .O(N__3634),
            .I(N__3628));
    Odrv4 I__756 (
            .O(N__3631),
            .I(un11_x_4));
    LocalMux I__755 (
            .O(N__3628),
            .I(un11_x_4));
    InMux I__754 (
            .O(N__3623),
            .I(N__3620));
    LocalMux I__753 (
            .O(N__3620),
            .I(un2_x_if_generate_plus_mult1_un47_sum_i));
    InMux I__752 (
            .O(N__3617),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__751 (
            .O(N__3614),
            .I(N__3610));
    InMux I__750 (
            .O(N__3613),
            .I(N__3607));
    LocalMux I__749 (
            .O(N__3610),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0));
    LocalMux I__748 (
            .O(N__3607),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0));
    CascadeMux I__747 (
            .O(N__3602),
            .I(N__3599));
    InMux I__746 (
            .O(N__3599),
            .I(N__3596));
    LocalMux I__745 (
            .O(N__3596),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0));
    InMux I__744 (
            .O(N__3593),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_5));
    CascadeMux I__743 (
            .O(N__3590),
            .I(N__3586));
    InMux I__742 (
            .O(N__3589),
            .I(N__3583));
    InMux I__741 (
            .O(N__3586),
            .I(N__3580));
    LocalMux I__740 (
            .O(N__3583),
            .I(un2_x_if_generate_plus_mult1_un47_sum_i_8));
    LocalMux I__739 (
            .O(N__3580),
            .I(un2_x_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__738 (
            .O(N__3575),
            .I(N__3572));
    InMux I__737 (
            .O(N__3572),
            .I(N__3569));
    LocalMux I__736 (
            .O(N__3569),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0));
    InMux I__735 (
            .O(N__3566),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__734 (
            .O(N__3563),
            .I(N__3560));
    LocalMux I__733 (
            .O(N__3560),
            .I(un2_x_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__732 (
            .O(N__3557),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__731 (
            .O(N__3554),
            .I(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_));
    InMux I__730 (
            .O(N__3551),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__729 (
            .O(N__3548),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7));
    CascadeMux I__728 (
            .O(N__3545),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_));
    CascadeMux I__727 (
            .O(N__3542),
            .I(N__3539));
    InMux I__726 (
            .O(N__3539),
            .I(N__3533));
    InMux I__725 (
            .O(N__3538),
            .I(N__3533));
    LocalMux I__724 (
            .O(N__3533),
            .I(N__3529));
    InMux I__723 (
            .O(N__3532),
            .I(N__3526));
    Odrv4 I__722 (
            .O(N__3529),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    LocalMux I__721 (
            .O(N__3526),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__720 (
            .O(N__3521),
            .I(N__3518));
    LocalMux I__719 (
            .O(N__3518),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0));
    InMux I__718 (
            .O(N__3515),
            .I(N__3512));
    LocalMux I__717 (
            .O(N__3512),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3));
    InMux I__716 (
            .O(N__3509),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__715 (
            .O(N__3506),
            .I(N__3503));
    InMux I__714 (
            .O(N__3503),
            .I(N__3500));
    LocalMux I__713 (
            .O(N__3500),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465));
    InMux I__712 (
            .O(N__3497),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__711 (
            .O(N__3494),
            .I(N__3491));
    LocalMux I__710 (
            .O(N__3491),
            .I(un2_x_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__709 (
            .O(N__3488),
            .I(un2_x_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__708 (
            .O(N__3485),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5));
    CascadeMux I__707 (
            .O(N__3482),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_));
    InMux I__706 (
            .O(N__3479),
            .I(N__3475));
    InMux I__705 (
            .O(N__3478),
            .I(N__3472));
    LocalMux I__704 (
            .O(N__3475),
            .I(un11_x_3_0));
    LocalMux I__703 (
            .O(N__3472),
            .I(un11_x_3_0));
    CascadeMux I__702 (
            .O(N__3467),
            .I(N__3464));
    InMux I__701 (
            .O(N__3464),
            .I(N__3451));
    InMux I__700 (
            .O(N__3463),
            .I(N__3451));
    InMux I__699 (
            .O(N__3462),
            .I(N__3451));
    CascadeMux I__698 (
            .O(N__3461),
            .I(N__3448));
    CascadeMux I__697 (
            .O(N__3460),
            .I(N__3445));
    InMux I__696 (
            .O(N__3459),
            .I(N__3442));
    InMux I__695 (
            .O(N__3458),
            .I(N__3439));
    LocalMux I__694 (
            .O(N__3451),
            .I(N__3436));
    InMux I__693 (
            .O(N__3448),
            .I(N__3433));
    InMux I__692 (
            .O(N__3445),
            .I(N__3430));
    LocalMux I__691 (
            .O(N__3442),
            .I(xZ0Z_4));
    LocalMux I__690 (
            .O(N__3439),
            .I(xZ0Z_4));
    Odrv4 I__689 (
            .O(N__3436),
            .I(xZ0Z_4));
    LocalMux I__688 (
            .O(N__3433),
            .I(xZ0Z_4));
    LocalMux I__687 (
            .O(N__3430),
            .I(xZ0Z_4));
    InMux I__686 (
            .O(N__3419),
            .I(N__3416));
    LocalMux I__685 (
            .O(N__3416),
            .I(un4_xlt9));
    CascadeMux I__684 (
            .O(N__3413),
            .I(N__3408));
    InMux I__683 (
            .O(N__3412),
            .I(N__3402));
    InMux I__682 (
            .O(N__3411),
            .I(N__3399));
    InMux I__681 (
            .O(N__3408),
            .I(N__3396));
    InMux I__680 (
            .O(N__3407),
            .I(N__3389));
    InMux I__679 (
            .O(N__3406),
            .I(N__3389));
    InMux I__678 (
            .O(N__3405),
            .I(N__3389));
    LocalMux I__677 (
            .O(N__3402),
            .I(xZ0Z_9));
    LocalMux I__676 (
            .O(N__3399),
            .I(xZ0Z_9));
    LocalMux I__675 (
            .O(N__3396),
            .I(xZ0Z_9));
    LocalMux I__674 (
            .O(N__3389),
            .I(xZ0Z_9));
    IoInMux I__673 (
            .O(N__3380),
            .I(N__3377));
    LocalMux I__672 (
            .O(N__3377),
            .I(N__3374));
    Span4Mux_s0_v I__671 (
            .O(N__3374),
            .I(N__3371));
    Span4Mux_h I__670 (
            .O(N__3371),
            .I(N__3368));
    Odrv4 I__669 (
            .O(N__3368),
            .I(HSync_c));
    CascadeMux I__668 (
            .O(N__3365),
            .I(N__3362));
    InMux I__667 (
            .O(N__3362),
            .I(N__3355));
    InMux I__666 (
            .O(N__3361),
            .I(N__3352));
    InMux I__665 (
            .O(N__3360),
            .I(N__3349));
    InMux I__664 (
            .O(N__3359),
            .I(N__3346));
    InMux I__663 (
            .O(N__3358),
            .I(N__3343));
    LocalMux I__662 (
            .O(N__3355),
            .I(N__3340));
    LocalMux I__661 (
            .O(N__3352),
            .I(xZ0Z_8));
    LocalMux I__660 (
            .O(N__3349),
            .I(xZ0Z_8));
    LocalMux I__659 (
            .O(N__3346),
            .I(xZ0Z_8));
    LocalMux I__658 (
            .O(N__3343),
            .I(xZ0Z_8));
    Odrv4 I__657 (
            .O(N__3340),
            .I(xZ0Z_8));
    InMux I__656 (
            .O(N__3329),
            .I(N__3326));
    LocalMux I__655 (
            .O(N__3326),
            .I(un1_xlto9_0));
    InMux I__654 (
            .O(N__3323),
            .I(N__3320));
    LocalMux I__653 (
            .O(N__3320),
            .I(un2_x_if_generate_plus_mult1_un40_sum_i));
    InMux I__652 (
            .O(N__3317),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__651 (
            .O(N__3314),
            .I(N__3311));
    LocalMux I__650 (
            .O(N__3311),
            .I(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8));
    IoInMux I__649 (
            .O(N__3308),
            .I(N__3302));
    CascadeMux I__648 (
            .O(N__3307),
            .I(N__3299));
    CascadeMux I__647 (
            .O(N__3306),
            .I(N__3295));
    CascadeMux I__646 (
            .O(N__3305),
            .I(N__3289));
    LocalMux I__645 (
            .O(N__3302),
            .I(N__3286));
    InMux I__644 (
            .O(N__3299),
            .I(N__3279));
    InMux I__643 (
            .O(N__3298),
            .I(N__3279));
    InMux I__642 (
            .O(N__3295),
            .I(N__3279));
    CascadeMux I__641 (
            .O(N__3294),
            .I(N__3276));
    CascadeMux I__640 (
            .O(N__3293),
            .I(N__3273));
    CascadeMux I__639 (
            .O(N__3292),
            .I(N__3270));
    InMux I__638 (
            .O(N__3289),
            .I(N__3267));
    Span4Mux_s0_v I__637 (
            .O(N__3286),
            .I(N__3264));
    LocalMux I__636 (
            .O(N__3279),
            .I(N__3261));
    InMux I__635 (
            .O(N__3276),
            .I(N__3258));
    InMux I__634 (
            .O(N__3273),
            .I(N__3253));
    InMux I__633 (
            .O(N__3270),
            .I(N__3253));
    LocalMux I__632 (
            .O(N__3267),
            .I(N__3250));
    Span4Mux_v I__631 (
            .O(N__3264),
            .I(N__3241));
    Span4Mux_s1_h I__630 (
            .O(N__3261),
            .I(N__3241));
    LocalMux I__629 (
            .O(N__3258),
            .I(N__3241));
    LocalMux I__628 (
            .O(N__3253),
            .I(N__3241));
    Odrv4 I__627 (
            .O(N__3250),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__626 (
            .O(N__3241),
            .I(CONSTANT_ONE_NET));
    InMux I__625 (
            .O(N__3236),
            .I(un2_x_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__624 (
            .O(N__3233),
            .I(N__3227));
    InMux I__623 (
            .O(N__3232),
            .I(N__3224));
    InMux I__622 (
            .O(N__3231),
            .I(N__3221));
    CascadeMux I__621 (
            .O(N__3230),
            .I(N__3218));
    LocalMux I__620 (
            .O(N__3227),
            .I(N__3211));
    LocalMux I__619 (
            .O(N__3224),
            .I(N__3211));
    LocalMux I__618 (
            .O(N__3221),
            .I(N__3208));
    InMux I__617 (
            .O(N__3218),
            .I(N__3203));
    InMux I__616 (
            .O(N__3217),
            .I(N__3203));
    InMux I__615 (
            .O(N__3216),
            .I(N__3200));
    Span4Mux_h I__614 (
            .O(N__3211),
            .I(N__3197));
    Odrv12 I__613 (
            .O(N__3208),
            .I(yZ0Z_3));
    LocalMux I__612 (
            .O(N__3203),
            .I(yZ0Z_3));
    LocalMux I__611 (
            .O(N__3200),
            .I(yZ0Z_3));
    Odrv4 I__610 (
            .O(N__3197),
            .I(yZ0Z_3));
    CascadeMux I__609 (
            .O(N__3188),
            .I(N__3185));
    InMux I__608 (
            .O(N__3185),
            .I(N__3179));
    InMux I__607 (
            .O(N__3184),
            .I(N__3175));
    CascadeMux I__606 (
            .O(N__3183),
            .I(N__3171));
    InMux I__605 (
            .O(N__3182),
            .I(N__3167));
    LocalMux I__604 (
            .O(N__3179),
            .I(N__3164));
    InMux I__603 (
            .O(N__3178),
            .I(N__3161));
    LocalMux I__602 (
            .O(N__3175),
            .I(N__3158));
    InMux I__601 (
            .O(N__3174),
            .I(N__3153));
    InMux I__600 (
            .O(N__3171),
            .I(N__3153));
    InMux I__599 (
            .O(N__3170),
            .I(N__3150));
    LocalMux I__598 (
            .O(N__3167),
            .I(N__3143));
    Span4Mux_v I__597 (
            .O(N__3164),
            .I(N__3143));
    LocalMux I__596 (
            .O(N__3161),
            .I(N__3143));
    Span4Mux_s3_h I__595 (
            .O(N__3158),
            .I(N__3140));
    LocalMux I__594 (
            .O(N__3153),
            .I(yZ0Z_2));
    LocalMux I__593 (
            .O(N__3150),
            .I(yZ0Z_2));
    Odrv4 I__592 (
            .O(N__3143),
            .I(yZ0Z_2));
    Odrv4 I__591 (
            .O(N__3140),
            .I(yZ0Z_2));
    InMux I__590 (
            .O(N__3131),
            .I(N__3124));
    InMux I__589 (
            .O(N__3130),
            .I(N__3124));
    CascadeMux I__588 (
            .O(N__3129),
            .I(N__3120));
    LocalMux I__587 (
            .O(N__3124),
            .I(N__3117));
    CascadeMux I__586 (
            .O(N__3123),
            .I(N__3113));
    InMux I__585 (
            .O(N__3120),
            .I(N__3110));
    Span4Mux_v I__584 (
            .O(N__3117),
            .I(N__3107));
    InMux I__583 (
            .O(N__3116),
            .I(N__3102));
    InMux I__582 (
            .O(N__3113),
            .I(N__3102));
    LocalMux I__581 (
            .O(N__3110),
            .I(yZ0Z_9));
    Odrv4 I__580 (
            .O(N__3107),
            .I(yZ0Z_9));
    LocalMux I__579 (
            .O(N__3102),
            .I(yZ0Z_9));
    InMux I__578 (
            .O(N__3095),
            .I(N__3088));
    InMux I__577 (
            .O(N__3094),
            .I(N__3088));
    InMux I__576 (
            .O(N__3093),
            .I(N__3083));
    LocalMux I__575 (
            .O(N__3088),
            .I(N__3080));
    InMux I__574 (
            .O(N__3087),
            .I(N__3077));
    InMux I__573 (
            .O(N__3086),
            .I(N__3074));
    LocalMux I__572 (
            .O(N__3083),
            .I(yZ0Z_8));
    Odrv4 I__571 (
            .O(N__3080),
            .I(yZ0Z_8));
    LocalMux I__570 (
            .O(N__3077),
            .I(yZ0Z_8));
    LocalMux I__569 (
            .O(N__3074),
            .I(yZ0Z_8));
    InMux I__568 (
            .O(N__3065),
            .I(N__3062));
    LocalMux I__567 (
            .O(N__3062),
            .I(y_12_5));
    CascadeMux I__566 (
            .O(N__3059),
            .I(y_12_6_cascade_));
    InMux I__565 (
            .O(N__3056),
            .I(N__3052));
    InMux I__564 (
            .O(N__3055),
            .I(N__3049));
    LocalMux I__563 (
            .O(N__3052),
            .I(N__3045));
    LocalMux I__562 (
            .O(N__3049),
            .I(N__3040));
    InMux I__561 (
            .O(N__3048),
            .I(N__3037));
    Span4Mux_h I__560 (
            .O(N__3045),
            .I(N__3034));
    InMux I__559 (
            .O(N__3044),
            .I(N__3029));
    InMux I__558 (
            .O(N__3043),
            .I(N__3029));
    Odrv4 I__557 (
            .O(N__3040),
            .I(yZ0Z_7));
    LocalMux I__556 (
            .O(N__3037),
            .I(yZ0Z_7));
    Odrv4 I__555 (
            .O(N__3034),
            .I(yZ0Z_7));
    LocalMux I__554 (
            .O(N__3029),
            .I(yZ0Z_7));
    InMux I__553 (
            .O(N__3020),
            .I(N__3017));
    LocalMux I__552 (
            .O(N__3017),
            .I(N__3012));
    InMux I__551 (
            .O(N__3016),
            .I(N__3007));
    InMux I__550 (
            .O(N__3015),
            .I(N__3007));
    Span4Mux_s3_h I__549 (
            .O(N__3012),
            .I(N__3004));
    LocalMux I__548 (
            .O(N__3007),
            .I(y_12_8));
    Odrv4 I__547 (
            .O(N__3004),
            .I(y_12_8));
    CascadeMux I__546 (
            .O(N__2999),
            .I(y_12_8_cascade_));
    InMux I__545 (
            .O(N__2996),
            .I(N__2992));
    CascadeMux I__544 (
            .O(N__2995),
            .I(N__2987));
    LocalMux I__543 (
            .O(N__2992),
            .I(N__2984));
    InMux I__542 (
            .O(N__2991),
            .I(N__2977));
    InMux I__541 (
            .O(N__2990),
            .I(N__2977));
    InMux I__540 (
            .O(N__2987),
            .I(N__2977));
    Odrv12 I__539 (
            .O(N__2984),
            .I(yZ0Z_0));
    LocalMux I__538 (
            .O(N__2977),
            .I(yZ0Z_0));
    CascadeMux I__537 (
            .O(N__2972),
            .I(un11_x_4_0_cascade_));
    InMux I__536 (
            .O(N__2969),
            .I(N__2959));
    InMux I__535 (
            .O(N__2968),
            .I(N__2959));
    InMux I__534 (
            .O(N__2967),
            .I(N__2959));
    InMux I__533 (
            .O(N__2966),
            .I(N__2950));
    LocalMux I__532 (
            .O(N__2959),
            .I(N__2947));
    InMux I__531 (
            .O(N__2958),
            .I(N__2942));
    InMux I__530 (
            .O(N__2957),
            .I(N__2942));
    InMux I__529 (
            .O(N__2956),
            .I(N__2933));
    InMux I__528 (
            .O(N__2955),
            .I(N__2933));
    InMux I__527 (
            .O(N__2954),
            .I(N__2933));
    InMux I__526 (
            .O(N__2953),
            .I(N__2933));
    LocalMux I__525 (
            .O(N__2950),
            .I(N__2930));
    Sp12to4 I__524 (
            .O(N__2947),
            .I(N__2922));
    LocalMux I__523 (
            .O(N__2942),
            .I(N__2922));
    LocalMux I__522 (
            .O(N__2933),
            .I(N__2919));
    Span4Mux_h I__521 (
            .O(N__2930),
            .I(N__2916));
    InMux I__520 (
            .O(N__2929),
            .I(N__2913));
    InMux I__519 (
            .O(N__2928),
            .I(N__2910));
    InMux I__518 (
            .O(N__2927),
            .I(N__2907));
    Span12Mux_s4_h I__517 (
            .O(N__2922),
            .I(N__2904));
    Span4Mux_v I__516 (
            .O(N__2919),
            .I(N__2899));
    Span4Mux_v I__515 (
            .O(N__2916),
            .I(N__2899));
    LocalMux I__514 (
            .O(N__2913),
            .I(x_RNID8R22Z0Z_9));
    LocalMux I__513 (
            .O(N__2910),
            .I(x_RNID8R22Z0Z_9));
    LocalMux I__512 (
            .O(N__2907),
            .I(x_RNID8R22Z0Z_9));
    Odrv12 I__511 (
            .O(N__2904),
            .I(x_RNID8R22Z0Z_9));
    Odrv4 I__510 (
            .O(N__2899),
            .I(x_RNID8R22Z0Z_9));
    InMux I__509 (
            .O(N__2888),
            .I(N__2884));
    InMux I__508 (
            .O(N__2887),
            .I(N__2881));
    LocalMux I__507 (
            .O(N__2884),
            .I(xZ0Z_2));
    LocalMux I__506 (
            .O(N__2881),
            .I(xZ0Z_2));
    CascadeMux I__505 (
            .O(N__2876),
            .I(N__2873));
    InMux I__504 (
            .O(N__2873),
            .I(N__2868));
    InMux I__503 (
            .O(N__2872),
            .I(N__2863));
    InMux I__502 (
            .O(N__2871),
            .I(N__2863));
    LocalMux I__501 (
            .O(N__2868),
            .I(xZ0Z_1));
    LocalMux I__500 (
            .O(N__2863),
            .I(xZ0Z_1));
    InMux I__499 (
            .O(N__2858),
            .I(N__2854));
    CascadeMux I__498 (
            .O(N__2857),
            .I(N__2850));
    LocalMux I__497 (
            .O(N__2854),
            .I(N__2847));
    InMux I__496 (
            .O(N__2853),
            .I(N__2844));
    InMux I__495 (
            .O(N__2850),
            .I(N__2841));
    Odrv4 I__494 (
            .O(N__2847),
            .I(xZ0Z_3));
    LocalMux I__493 (
            .O(N__2844),
            .I(xZ0Z_3));
    LocalMux I__492 (
            .O(N__2841),
            .I(xZ0Z_3));
    InMux I__491 (
            .O(N__2834),
            .I(N__2828));
    InMux I__490 (
            .O(N__2833),
            .I(N__2821));
    InMux I__489 (
            .O(N__2832),
            .I(N__2821));
    InMux I__488 (
            .O(N__2831),
            .I(N__2821));
    LocalMux I__487 (
            .O(N__2828),
            .I(xZ0Z_0));
    LocalMux I__486 (
            .O(N__2821),
            .I(xZ0Z_0));
    InMux I__485 (
            .O(N__2816),
            .I(N__2810));
    InMux I__484 (
            .O(N__2815),
            .I(N__2810));
    LocalMux I__483 (
            .O(N__2810),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747));
    InMux I__482 (
            .O(N__2807),
            .I(N__2804));
    LocalMux I__481 (
            .O(N__2804),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0));
    InMux I__480 (
            .O(N__2801),
            .I(N__2798));
    LocalMux I__479 (
            .O(N__2798),
            .I(N__2795));
    Odrv12 I__478 (
            .O(N__2795),
            .I(un13lt10));
    CascadeMux I__477 (
            .O(N__2792),
            .I(un1_ylto9_5_cascade_));
    InMux I__476 (
            .O(N__2789),
            .I(N__2786));
    LocalMux I__475 (
            .O(N__2786),
            .I(N__2783));
    Odrv12 I__474 (
            .O(N__2783),
            .I(un4_y_cry_2_THRU_CO));
    InMux I__473 (
            .O(N__2780),
            .I(N__2776));
    InMux I__472 (
            .O(N__2779),
            .I(N__2770));
    LocalMux I__471 (
            .O(N__2776),
            .I(N__2767));
    InMux I__470 (
            .O(N__2775),
            .I(N__2762));
    InMux I__469 (
            .O(N__2774),
            .I(N__2762));
    InMux I__468 (
            .O(N__2773),
            .I(N__2759));
    LocalMux I__467 (
            .O(N__2770),
            .I(N__2756));
    Span4Mux_h I__466 (
            .O(N__2767),
            .I(N__2753));
    LocalMux I__465 (
            .O(N__2762),
            .I(N__2750));
    LocalMux I__464 (
            .O(N__2759),
            .I(yZ0Z_5));
    Odrv4 I__463 (
            .O(N__2756),
            .I(yZ0Z_5));
    Odrv4 I__462 (
            .O(N__2753),
            .I(yZ0Z_5));
    Odrv4 I__461 (
            .O(N__2750),
            .I(yZ0Z_5));
    InMux I__460 (
            .O(N__2741),
            .I(N__2737));
    InMux I__459 (
            .O(N__2740),
            .I(N__2731));
    LocalMux I__458 (
            .O(N__2737),
            .I(N__2728));
    InMux I__457 (
            .O(N__2736),
            .I(N__2723));
    InMux I__456 (
            .O(N__2735),
            .I(N__2723));
    InMux I__455 (
            .O(N__2734),
            .I(N__2720));
    LocalMux I__454 (
            .O(N__2731),
            .I(N__2717));
    Span4Mux_h I__453 (
            .O(N__2728),
            .I(N__2714));
    LocalMux I__452 (
            .O(N__2723),
            .I(N__2711));
    LocalMux I__451 (
            .O(N__2720),
            .I(yZ0Z_6));
    Odrv4 I__450 (
            .O(N__2717),
            .I(yZ0Z_6));
    Odrv4 I__449 (
            .O(N__2714),
            .I(yZ0Z_6));
    Odrv4 I__448 (
            .O(N__2711),
            .I(yZ0Z_6));
    InMux I__447 (
            .O(N__2702),
            .I(N__2698));
    CascadeMux I__446 (
            .O(N__2701),
            .I(N__2695));
    LocalMux I__445 (
            .O(N__2698),
            .I(N__2692));
    InMux I__444 (
            .O(N__2695),
            .I(N__2688));
    Span4Mux_s3_h I__443 (
            .O(N__2692),
            .I(N__2683));
    InMux I__442 (
            .O(N__2691),
            .I(N__2680));
    LocalMux I__441 (
            .O(N__2688),
            .I(N__2677));
    InMux I__440 (
            .O(N__2687),
            .I(N__2672));
    InMux I__439 (
            .O(N__2686),
            .I(N__2672));
    Odrv4 I__438 (
            .O(N__2683),
            .I(yZ0Z_1));
    LocalMux I__437 (
            .O(N__2680),
            .I(yZ0Z_1));
    Odrv12 I__436 (
            .O(N__2677),
            .I(yZ0Z_1));
    LocalMux I__435 (
            .O(N__2672),
            .I(yZ0Z_1));
    InMux I__434 (
            .O(N__2663),
            .I(N__2660));
    LocalMux I__433 (
            .O(N__2660),
            .I(un1_ylto9_4));
    CascadeMux I__432 (
            .O(N__2657),
            .I(N__2654));
    InMux I__431 (
            .O(N__2654),
            .I(N__2651));
    LocalMux I__430 (
            .O(N__2651),
            .I(N__2648));
    Odrv4 I__429 (
            .O(N__2648),
            .I(un4_y_cry_1_THRU_CO));
    CascadeMux I__428 (
            .O(N__2645),
            .I(N__2642));
    InMux I__427 (
            .O(N__2642),
            .I(N__2636));
    InMux I__426 (
            .O(N__2641),
            .I(N__2633));
    CascadeMux I__425 (
            .O(N__2640),
            .I(N__2630));
    InMux I__424 (
            .O(N__2639),
            .I(N__2626));
    LocalMux I__423 (
            .O(N__2636),
            .I(N__2623));
    LocalMux I__422 (
            .O(N__2633),
            .I(N__2620));
    InMux I__421 (
            .O(N__2630),
            .I(N__2617));
    InMux I__420 (
            .O(N__2629),
            .I(N__2614));
    LocalMux I__419 (
            .O(N__2626),
            .I(N__2611));
    Span4Mux_h I__418 (
            .O(N__2623),
            .I(N__2608));
    Span4Mux_s1_h I__417 (
            .O(N__2620),
            .I(N__2603));
    LocalMux I__416 (
            .O(N__2617),
            .I(N__2603));
    LocalMux I__415 (
            .O(N__2614),
            .I(yZ0Z_4));
    Odrv4 I__414 (
            .O(N__2611),
            .I(yZ0Z_4));
    Odrv4 I__413 (
            .O(N__2608),
            .I(yZ0Z_4));
    Odrv4 I__412 (
            .O(N__2603),
            .I(yZ0Z_4));
    CascadeMux I__411 (
            .O(N__2594),
            .I(Pixel_0_sqmuxa_0_cascade_));
    InMux I__410 (
            .O(N__2591),
            .I(N__2588));
    LocalMux I__409 (
            .O(N__2588),
            .I(N__2585));
    Span4Mux_s3_h I__408 (
            .O(N__2585),
            .I(N__2582));
    Odrv4 I__407 (
            .O(N__2582),
            .I(Pixel_0_sqmuxa_1));
    InMux I__406 (
            .O(N__2579),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__405 (
            .O(N__2576),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__404 (
            .O(N__2573),
            .I(N__2567));
    InMux I__403 (
            .O(N__2572),
            .I(N__2567));
    LocalMux I__402 (
            .O(N__2567),
            .I(un2_x_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__401 (
            .O(N__2564),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__400 (
            .O(N__2561),
            .I(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_));
    InMux I__399 (
            .O(N__2558),
            .I(N__2555));
    LocalMux I__398 (
            .O(N__2555),
            .I(Pixel_RNOZ0Z_5));
    InMux I__397 (
            .O(N__2552),
            .I(N__2549));
    LocalMux I__396 (
            .O(N__2549),
            .I(N__2546));
    Odrv12 I__395 (
            .O(N__2546),
            .I(un2_x_27));
    CascadeMux I__394 (
            .O(N__2543),
            .I(N__2540));
    InMux I__393 (
            .O(N__2540),
            .I(N__2537));
    LocalMux I__392 (
            .O(N__2537),
            .I(un2_x_if_generate_plus_mult1_un68_sum_i));
    InMux I__391 (
            .O(N__2534),
            .I(un16_x_cry_1));
    InMux I__390 (
            .O(N__2531),
            .I(un16_x_cry_2));
    InMux I__389 (
            .O(N__2528),
            .I(un16_x_cry_3));
    InMux I__388 (
            .O(N__2525),
            .I(un16_x_cry_4));
    InMux I__387 (
            .O(N__2522),
            .I(un16_x_cry_5));
    InMux I__386 (
            .O(N__2519),
            .I(un16_x_cry_6));
    InMux I__385 (
            .O(N__2516),
            .I(un16_x_cry_7));
    InMux I__384 (
            .O(N__2513),
            .I(bfn_4_2_0_));
    CascadeMux I__383 (
            .O(N__2510),
            .I(N__2507));
    InMux I__382 (
            .O(N__2507),
            .I(N__2504));
    LocalMux I__381 (
            .O(N__2504),
            .I(un8_xlt9_0));
    InMux I__380 (
            .O(N__2501),
            .I(un4_y_cry_1));
    InMux I__379 (
            .O(N__2498),
            .I(un4_y_cry_2));
    InMux I__378 (
            .O(N__2495),
            .I(un4_y_cry_3));
    InMux I__377 (
            .O(N__2492),
            .I(un4_y_cry_4));
    InMux I__376 (
            .O(N__2489),
            .I(un4_y_cry_5));
    InMux I__375 (
            .O(N__2486),
            .I(un4_y_cry_6));
    InMux I__374 (
            .O(N__2483),
            .I(un4_y_cry_7));
    InMux I__373 (
            .O(N__2480),
            .I(bfn_2_7_0_));
    InMux I__372 (
            .O(N__2477),
            .I(N__2474));
    LocalMux I__371 (
            .O(N__2474),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0));
    InMux I__370 (
            .O(N__2471),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__369 (
            .O(N__2468),
            .I(N__2465));
    LocalMux I__368 (
            .O(N__2465),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0));
    CascadeMux I__367 (
            .O(N__2462),
            .I(N__2459));
    InMux I__366 (
            .O(N__2459),
            .I(N__2456));
    LocalMux I__365 (
            .O(N__2456),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0));
    InMux I__364 (
            .O(N__2453),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__363 (
            .O(N__2450),
            .I(N__2447));
    LocalMux I__362 (
            .O(N__2447),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0));
    InMux I__361 (
            .O(N__2444),
            .I(N__2441));
    LocalMux I__360 (
            .O(N__2441),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0));
    InMux I__359 (
            .O(N__2438),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__358 (
            .O(N__2435),
            .I(N__2431));
    InMux I__357 (
            .O(N__2434),
            .I(N__2422));
    InMux I__356 (
            .O(N__2431),
            .I(N__2422));
    InMux I__355 (
            .O(N__2430),
            .I(N__2422));
    InMux I__354 (
            .O(N__2429),
            .I(N__2419));
    LocalMux I__353 (
            .O(N__2422),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0));
    LocalMux I__352 (
            .O(N__2419),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0));
    InMux I__351 (
            .O(N__2414),
            .I(N__2409));
    InMux I__350 (
            .O(N__2413),
            .I(N__2406));
    InMux I__349 (
            .O(N__2412),
            .I(N__2403));
    LocalMux I__348 (
            .O(N__2409),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2));
    LocalMux I__347 (
            .O(N__2406),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2));
    LocalMux I__346 (
            .O(N__2403),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2));
    CascadeMux I__345 (
            .O(N__2396),
            .I(N__2393));
    InMux I__344 (
            .O(N__2393),
            .I(N__2390));
    LocalMux I__343 (
            .O(N__2390),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5));
    InMux I__342 (
            .O(N__2387),
            .I(N__2384));
    LocalMux I__341 (
            .O(N__2384),
            .I(un2_y_if_generate_plus_mult1_un47_sum_axb_7));
    InMux I__340 (
            .O(N__2381),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__339 (
            .O(N__2378),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__338 (
            .O(N__2375),
            .I(N__2372));
    InMux I__337 (
            .O(N__2372),
            .I(N__2369));
    LocalMux I__336 (
            .O(N__2369),
            .I(un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__335 (
            .O(N__2366),
            .I(N__2363));
    LocalMux I__334 (
            .O(N__2363),
            .I(y_RNI94P7Z0Z_8));
    CascadeMux I__333 (
            .O(N__2360),
            .I(N__2357));
    InMux I__332 (
            .O(N__2357),
            .I(N__2354));
    LocalMux I__331 (
            .O(N__2354),
            .I(un2_y_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__330 (
            .O(N__2351),
            .I(N__2348));
    LocalMux I__329 (
            .O(N__2348),
            .I(N__2345));
    Odrv12 I__328 (
            .O(N__2345),
            .I(G_7_i_a4_0_0));
    InMux I__327 (
            .O(N__2342),
            .I(N__2339));
    LocalMux I__326 (
            .O(N__2339),
            .I(un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21));
    InMux I__325 (
            .O(N__2336),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__324 (
            .O(N__2333),
            .I(N__2330));
    InMux I__323 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__322 (
            .O(N__2327),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81));
    InMux I__321 (
            .O(N__2324),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__320 (
            .O(N__2321),
            .I(N__2318));
    LocalMux I__319 (
            .O(N__2318),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1));
    InMux I__318 (
            .O(N__2315),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__317 (
            .O(N__2312),
            .I(N__2309));
    InMux I__316 (
            .O(N__2309),
            .I(N__2306));
    LocalMux I__315 (
            .O(N__2306),
            .I(un2_y_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__314 (
            .O(N__2303),
            .I(N__2300));
    LocalMux I__313 (
            .O(N__2300),
            .I(un2_y_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__312 (
            .O(N__2297),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__311 (
            .O(N__2294),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__310 (
            .O(N__2291),
            .I(N__2287));
    InMux I__309 (
            .O(N__2290),
            .I(N__2278));
    InMux I__308 (
            .O(N__2287),
            .I(N__2278));
    InMux I__307 (
            .O(N__2286),
            .I(N__2278));
    InMux I__306 (
            .O(N__2285),
            .I(N__2275));
    LocalMux I__305 (
            .O(N__2278),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91));
    LocalMux I__304 (
            .O(N__2275),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91));
    CascadeMux I__303 (
            .O(N__2270),
            .I(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_));
    CascadeMux I__302 (
            .O(N__2267),
            .I(N__2264));
    InMux I__301 (
            .O(N__2264),
            .I(N__2261));
    LocalMux I__300 (
            .O(N__2261),
            .I(un2_y_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__299 (
            .O(N__2258),
            .I(N__2255));
    InMux I__298 (
            .O(N__2255),
            .I(N__2252));
    LocalMux I__297 (
            .O(N__2252),
            .I(un2_y_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__296 (
            .O(N__2249),
            .I(N__2246));
    LocalMux I__295 (
            .O(N__2246),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9));
    InMux I__294 (
            .O(N__2243),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__293 (
            .O(N__2240),
            .I(N__2237));
    LocalMux I__292 (
            .O(N__2237),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0));
    CascadeMux I__291 (
            .O(N__2234),
            .I(N__2229));
    CascadeMux I__290 (
            .O(N__2233),
            .I(N__2225));
    InMux I__289 (
            .O(N__2232),
            .I(N__2221));
    InMux I__288 (
            .O(N__2229),
            .I(N__2212));
    InMux I__287 (
            .O(N__2228),
            .I(N__2212));
    InMux I__286 (
            .O(N__2225),
            .I(N__2212));
    InMux I__285 (
            .O(N__2224),
            .I(N__2212));
    LocalMux I__284 (
            .O(N__2221),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0));
    LocalMux I__283 (
            .O(N__2212),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0));
    CascadeMux I__282 (
            .O(N__2207),
            .I(N__2204));
    InMux I__281 (
            .O(N__2204),
            .I(N__2201));
    LocalMux I__280 (
            .O(N__2201),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0));
    InMux I__279 (
            .O(N__2198),
            .I(N__2195));
    LocalMux I__278 (
            .O(N__2195),
            .I(un2_y_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__277 (
            .O(N__2192),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6));
    CascadeMux I__276 (
            .O(N__2189),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_));
    InMux I__275 (
            .O(N__2186),
            .I(N__2183));
    LocalMux I__274 (
            .O(N__2183),
            .I(un2_y_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__273 (
            .O(N__2180),
            .I(N__2176));
    InMux I__272 (
            .O(N__2179),
            .I(N__2173));
    LocalMux I__271 (
            .O(N__2176),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0));
    LocalMux I__270 (
            .O(N__2173),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0));
    InMux I__269 (
            .O(N__2168),
            .I(N__2164));
    InMux I__268 (
            .O(N__2167),
            .I(N__2161));
    LocalMux I__267 (
            .O(N__2164),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0));
    LocalMux I__266 (
            .O(N__2161),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0));
    InMux I__265 (
            .O(N__2156),
            .I(N__2153));
    LocalMux I__264 (
            .O(N__2153),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0));
    InMux I__263 (
            .O(N__2150),
            .I(N__2147));
    LocalMux I__262 (
            .O(N__2147),
            .I(Pixel_RNOZ0Z_8));
    CascadeMux I__261 (
            .O(N__2144),
            .I(N_8_cascade_));
    InMux I__260 (
            .O(N__2141),
            .I(N__2138));
    LocalMux I__259 (
            .O(N__2138),
            .I(N_11));
    CascadeMux I__258 (
            .O(N__2135),
            .I(un12_0_1_cascade_));
    IoInMux I__257 (
            .O(N__2132),
            .I(N__2129));
    LocalMux I__256 (
            .O(N__2129),
            .I(N__2126));
    IoSpan4Mux I__255 (
            .O(N__2126),
            .I(N__2123));
    Span4Mux_s1_v I__254 (
            .O(N__2123),
            .I(N__2120));
    Span4Mux_h I__253 (
            .O(N__2120),
            .I(N__2117));
    Odrv4 I__252 (
            .O(N__2117),
            .I(Pixel_c));
    InMux I__251 (
            .O(N__2114),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_5));
    CascadeMux I__250 (
            .O(N__2111),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_));
    InMux I__249 (
            .O(N__2108),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_2));
    CascadeMux I__248 (
            .O(N__2105),
            .I(N__2102));
    InMux I__247 (
            .O(N__2102),
            .I(N__2099));
    LocalMux I__246 (
            .O(N__2099),
            .I(un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO));
    InMux I__245 (
            .O(N__2096),
            .I(N__2093));
    LocalMux I__244 (
            .O(N__2093),
            .I(y_RNIA5P7Z0Z_9));
    InMux I__243 (
            .O(N__2090),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__242 (
            .O(N__2087),
            .I(N__2084));
    InMux I__241 (
            .O(N__2084),
            .I(N__2081));
    LocalMux I__240 (
            .O(N__2081),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6));
    InMux I__239 (
            .O(N__2078),
            .I(un2_y_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__238 (
            .O(N__2075),
            .I(N__2072));
    LocalMux I__237 (
            .O(N__2072),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2));
    InMux I__236 (
            .O(N__2069),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__235 (
            .O(N__2066),
            .I(N__2063));
    LocalMux I__234 (
            .O(N__2063),
            .I(un2_y_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__233 (
            .O(N__2060),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__232 (
            .O(N__2057),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__231 (
            .O(N__2054),
            .I(N__2050));
    InMux I__230 (
            .O(N__2053),
            .I(N__2041));
    InMux I__229 (
            .O(N__2050),
            .I(N__2041));
    InMux I__228 (
            .O(N__2049),
            .I(N__2041));
    InMux I__227 (
            .O(N__2048),
            .I(N__2038));
    LocalMux I__226 (
            .O(N__2041),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2));
    LocalMux I__225 (
            .O(N__2038),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2));
    CascadeMux I__224 (
            .O(N__2033),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_));
    CascadeMux I__223 (
            .O(N__2030),
            .I(N__2027));
    InMux I__222 (
            .O(N__2027),
            .I(N__2024));
    LocalMux I__221 (
            .O(N__2024),
            .I(un2_y_if_generate_plus_mult1_un54_sum_i_7));
    CascadeMux I__220 (
            .O(N__2021),
            .I(N__2018));
    InMux I__219 (
            .O(N__2018),
            .I(N__2015));
    LocalMux I__218 (
            .O(N__2015),
            .I(un2_y_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__217 (
            .O(N__2012),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__216 (
            .O(N__2009),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__215 (
            .O(N__2006),
            .I(un2_y_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__214 (
            .O(N__2003),
            .I(N__2000));
    InMux I__213 (
            .O(N__2000),
            .I(N__1997));
    LocalMux I__212 (
            .O(N__1997),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4));
    InMux I__211 (
            .O(N__1994),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__210 (
            .O(N__1991),
            .I(N__1988));
    LocalMux I__209 (
            .O(N__1988),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5));
    InMux I__208 (
            .O(N__1985),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__207 (
            .O(N__1982),
            .I(N__1979));
    LocalMux I__206 (
            .O(N__1979),
            .I(un2_y_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__205 (
            .O(N__1976),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__204 (
            .O(N__1973),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__203 (
            .O(N__1970),
            .I(N__1966));
    InMux I__202 (
            .O(N__1969),
            .I(N__1957));
    InMux I__201 (
            .O(N__1966),
            .I(N__1957));
    InMux I__200 (
            .O(N__1965),
            .I(N__1957));
    InMux I__199 (
            .O(N__1964),
            .I(N__1954));
    LocalMux I__198 (
            .O(N__1957),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5));
    LocalMux I__197 (
            .O(N__1954),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5));
    CascadeMux I__196 (
            .O(N__1949),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_));
    CascadeMux I__195 (
            .O(N__1946),
            .I(N__1943));
    InMux I__194 (
            .O(N__1943),
            .I(N__1940));
    LocalMux I__193 (
            .O(N__1940),
            .I(un2_y_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__192 (
            .O(N__1937),
            .I(N__1934));
    LocalMux I__191 (
            .O(N__1934),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1));
    InMux I__190 (
            .O(N__1931),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__189 (
            .O(N__1928),
            .I(N__1925));
    InMux I__188 (
            .O(N__1925),
            .I(N__1922));
    LocalMux I__187 (
            .O(N__1922),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2));
    InMux I__186 (
            .O(N__1919),
            .I(un2_y_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__185 (
            .O(N__1916),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__184 (
            .O(N__1913),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__183 (
            .O(N__1910),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__182 (
            .O(N__1907),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__181 (
            .O(N__1904),
            .I(un2_y_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__180 (
            .O(N__1901),
            .I(N__1898));
    InMux I__179 (
            .O(N__1898),
            .I(N__1895));
    LocalMux I__178 (
            .O(N__1895),
            .I(un2_y_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__177 (
            .O(N__1892),
            .I(N__1889));
    LocalMux I__176 (
            .O(N__1889),
            .I(un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083));
    InMux I__175 (
            .O(N__1886),
            .I(un2_y_if_generate_plus_mult1_un61_sum_cry_2));
    IoInMux I__174 (
            .O(N__1883),
            .I(N__1880));
    LocalMux I__173 (
            .O(N__1880),
            .I(N__1877));
    Span4Mux_s1_h I__172 (
            .O(N__1877),
            .I(N__1874));
    Span4Mux_h I__171 (
            .O(N__1874),
            .I(N__1871));
    Sp12to4 I__170 (
            .O(N__1871),
            .I(N__1868));
    Odrv12 I__169 (
            .O(N__1868),
            .I(\VGAClock.PixelClock ));
    IoInMux I__168 (
            .O(N__1865),
            .I(N__1862));
    LocalMux I__167 (
            .O(N__1862),
            .I(N__1859));
    IoSpan4Mux I__166 (
            .O(N__1859),
            .I(N__1856));
    Odrv4 I__165 (
            .O(N__1856),
            .I(Clock12MHz_c));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_4_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_1_0_));
    defparam IN_MUX_bfv_4_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_2_0_ (
            .carryinitin(un16_x_cry_8),
            .carryinitout(bfn_4_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(un4_y_cry_8),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    ICE_GB \VGAClock.PLLOUTCORE_derived_clock_RNIE579  (
            .USERSIGNALTOGLOBALBUFFER(N__1883),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_2_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_2_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_2_0 (
            .in0(_gnd_net_),
            .in1(N__3232),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJ6_LC_1_2_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJ6_LC_1_2_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJ6_LC_1_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJ6_LC_1_2_1 (
            .in0(_gnd_net_),
            .in1(N__1965),
            .in2(N__1901),
            .in3(N__1916),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_2_c_RNILCRJZ0Z6),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8E9_LC_1_2_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8E9_LC_1_2_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8E9_LC_1_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8E9_LC_1_2_2 (
            .in0(_gnd_net_),
            .in1(N__1892),
            .in2(N__1970),
            .in3(N__1913),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_3_c_RNIGA8EZ0Z9),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10B_LC_1_2_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10B_LC_1_2_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10B_LC_1_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10B_LC_1_2_3 (
            .in0(_gnd_net_),
            .in1(N__1969),
            .in2(N__2003),
            .in3(N__1910),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_4_c_RNIKA10BZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAIONN_LC_1_2_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAIONN_LC_1_2_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAIONN_LC_1_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAIONN_LC_1_2_4 (
            .in0(N__2232),
            .in1(N__1991),
            .in2(N__1946),
            .in3(N__1907),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUB_LC_1_2_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUB_LC_1_2_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUB_LC_1_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUB_LC_1_2_5 (
            .in0(_gnd_net_),
            .in1(N__1982),
            .in2(_gnd_net_),
            .in3(N__1904),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_cry_6_c_RNI1NVUBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_2_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_2_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2641),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_3_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_3_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2640),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILP083_LC_1_3_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILP083_LC_1_3_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILP083_LC_1_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILP083_LC_1_3_1 (
            .in0(_gnd_net_),
            .in1(N__2049),
            .in2(N__2021),
            .in3(N__1886),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_sbtinv_RNILPZ0Z083),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOP4_LC_1_3_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOP4_LC_1_3_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOP4_LC_1_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOP4_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(N__1937),
            .in2(N__2054),
            .in3(N__1994),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_3_c_RNIONOPZ0Z4),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FI5_LC_1_3_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FI5_LC_1_3_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FI5_LC_1_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FI5_LC_1_3_3 (
            .in0(_gnd_net_),
            .in1(N__2053),
            .in2(N__1928),
            .in3(N__1985),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_4_c_RNIC6FIZ0Z5),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGA9KB_LC_1_3_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGA9KB_LC_1_3_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGA9KB_LC_1_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGA9KB_LC_1_3_4 (
            .in0(N__1964),
            .in1(N__2075),
            .in2(N__2030),
            .in3(N__1976),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_LC_1_3_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_LC_1_3_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_LC_1_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_LC_1_3_5 (
            .in0(_gnd_net_),
            .in1(N__2066),
            .in2(_gnd_net_),
            .in3(N__1973),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5),
            .ltout(un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKRZ0Z5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_0_LC_1_3_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_0_LC_1_3_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_0_LC_1_3_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un61_sum_cry_6_c_RNIDAKR5_0_LC_1_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1949),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(N__2774),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFL1_LC_1_4_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFL1_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFL1_LC_1_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFL1_LC_1_4_1 (
            .in0(_gnd_net_),
            .in1(N__2286),
            .in2(N__2258),
            .in3(N__1931),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_2_c_RNIVEFLZ0Z1),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4E2_LC_1_4_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4E2_LC_1_4_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4E2_LC_1_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4E2_LC_1_4_2 (
            .in0(_gnd_net_),
            .in1(N__2342),
            .in2(N__2291),
            .in3(N__1919),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIR4EZ0Z2),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9K2_LC_1_4_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9K2_LC_1_4_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9K2_LC_1_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9K2_LC_1_4_3 (
            .in0(_gnd_net_),
            .in1(N__2290),
            .in2(N__2333),
            .in3(N__2069),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_4_c_RNI8J9KZ0Z2),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNI3IEJ5_LC_1_4_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNI3IEJ5_LC_1_4_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNI3IEJ5_LC_1_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_5_c_RNI3IEJ5_LC_1_4_4 (
            .in0(N__2048),
            .in1(N__2321),
            .in2(N__2267),
            .in3(N__2060),
            .lcout(un2_y_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_LC_1_4_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_LC_1_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(N__2303),
            .in2(_gnd_net_),
            .in3(N__2057),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2),
            .ltout(un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6SZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_0_LC_1_4_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_0_LC_1_4_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_0_LC_1_4_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_cry_6_c_RNIIM6S2_0_LC_1_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2033),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_4_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_4_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_4_7 (
            .in0(N__2775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_5_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_LC_1_5_0 (
            .in0(_gnd_net_),
            .in1(N__3086),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_5_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KA_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__2096),
            .in2(N__3306),
            .in3(N__2012),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_2_c_RNIF6KAZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_5_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFF_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(N__3298),
            .in2(N__2105),
            .in3(N__2009),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_3_c_RNIDRFFZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75T2_LC_1_5_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75T2_LC_1_5_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75T2_LC_1_5_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75T2_LC_1_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3307),
            .in3(N__2006),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNI75TZ0Z2),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un33_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_LC_1_5_4.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_LC_1_5_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_LC_1_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2375),
            .in3(N__2114),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0),
            .ltout(un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4CZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_0_LC_1_5_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_0_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_0_LC_1_5_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_5_c_RNIFP4C_0_LC_1_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2111),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQ5_LC_1_5_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQ5_LC_1_5_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQ5_LC_1_5_6.LUT_INIT=16'b0110011001100110;
    LogicCell40 un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQ5_LC_1_5_6 (
            .in0(N__2412),
            .in1(N__2413),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEAQZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_1_6_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_1_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_2_c_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3123),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(un2_y_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_1_6_1.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_1_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2108),
            .lcout(un2_y_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIA5P7_9_LC_1_6_3.C_ON=1'b0;
    defparam y_RNIA5P7_9_LC_1_6_3.SEQ_MODE=4'b0000;
    defparam y_RNIA5P7_9_LC_1_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 y_RNIA5P7_9_LC_1_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3116),
            .lcout(y_RNIA5P7Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_2_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_2_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_2_0 (
            .in0(_gnd_net_),
            .in1(N__3184),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCC_LC_2_2_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCC_LC_2_2_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCC_LC_2_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCC_LC_2_2_1 (
            .in0(_gnd_net_),
            .in1(N__2186),
            .in2(N__2233),
            .in3(N__2090),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_2_c_RNIEFHCCZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJI_LC_2_2_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJI_LC_2_2_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJI_LC_2_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJI_LC_2_2_2 (
            .in0(_gnd_net_),
            .in1(N__2228),
            .in2(N__2087),
            .in3(N__2078),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2JLJIZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_8_LC_2_2_3.C_ON=1'b1;
    defparam Pixel_RNO_8_LC_2_2_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_8_LC_2_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_8_LC_2_2_3 (
            .in0(_gnd_net_),
            .in1(N__2249),
            .in2(N__2234),
            .in3(N__2243),
            .lcout(Pixel_RNOZ0Z_8),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_2_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_2_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_2_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_2_4 (
            .in0(_gnd_net_),
            .in1(N__2240),
            .in2(N__2207),
            .in3(N__2224),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MON_LC_2_2_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MON_LC_2_2_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MON_LC_2_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MON_LC_2_2_5 (
            .in0(_gnd_net_),
            .in1(N__2198),
            .in2(_gnd_net_),
            .in3(N__2192),
            .lcout(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0),
            .ltout(un2_y_if_generate_plus_mult1_un75_sum_cry_6_c_RNIP7MONZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_7_LC_2_2_6.C_ON=1'b0;
    defparam Pixel_RNO_7_LC_2_2_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_7_LC_2_2_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_RNO_7_LC_2_2_6 (
            .in0(N__2351),
            .in1(N__2180),
            .in2(N__2189),
            .in3(N__2167),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_2_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_2_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_2_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_2_7 (
            .in0(N__3233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_6_LC_2_3_3.C_ON=1'b0;
    defparam Pixel_RNO_6_LC_2_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_6_LC_2_3_3.LUT_INIT=16'b1110111111111111;
    LogicCell40 Pixel_RNO_6_LC_2_3_3 (
            .in0(N__2179),
            .in1(N__2168),
            .in2(N__3188),
            .in3(N__2156),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_2_LC_2_3_4.C_ON=1'b0;
    defparam Pixel_RNO_2_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_2_LC_2_3_4.LUT_INIT=16'b0000000000110100;
    LogicCell40 Pixel_RNO_2_LC_2_3_4 (
            .in0(N__2702),
            .in1(N__2150),
            .in2(N__2144),
            .in3(N__2141),
            .lcout(),
            .ltout(un12_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_2_3_5.C_ON=1'b0;
    defparam PixelZ0_LC_2_3_5.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_2_3_5.LUT_INIT=16'b1100000010000100;
    LogicCell40 PixelZ0_LC_2_3_5 (
            .in0(N__2801),
            .in1(N__2591),
            .in2(N__2135),
            .in3(N__2552),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3714),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0 (
            .in0(_gnd_net_),
            .in1(N__2735),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIG21_LC_2_4_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIG21_LC_2_4_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIG21_LC_2_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIG21_LC_2_4_1 (
            .in0(_gnd_net_),
            .in1(N__2430),
            .in2(N__2360),
            .in3(N__2336),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_sbtinv_RNIHIGZ0Z21),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68K81_LC_2_4_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68K81_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68K81_LC_2_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68K81_LC_2_4_2 (
            .in0(_gnd_net_),
            .in1(N__2477),
            .in2(N__2435),
            .in3(N__2324),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_3_c_RNI68KZ0Z81),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHB1_LC_2_4_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHB1_LC_2_4_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHB1_LC_2_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHB1_LC_2_4_3 (
            .in0(_gnd_net_),
            .in1(N__2434),
            .in2(N__2462),
            .in3(N__2315),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEEHBZ0Z1),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI678Q2_LC_2_4_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI678Q2_LC_2_4_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI678Q2_LC_2_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_5_c_RNI678Q2_LC_2_4_4 (
            .in0(N__2285),
            .in1(N__2444),
            .in2(N__2312),
            .in3(N__2297),
            .lcout(un2_y_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_LC_2_4_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_LC_2_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_LC_2_4_5 (
            .in0(_gnd_net_),
            .in1(N__2387),
            .in2(_gnd_net_),
            .in3(N__2294),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91),
            .ltout(un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVOZ0Z91_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_0_LC_2_4_6.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_0_LC_2_4_6.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_0_LC_2_4_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_cry_6_c_RNIOVO91_0_LC_2_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2270),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_4_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_4_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un47_sum_sbtinv_LC_2_4_7 (
            .in0(N__2736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_5_0.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_5_0 (
            .in0(_gnd_net_),
            .in1(N__3043),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERG_LC_2_5_1.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERG_LC_2_5_1.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERG_LC_2_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERG_LC_2_5_1 (
            .in0(_gnd_net_),
            .in1(N__2366),
            .in2(N__3292),
            .in3(N__2471),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_2_c_RNICERGZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJ_LC_2_5_2.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJ_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJ_LC_2_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJ_LC_2_5_2 (
            .in0(_gnd_net_),
            .in1(N__2468),
            .in2(N__3294),
            .in3(N__2453),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_3_c_RNIJINJZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KO_LC_2_5_3.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KO_LC_2_5_3.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KO_LC_2_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KO_LC_2_5_3 (
            .in0(_gnd_net_),
            .in1(N__2450),
            .in2(N__3293),
            .in3(N__2438),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_4_c_RNII9KOZ0),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNIAP1U_LC_2_5_4.C_ON=1'b1;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNIAP1U_LC_2_5_4.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNIAP1U_LC_2_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_5_c_RNIAP1U_LC_2_5_4 (
            .in0(N__2429),
            .in1(N__2414),
            .in2(N__2396),
            .in3(N__2381),
            .lcout(un2_y_if_generate_plus_mult1_un47_sum_axb_7),
            .ltout(),
            .carryin(un2_y_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un2_y_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_5_5.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_5_5.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_2_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2378),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNI94P7_8_LC_2_5_6.C_ON=1'b0;
    defparam y_RNI94P7_8_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam y_RNI94P7_8_LC_2_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 y_RNI94P7_8_LC_2_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3087),
            .lcout(y_RNI94P7Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_7.C_ON=1'b0;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un2_y_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_7 (
            .in0(N__3044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_y_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_11_LC_2_6_0.C_ON=1'b1;
    defparam Pixel_RNO_11_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_11_LC_2_6_0.LUT_INIT=16'b0000000011110000;
    LogicCell40 Pixel_RNO_11_LC_2_6_0 (
            .in0(_gnd_net_),
            .in1(N__2996),
            .in2(N__2701),
            .in3(N__3178),
            .lcout(G_7_i_a4_0_0),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(un4_y_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_y_cry_1_THRU_LUT4_0_LC_2_6_1.C_ON=1'b1;
    defparam un4_y_cry_1_THRU_LUT4_0_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam un4_y_cry_1_THRU_LUT4_0_LC_2_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_y_cry_1_THRU_LUT4_0_LC_2_6_1 (
            .in0(_gnd_net_),
            .in1(N__3182),
            .in2(_gnd_net_),
            .in3(N__2501),
            .lcout(un4_y_cry_1_THRU_CO),
            .ltout(),
            .carryin(un4_y_cry_1),
            .carryout(un4_y_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_y_cry_2_THRU_LUT4_0_LC_2_6_2.C_ON=1'b1;
    defparam un4_y_cry_2_THRU_LUT4_0_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam un4_y_cry_2_THRU_LUT4_0_LC_2_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_y_cry_2_THRU_LUT4_0_LC_2_6_2 (
            .in0(_gnd_net_),
            .in1(N__3231),
            .in2(_gnd_net_),
            .in3(N__2498),
            .lcout(un4_y_cry_2_THRU_CO),
            .ltout(),
            .carryin(un4_y_cry_2),
            .carryout(un4_y_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_4_LC_2_6_3.C_ON=1'b1;
    defparam y_4_LC_2_6_3.SEQ_MODE=4'b1000;
    defparam y_4_LC_2_6_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_4_LC_2_6_3 (
            .in0(N__2967),
            .in1(N__2629),
            .in2(_gnd_net_),
            .in3(N__2495),
            .lcout(yZ0Z_4),
            .ltout(),
            .carryin(un4_y_cry_3),
            .carryout(un4_y_cry_4),
            .clk(N__3712),
            .ce(),
            .sr(_gnd_net_));
    defparam y_5_LC_2_6_4.C_ON=1'b1;
    defparam y_5_LC_2_6_4.SEQ_MODE=4'b1000;
    defparam y_5_LC_2_6_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_5_LC_2_6_4 (
            .in0(N__2957),
            .in1(N__2773),
            .in2(_gnd_net_),
            .in3(N__2492),
            .lcout(yZ0Z_5),
            .ltout(),
            .carryin(un4_y_cry_4),
            .carryout(un4_y_cry_5),
            .clk(N__3712),
            .ce(),
            .sr(_gnd_net_));
    defparam y_6_LC_2_6_5.C_ON=1'b1;
    defparam y_6_LC_2_6_5.SEQ_MODE=4'b1000;
    defparam y_6_LC_2_6_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_6_LC_2_6_5 (
            .in0(N__2968),
            .in1(N__2734),
            .in2(_gnd_net_),
            .in3(N__2489),
            .lcout(yZ0Z_6),
            .ltout(),
            .carryin(un4_y_cry_5),
            .carryout(un4_y_cry_6),
            .clk(N__3712),
            .ce(),
            .sr(_gnd_net_));
    defparam y_7_LC_2_6_6.C_ON=1'b1;
    defparam y_7_LC_2_6_6.SEQ_MODE=4'b1000;
    defparam y_7_LC_2_6_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_7_LC_2_6_6 (
            .in0(N__2958),
            .in1(N__3048),
            .in2(_gnd_net_),
            .in3(N__2486),
            .lcout(yZ0Z_7),
            .ltout(),
            .carryin(un4_y_cry_6),
            .carryout(un4_y_cry_7),
            .clk(N__3712),
            .ce(),
            .sr(_gnd_net_));
    defparam y_8_LC_2_6_7.C_ON=1'b1;
    defparam y_8_LC_2_6_7.SEQ_MODE=4'b1000;
    defparam y_8_LC_2_6_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_8_LC_2_6_7 (
            .in0(N__2969),
            .in1(N__3093),
            .in2(_gnd_net_),
            .in3(N__2483),
            .lcout(yZ0Z_8),
            .ltout(),
            .carryin(un4_y_cry_7),
            .carryout(un4_y_cry_8),
            .clk(N__3712),
            .ce(),
            .sr(_gnd_net_));
    defparam y_9_LC_2_7_0.C_ON=1'b0;
    defparam y_9_LC_2_7_0.SEQ_MODE=4'b1000;
    defparam y_9_LC_2_7_0.LUT_INIT=16'b0011010001110000;
    LogicCell40 y_9_LC_2_7_0 (
            .in0(N__3020),
            .in1(N__2966),
            .in2(N__3129),
            .in3(N__2480),
            .lcout(yZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3711),
            .ce(),
            .sr(_gnd_net_));
    defparam un16_x_cry_1_c_LC_4_1_0.C_ON=1'b1;
    defparam un16_x_cry_1_c_LC_4_1_0.SEQ_MODE=4'b0000;
    defparam un16_x_cry_1_c_LC_4_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un16_x_cry_1_c_LC_4_1_0 (
            .in0(_gnd_net_),
            .in1(N__2834),
            .in2(N__2876),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_1_0_),
            .carryout(un16_x_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_2_LC_4_1_1.C_ON=1'b1;
    defparam x_2_LC_4_1_1.SEQ_MODE=4'b1000;
    defparam x_2_LC_4_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_2_LC_4_1_1 (
            .in0(_gnd_net_),
            .in1(N__2888),
            .in2(_gnd_net_),
            .in3(N__2534),
            .lcout(xZ0Z_2),
            .ltout(),
            .carryin(un16_x_cry_1),
            .carryout(un16_x_cry_2),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_3_LC_4_1_2.C_ON=1'b1;
    defparam x_3_LC_4_1_2.SEQ_MODE=4'b1000;
    defparam x_3_LC_4_1_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_3_LC_4_1_2 (
            .in0(_gnd_net_),
            .in1(N__2853),
            .in2(_gnd_net_),
            .in3(N__2531),
            .lcout(xZ0Z_3),
            .ltout(),
            .carryin(un16_x_cry_2),
            .carryout(un16_x_cry_3),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_4_LC_4_1_3.C_ON=1'b1;
    defparam x_4_LC_4_1_3.SEQ_MODE=4'b1000;
    defparam x_4_LC_4_1_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_4_LC_4_1_3 (
            .in0(_gnd_net_),
            .in1(N__3459),
            .in2(_gnd_net_),
            .in3(N__2528),
            .lcout(xZ0Z_4),
            .ltout(),
            .carryin(un16_x_cry_3),
            .carryout(un16_x_cry_4),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_5_LC_4_1_4.C_ON=1'b1;
    defparam x_5_LC_4_1_4.SEQ_MODE=4'b1000;
    defparam x_5_LC_4_1_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 x_5_LC_4_1_4 (
            .in0(N__2928),
            .in1(N__3676),
            .in2(_gnd_net_),
            .in3(N__2525),
            .lcout(xZ0Z_5),
            .ltout(),
            .carryin(un16_x_cry_4),
            .carryout(un16_x_cry_5),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_6_LC_4_1_5.C_ON=1'b1;
    defparam x_6_LC_4_1_5.SEQ_MODE=4'b1000;
    defparam x_6_LC_4_1_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_6_LC_4_1_5 (
            .in0(_gnd_net_),
            .in1(N__3936),
            .in2(_gnd_net_),
            .in3(N__2522),
            .lcout(xZ0Z_6),
            .ltout(),
            .carryin(un16_x_cry_5),
            .carryout(un16_x_cry_6),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_7_LC_4_1_6.C_ON=1'b1;
    defparam x_7_LC_4_1_6.SEQ_MODE=4'b1000;
    defparam x_7_LC_4_1_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 x_7_LC_4_1_6 (
            .in0(_gnd_net_),
            .in1(N__3972),
            .in2(_gnd_net_),
            .in3(N__2519),
            .lcout(xZ0Z_7),
            .ltout(),
            .carryin(un16_x_cry_6),
            .carryout(un16_x_cry_7),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_8_LC_4_1_7.C_ON=1'b1;
    defparam x_8_LC_4_1_7.SEQ_MODE=4'b1000;
    defparam x_8_LC_4_1_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 x_8_LC_4_1_7 (
            .in0(N__2927),
            .in1(N__3361),
            .in2(_gnd_net_),
            .in3(N__2516),
            .lcout(xZ0Z_8),
            .ltout(),
            .carryin(un16_x_cry_7),
            .carryout(un16_x_cry_8),
            .clk(N__3716),
            .ce(),
            .sr(_gnd_net_));
    defparam x_9_LC_4_2_0.C_ON=1'b0;
    defparam x_9_LC_4_2_0.SEQ_MODE=4'b1000;
    defparam x_9_LC_4_2_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 x_9_LC_4_2_0 (
            .in0(N__3412),
            .in1(N__2929),
            .in2(_gnd_net_),
            .in3(N__2513),
            .lcout(xZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3715),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_10_LC_4_2_5.C_ON=1'b0;
    defparam Pixel_RNO_10_LC_4_2_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_10_LC_4_2_5.LUT_INIT=16'b1111111000000000;
    LogicCell40 Pixel_RNO_10_LC_4_2_5 (
            .in0(N__3675),
            .in1(N__3932),
            .in2(N__3460),
            .in3(N__3968),
            .lcout(un8_xlt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_4_LC_4_2_6.C_ON=1'b0;
    defparam Pixel_RNO_4_LC_4_2_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_4_LC_4_2_6.LUT_INIT=16'b1011101111111100;
    LogicCell40 Pixel_RNO_4_LC_4_2_6 (
            .in0(N__3419),
            .in1(N__3359),
            .in2(N__2510),
            .in3(N__3411),
            .lcout(),
            .ltout(Pixel_0_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_0_LC_4_2_7.C_ON=1'b0;
    defparam Pixel_RNO_0_LC_4_2_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_0_LC_4_2_7.LUT_INIT=16'b0101000001010000;
    LogicCell40 Pixel_RNO_0_LC_4_2_7 (
            .in0(N__3748),
            .in1(_gnd_net_),
            .in2(N__2594),
            .in3(_gnd_net_),
            .lcout(Pixel_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_4_3_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_4_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(N__3462),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_4_3_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_4_3_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_4_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIH747_LC_4_3_1 (
            .in0(_gnd_net_),
            .in1(N__2572),
            .in2(N__2543),
            .in3(N__2579),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_cry_4_c_RNIHZ0Z747),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_5_LC_4_3_2.C_ON=1'b1;
    defparam Pixel_RNO_5_LC_4_3_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_5_LC_4_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_5_LC_4_3_2 (
            .in0(_gnd_net_),
            .in1(N__3515),
            .in2(N__3781),
            .in3(N__2576),
            .lcout(Pixel_RNOZ0Z_5),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_4_3_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_4_3_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_4_3_3 (
            .in0(_gnd_net_),
            .in1(N__2573),
            .in2(N__3506),
            .in3(N__3774),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_4_3_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_4_3_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_4_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THB_LC_4_3_4 (
            .in0(_gnd_net_),
            .in1(N__3494),
            .in2(_gnd_net_),
            .in3(N__2564),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0),
            .ltout(un2_x_if_generate_plus_mult1_un75_sum_cry_7_c_RNIU3THBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_1_LC_4_3_5.C_ON=1'b0;
    defparam Pixel_RNO_1_LC_4_3_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_1_LC_4_3_5.LUT_INIT=16'b0100111110110000;
    LogicCell40 Pixel_RNO_1_LC_4_3_5 (
            .in0(N__3463),
            .in1(N__2815),
            .in2(N__2561),
            .in3(N__2558),
            .lcout(un2_x_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI5UL6_5_LC_4_3_6.C_ON=1'b0;
    defparam x_RNI5UL6_5_LC_4_3_6.SEQ_MODE=4'b0000;
    defparam x_RNI5UL6_5_LC_4_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI5UL6_5_LC_4_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3684),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_3_LC_4_3_7.C_ON=1'b0;
    defparam Pixel_RNO_3_LC_4_3_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_3_LC_4_3_7.LUT_INIT=16'b1100001010001100;
    LogicCell40 Pixel_RNO_3_LC_4_3_7 (
            .in0(N__2858),
            .in1(N__2816),
            .in2(N__3467),
            .in3(N__2807),
            .lcout(un13lt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_5_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_5_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIQ64V_4_LC_4_5_2.C_ON=1'b0;
    defparam y_RNIQ64V_4_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam y_RNIQ64V_4_LC_4_5_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 y_RNIQ64V_4_LC_4_5_2 (
            .in0(N__2780),
            .in1(N__2741),
            .in2(N__2645),
            .in3(N__3056),
            .lcout(),
            .ltout(un1_ylto9_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIMA162_3_LC_4_5_3.C_ON=1'b0;
    defparam y_RNIMA162_3_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam y_RNIMA162_3_LC_4_5_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 y_RNIMA162_3_LC_4_5_3 (
            .in0(N__2663),
            .in1(N__3216),
            .in2(N__2792),
            .in3(N__3170),
            .lcout(un1_y),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_3_LC_4_6_0.C_ON=1'b0;
    defparam y_3_LC_4_6_0.SEQ_MODE=4'b1000;
    defparam y_3_LC_4_6_0.LUT_INIT=16'b0101000001111000;
    LogicCell40 y_3_LC_4_6_0 (
            .in0(N__2954),
            .in1(N__2789),
            .in2(N__3230),
            .in3(N__3016),
            .lcout(yZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3713),
            .ce(),
            .sr(_gnd_net_));
    defparam y_1_LC_4_6_1.C_ON=1'b0;
    defparam y_1_LC_4_6_1.SEQ_MODE=4'b1000;
    defparam y_1_LC_4_6_1.LUT_INIT=16'b0110011010101010;
    LogicCell40 y_1_LC_4_6_1 (
            .in0(N__2687),
            .in1(N__2955),
            .in2(_gnd_net_),
            .in3(N__2991),
            .lcout(yZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3713),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIGS3V_0_LC_4_6_2.C_ON=1'b0;
    defparam y_RNIGS3V_0_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam y_RNIGS3V_0_LC_4_6_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 y_RNIGS3V_0_LC_4_6_2 (
            .in0(N__2691),
            .in1(N__2779),
            .in2(N__2995),
            .in3(N__2740),
            .lcout(y_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIL6BN_9_LC_4_6_3.C_ON=1'b0;
    defparam y_RNIL6BN_9_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam y_RNIL6BN_9_LC_4_6_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 y_RNIL6BN_9_LC_4_6_3 (
            .in0(N__2686),
            .in1(N__3094),
            .in2(_gnd_net_),
            .in3(N__3130),
            .lcout(un1_ylto9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_2_LC_4_6_4.C_ON=1'b0;
    defparam y_2_LC_4_6_4.SEQ_MODE=4'b1000;
    defparam y_2_LC_4_6_4.LUT_INIT=16'b0101011100100000;
    LogicCell40 y_2_LC_4_6_4 (
            .in0(N__2953),
            .in1(N__3015),
            .in2(N__2657),
            .in3(N__3174),
            .lcout(yZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3713),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIM24V_9_LC_4_6_5.C_ON=1'b0;
    defparam y_RNIM24V_9_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam y_RNIM24V_9_LC_4_6_5.LUT_INIT=16'b0100000000000000;
    LogicCell40 y_RNIM24V_9_LC_4_6_5 (
            .in0(N__2639),
            .in1(N__3217),
            .in2(N__3183),
            .in3(N__3131),
            .lcout(),
            .ltout(y_12_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_RNIN6QD2_7_LC_4_6_6.C_ON=1'b0;
    defparam y_RNIN6QD2_7_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam y_RNIN6QD2_7_LC_4_6_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 y_RNIN6QD2_7_LC_4_6_6 (
            .in0(N__3095),
            .in1(N__3065),
            .in2(N__3059),
            .in3(N__3055),
            .lcout(y_12_8),
            .ltout(y_12_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_0_LC_4_6_7.C_ON=1'b0;
    defparam y_0_LC_4_6_7.SEQ_MODE=4'b1000;
    defparam y_0_LC_4_6_7.LUT_INIT=16'b0000001111001100;
    LogicCell40 y_0_LC_4_6_7 (
            .in0(_gnd_net_),
            .in1(N__2990),
            .in2(N__2999),
            .in3(N__2956),
            .lcout(yZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3713),
            .ce(),
            .sr(_gnd_net_));
    defparam x_0_LC_5_1_1.C_ON=1'b0;
    defparam x_0_LC_5_1_1.SEQ_MODE=4'b1000;
    defparam x_0_LC_5_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_0_LC_5_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2832),
            .lcout(xZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3718),
            .ce(),
            .sr(_gnd_net_));
    defparam x_1_LC_5_1_3.C_ON=1'b0;
    defparam x_1_LC_5_1_3.SEQ_MODE=4'b1000;
    defparam x_1_LC_5_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 x_1_LC_5_1_3 (
            .in0(_gnd_net_),
            .in1(N__2872),
            .in2(_gnd_net_),
            .in3(N__2833),
            .lcout(xZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3718),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNIRVNQ_9_LC_5_1_4.C_ON=1'b0;
    defparam x_RNIRVNQ_9_LC_5_1_4.SEQ_MODE=4'b0000;
    defparam x_RNIRVNQ_9_LC_5_1_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 x_RNIRVNQ_9_LC_5_1_4 (
            .in0(N__3935),
            .in1(N__3360),
            .in2(N__3413),
            .in3(N__3458),
            .lcout(),
            .ltout(un11_x_4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNID8R22_9_LC_5_1_5.C_ON=1'b0;
    defparam x_RNID8R22_9_LC_5_1_5.SEQ_MODE=4'b0000;
    defparam x_RNID8R22_9_LC_5_1_5.LUT_INIT=16'b1100000000000000;
    LogicCell40 x_RNID8R22_9_LC_5_1_5 (
            .in0(_gnd_net_),
            .in1(N__3638),
            .in2(N__2972),
            .in3(N__3479),
            .lcout(x_RNID8R22Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI6ANQ_1_LC_5_1_7.C_ON=1'b0;
    defparam x_RNI6ANQ_1_LC_5_1_7.SEQ_MODE=4'b0000;
    defparam x_RNI6ANQ_1_LC_5_1_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 x_RNI6ANQ_1_LC_5_1_7 (
            .in0(N__2887),
            .in1(N__2871),
            .in2(N__2857),
            .in3(N__2831),
            .lcout(un11_x_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_LC_5_2_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_LC_5_2_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_LC_5_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_LC_5_2_0 (
            .in0(_gnd_net_),
            .in1(N__3405),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(un2_x_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_5_2_1.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_5_2_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_5_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_5_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3485),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(un2_x_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_5_2_2.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_5_2_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_5_2_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46N8_LC_5_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3482),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI46NZ0Z8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_9_LC_5_2_3.C_ON=1'b0;
    defparam Pixel_RNO_9_LC_5_2_3.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_9_LC_5_2_3.LUT_INIT=16'b0000000000000010;
    LogicCell40 Pixel_RNO_9_LC_5_2_3 (
            .in0(N__3634),
            .in1(N__3478),
            .in2(N__3461),
            .in3(N__3933),
            .lcout(un4_xlt9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI81M6_8_LC_5_2_4.C_ON=1'b0;
    defparam x_RNI81M6_8_LC_5_2_4.SEQ_MODE=4'b0000;
    defparam x_RNI81M6_8_LC_5_2_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI81M6_8_LC_5_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3358),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI92M6_9_LC_5_2_5.C_ON=1'b0;
    defparam x_RNI92M6_9_LC_5_2_5.SEQ_MODE=4'b0000;
    defparam x_RNI92M6_9_LC_5_2_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 x_RNI92M6_9_LC_5_2_5 (
            .in0(N__3406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSyncZ0_LC_5_2_7.C_ON=1'b0;
    defparam HSyncZ0_LC_5_2_7.SEQ_MODE=4'b1000;
    defparam HSyncZ0_LC_5_2_7.LUT_INIT=16'b1111101110111011;
    LogicCell40 HSyncZ0_LC_5_2_7 (
            .in0(N__3407),
            .in1(N__3329),
            .in2(N__3685),
            .in3(N__3934),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3717),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_RNO_0_LC_5_3_0.C_ON=1'b1;
    defparam HSync_RNO_0_LC_5_3_0.SEQ_MODE=4'b0000;
    defparam HSync_RNO_0_LC_5_3_0.LUT_INIT=16'b0000000000001111;
    LogicCell40 HSync_RNO_0_LC_5_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3365),
            .in3(N__3978),
            .lcout(un1_xlto9_0),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_5_3_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_5_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTH_LC_5_3_1 (
            .in0(_gnd_net_),
            .in1(N__3323),
            .in2(_gnd_net_),
            .in3(N__3317),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_4_c_RNIKSTHZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_5_3_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_5_3_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_5_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20K_LC_5_3_2 (
            .in0(_gnd_net_),
            .in1(N__3314),
            .in2(N__3305),
            .in3(N__3236),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_5_c_RNIG20KZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_5_3_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_5_3_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_5_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_6_c_RNI7HQG1_LC_5_3_3 (
            .in0(N__3613),
            .in1(N__3521),
            .in2(N__3542),
            .in3(N__3551),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_5_3_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_5_3_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_5_3_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_LC_5_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3548),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0),
            .ltout(un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_5_3_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_5_3_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_5_3_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un47_sum_cry_7_c_RNIE0BB_0_LC_5_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3545),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_5_3_6.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_5_3_6.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_5_3_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEH_LC_5_3_6 (
            .in0(_gnd_net_),
            .in1(N__3532),
            .in2(_gnd_net_),
            .in3(N__3538),
            .lcout(un2_x_if_generate_plus_mult1_un40_sum_cry_4_c_RNI8CEHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0 (
            .in0(_gnd_net_),
            .in1(N__3680),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_5_4_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_5_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVB3_LC_5_4_1 (
            .in0(_gnd_net_),
            .in1(N__3793),
            .in2(N__3761),
            .in3(N__3509),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_4_c_RNIQMVBZ0Z3),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_5_4_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_5_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIM0465_LC_5_4_2 (
            .in0(_gnd_net_),
            .in1(N__3809),
            .in2(N__3890),
            .in3(N__3497),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_5_c_RNIMZ0Z0465),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_5_4_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_5_4_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_5_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFKBHB_LC_5_4_3 (
            .in0(N__3782),
            .in1(N__3794),
            .in2(N__3857),
            .in3(N__3488),
            .lcout(un2_x_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_5_4_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_5_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABU5_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__3827),
            .in2(_gnd_net_),
            .in3(N__3785),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_cry_7_c_RNIVABUZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI6VL6_6_LC_5_4_6.C_ON=1'b0;
    defparam x_RNI6VL6_6_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam x_RNI6VL6_6_LC_5_4_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI6VL6_6_LC_5_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3944),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSyncZ0_LC_6_2_3.C_ON=1'b0;
    defparam VSyncZ0_LC_6_2_3.SEQ_MODE=4'b1000;
    defparam VSyncZ0_LC_6_2_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 VSyncZ0_LC_6_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3752),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3719),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNICUBD_5_LC_6_3_0.C_ON=1'b1;
    defparam x_RNICUBD_5_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam x_RNICUBD_5_LC_6_3_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 x_RNICUBD_5_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(N__3979),
            .in2(_gnd_net_),
            .in3(N__3686),
            .lcout(un11_x_4),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_6_3_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_6_3_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_6_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJ_LC_6_3_1 (
            .in0(_gnd_net_),
            .in1(N__3623),
            .in2(N__3590),
            .in3(N__3617),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_4_c_RNIV4GJZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_6_3_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_6_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PU_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(N__3614),
            .in2(N__3602),
            .in3(N__3593),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC2PUZ0),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_6_3_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_6_3_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_6_3_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_6_c_RNIS49J2_LC_6_3_3 (
            .in0(N__3877),
            .in1(N__3589),
            .in2(N__3575),
            .in3(N__3566),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_6_3_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_6_3_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_6_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_LC_6_3_4 (
            .in0(_gnd_net_),
            .in1(N__3563),
            .in2(_gnd_net_),
            .in3(N__3557),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1),
            .ltout(un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCIZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_6_3_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_6_3_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un54_sum_cry_7_c_RNIJQCI1_0_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3554),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam x_RNI70M6_7_LC_6_3_6.C_ON=1'b0;
    defparam x_RNI70M6_7_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam x_RNI70M6_7_LC_6_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 x_RNI70M6_7_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3980),
            .lcout(un2_x_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0 (
            .in0(_gnd_net_),
            .in1(N__3943),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_4_1.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17P02_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(N__3844),
            .in2(N__3899),
            .in3(N__3881),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_4_c_RNI17PZ0Z02),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_4_2.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_4_2.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKD2_LC_6_4_2 (
            .in0(_gnd_net_),
            .in1(N__3878),
            .in2(N__3866),
            .in3(N__3848),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_5_c_RNIQDKDZ0Z2),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_4_3.C_ON=1'b1;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_4_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_6_c_RNIE41K5_LC_6_4_3 (
            .in0(N__3808),
            .in1(N__3845),
            .in2(N__3836),
            .in3(N__3821),
            .lcout(un2_x_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un2_x_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un2_x_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_4_4.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_LC_6_4_4 (
            .in0(_gnd_net_),
            .in1(N__3818),
            .in2(_gnd_net_),
            .in3(N__3812),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2),
            .ltout(un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2RZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_4_5.C_ON=1'b0;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_4_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un2_x_if_generate_plus_mult1_un61_sum_cry_7_c_RNI6N2R2_0_LC_6_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3797),
            .in3(_gnd_net_),
            .lcout(un2_x_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
