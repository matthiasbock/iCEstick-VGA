// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 19 2015 15:42:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__11180;
    wire N__11179;
    wire N__11178;
    wire N__11171;
    wire N__11170;
    wire N__11169;
    wire N__11162;
    wire N__11161;
    wire N__11160;
    wire N__11153;
    wire N__11152;
    wire N__11151;
    wire N__11144;
    wire N__11143;
    wire N__11142;
    wire N__11135;
    wire N__11134;
    wire N__11133;
    wire N__11126;
    wire N__11125;
    wire N__11124;
    wire N__11107;
    wire N__11106;
    wire N__11105;
    wire N__11104;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11074;
    wire N__11067;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11048;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10962;
    wire N__10959;
    wire N__10958;
    wire N__10955;
    wire N__10950;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10934;
    wire N__10933;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10921;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10882;
    wire N__10879;
    wire N__10872;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10829;
    wire N__10824;
    wire N__10821;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10810;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10772;
    wire N__10765;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10728;
    wire N__10727;
    wire N__10726;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10705;
    wire N__10700;
    wire N__10697;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10681;
    wire N__10678;
    wire N__10677;
    wire N__10676;
    wire N__10675;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10659;
    wire N__10656;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10645;
    wire N__10640;
    wire N__10637;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10617;
    wire N__10610;
    wire N__10607;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10578;
    wire N__10577;
    wire N__10576;
    wire N__10575;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10558;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10516;
    wire N__10513;
    wire N__10506;
    wire N__10501;
    wire N__10498;
    wire N__10493;
    wire N__10492;
    wire N__10489;
    wire N__10482;
    wire N__10479;
    wire N__10474;
    wire N__10469;
    wire N__10466;
    wire N__10461;
    wire N__10450;
    wire N__10449;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10443;
    wire N__10442;
    wire N__10439;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10431;
    wire N__10430;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10422;
    wire N__10419;
    wire N__10412;
    wire N__10407;
    wire N__10400;
    wire N__10395;
    wire N__10388;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10364;
    wire N__10363;
    wire N__10360;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10356;
    wire N__10355;
    wire N__10354;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10347;
    wire N__10346;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10316;
    wire N__10311;
    wire N__10306;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10280;
    wire N__10277;
    wire N__10272;
    wire N__10265;
    wire N__10262;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10247;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10219;
    wire N__10218;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10213;
    wire N__10212;
    wire N__10211;
    wire N__10210;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10193;
    wire N__10192;
    wire N__10191;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10176;
    wire N__10175;
    wire N__10172;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10134;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10119;
    wire N__10116;
    wire N__10111;
    wire N__10108;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10092;
    wire N__10087;
    wire N__10078;
    wire N__10077;
    wire N__10076;
    wire N__10075;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10065;
    wire N__10064;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10047;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10035;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10027;
    wire N__10022;
    wire N__10019;
    wire N__10012;
    wire N__10009;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9942;
    wire N__9937;
    wire N__9934;
    wire N__9933;
    wire N__9928;
    wire N__9925;
    wire N__9924;
    wire N__9923;
    wire N__9922;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9905;
    wire N__9902;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9859;
    wire N__9856;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9813;
    wire N__9812;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9759;
    wire N__9758;
    wire N__9755;
    wire N__9754;
    wire N__9753;
    wire N__9752;
    wire N__9749;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9720;
    wire N__9719;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9690;
    wire N__9685;
    wire N__9680;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9639;
    wire N__9638;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9586;
    wire N__9585;
    wire N__9584;
    wire N__9581;
    wire N__9580;
    wire N__9579;
    wire N__9576;
    wire N__9569;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9563;
    wire N__9562;
    wire N__9561;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9546;
    wire N__9545;
    wire N__9544;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9513;
    wire N__9508;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9444;
    wire N__9443;
    wire N__9440;
    wire N__9439;
    wire N__9436;
    wire N__9435;
    wire N__9432;
    wire N__9423;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9111;
    wire N__9110;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9091;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9072;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9039;
    wire N__9036;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__8997;
    wire N__8996;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8954;
    wire N__8949;
    wire N__8946;
    wire N__8945;
    wire N__8942;
    wire N__8933;
    wire N__8930;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8920;
    wire N__8915;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8887;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8875;
    wire N__8872;
    wire N__8865;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8828;
    wire N__8827;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8813;
    wire N__8812;
    wire N__8809;
    wire N__8808;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8778;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8760;
    wire N__8755;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8747;
    wire N__8742;
    wire N__8741;
    wire N__8738;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8714;
    wire N__8701;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8603;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8573;
    wire N__8570;
    wire N__8565;
    wire N__8560;
    wire N__8559;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8505;
    wire N__8504;
    wire N__8501;
    wire N__8500;
    wire N__8499;
    wire N__8496;
    wire N__8487;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8470;
    wire N__8469;
    wire N__8466;
    wire N__8465;
    wire N__8462;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8429;
    wire N__8416;
    wire N__8415;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8410;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8403;
    wire N__8402;
    wire N__8399;
    wire N__8394;
    wire N__8385;
    wire N__8378;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8366;
    wire N__8361;
    wire N__8358;
    wire N__8353;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8341;
    wire N__8340;
    wire N__8339;
    wire N__8334;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8308;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8288;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8225;
    wire N__8224;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8203;
    wire N__8196;
    wire N__8195;
    wire N__8192;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8167;
    wire N__8158;
    wire N__8157;
    wire N__8156;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8139;
    wire N__8134;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8128;
    wire N__8123;
    wire N__8120;
    wire N__8113;
    wire N__8104;
    wire N__8103;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8092;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8065;
    wire N__8062;
    wire N__8061;
    wire N__8060;
    wire N__8059;
    wire N__8056;
    wire N__8049;
    wire N__8048;
    wire N__8047;
    wire N__8046;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8034;
    wire N__8033;
    wire N__8030;
    wire N__8023;
    wire N__8020;
    wire N__8019;
    wire N__8018;
    wire N__8017;
    wire N__8014;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7993;
    wire N__7990;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7965;
    wire N__7962;
    wire N__7961;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7943;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7933;
    wire N__7932;
    wire N__7931;
    wire N__7930;
    wire N__7927;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7902;
    wire N__7893;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7855;
    wire N__7854;
    wire N__7853;
    wire N__7850;
    wire N__7849;
    wire N__7846;
    wire N__7837;
    wire N__7832;
    wire N__7829;
    wire N__7824;
    wire N__7813;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7805;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7782;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7677;
    wire N__7674;
    wire N__7673;
    wire N__7672;
    wire N__7669;
    wire N__7668;
    wire N__7667;
    wire N__7666;
    wire N__7659;
    wire N__7654;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7636;
    wire N__7635;
    wire N__7626;
    wire N__7623;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7572;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7555;
    wire N__7552;
    wire N__7551;
    wire N__7550;
    wire N__7545;
    wire N__7542;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7521;
    wire N__7520;
    wire N__7519;
    wire N__7518;
    wire N__7517;
    wire N__7516;
    wire N__7511;
    wire N__7510;
    wire N__7509;
    wire N__7508;
    wire N__7507;
    wire N__7506;
    wire N__7499;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7484;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7466;
    wire N__7463;
    wire N__7452;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7425;
    wire N__7422;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7347;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7326;
    wire N__7323;
    wire N__7322;
    wire N__7319;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7307;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7212;
    wire N__7211;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7120;
    wire N__7119;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7035;
    wire N__7030;
    wire N__7027;
    wire N__7026;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7016;
    wire N__7011;
    wire N__7008;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6996;
    wire N__6995;
    wire N__6994;
    wire N__6985;
    wire N__6982;
    wire N__6977;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6954;
    wire N__6949;
    wire N__6946;
    wire N__6945;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6912;
    wire N__6911;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6903;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6888;
    wire N__6885;
    wire N__6874;
    wire N__6873;
    wire N__6872;
    wire N__6869;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6846;
    wire N__6843;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6820;
    wire N__6819;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6802;
    wire N__6799;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6769;
    wire N__6768;
    wire N__6763;
    wire N__6762;
    wire N__6759;
    wire N__6758;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6736;
    wire N__6735;
    wire N__6734;
    wire N__6733;
    wire N__6730;
    wire N__6729;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6691;
    wire N__6690;
    wire N__6689;
    wire N__6686;
    wire N__6685;
    wire N__6684;
    wire N__6681;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6649;
    wire N__6646;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6638;
    wire N__6637;
    wire N__6632;
    wire N__6627;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6519;
    wire N__6518;
    wire N__6515;
    wire N__6514;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6489;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6423;
    wire N__6420;
    wire N__6419;
    wire N__6418;
    wire N__6411;
    wire N__6408;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6300;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6263;
    wire N__6262;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6249;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6230;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6194;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6181;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6130;
    wire N__6127;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6060;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5982;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5919;
    wire N__5918;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5906;
    wire N__5899;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5887;
    wire N__5884;
    wire N__5879;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5853;
    wire N__5848;
    wire N__5845;
    wire N__5844;
    wire N__5839;
    wire N__5836;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5757;
    wire N__5756;
    wire N__5751;
    wire N__5748;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5701;
    wire N__5698;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5690;
    wire N__5689;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5675;
    wire N__5668;
    wire N__5667;
    wire N__5662;
    wire N__5661;
    wire N__5660;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5638;
    wire N__5637;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5629;
    wire N__5624;
    wire N__5619;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5566;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5484;
    wire N__5483;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5471;
    wire N__5464;
    wire N__5455;
    wire N__5452;
    wire N__5451;
    wire N__5450;
    wire N__5449;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5440;
    wire N__5435;
    wire N__5432;
    wire N__5425;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5358;
    wire N__5357;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5274;
    wire N__5273;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5261;
    wire N__5258;
    wire N__5251;
    wire N__5248;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5231;
    wire N__5228;
    wire N__5221;
    wire N__5218;
    wire N__5217;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5200;
    wire N__5197;
    wire N__5188;
    wire N__5185;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5179;
    wire N__5178;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5160;
    wire N__5157;
    wire N__5146;
    wire N__5143;
    wire N__5142;
    wire N__5141;
    wire N__5140;
    wire N__5139;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5127;
    wire N__5122;
    wire N__5119;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5077;
    wire N__5074;
    wire N__5073;
    wire N__5070;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5051;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5019;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5011;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4996;
    wire N__4993;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4936;
    wire N__4933;
    wire N__4932;
    wire N__4921;
    wire N__4918;
    wire N__4917;
    wire N__4914;
    wire N__4913;
    wire N__4910;
    wire N__4909;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4886;
    wire N__4883;
    wire N__4878;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4825;
    wire N__4824;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire \Clock50MHz.PixelClock ;
    wire Clock12MHz_c;
    wire VCCG0;
    wire GNDG0;
    wire bfn_4_3_0_;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire bfn_4_4_0_;
    wire un5_beamx_3;
    wire un5_beamx_4_cascade_;
    wire beamY_RNIMA24P1Z0Z_5;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_;
    wire un3_beamx_5_cascade_;
    wire un3_beamx_7_cascade_;
    wire beamX_RNI5457Z0Z_5_cascade_;
    wire un13_beamylto2_0_cascade_;
    wire bfn_4_9_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_4_10_0_;
    wire un8_beamx_cry_9;
    wire N_7_1_cascade_;
    wire g2_1_0;
    wire N_14_cascade_;
    wire beamY_fast_RNIG57DZ0Z_4_cascade_;
    wire un5_visibley_c5_cascade_;
    wire un21_beamy_cry_2_c_RNICOZ0Z83;
    wire un21_beamy_cry_3_c_RNIERZ0Z93;
    wire un21_beamy_cry_1_c_RNIALZ0Z73;
    wire un5_visibley_ac0_11_d_cascade_;
    wire beamY_fastZ0Z_8;
    wire beamY_fastZ0Z_4;
    wire beamY_fast_RNI24GAZ0Z_2_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cascade_;
    wire beamY_RNI2GUN3Z0Z_9;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_;
    wire beamY_RNI2GUN3_0Z0Z_9;
    wire d_i4_mux;
    wire beamY_RNICDD7FZ0Z_5_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3;
    wire beamY_RNIUBM4FZ0Z_7_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_c5;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i;
    wire beamY_RNIID28F1_0Z0Z_3_cascade_;
    wire un18_beamylt5_0;
    wire un18_beamylto9_2_cascade_;
    wire beamY_RNIID28F1Z0Z_3;
    wire bfn_5_9_0_;
    wire beamXZ0Z_1;
    wire un5_visiblex_cry_0;
    wire beamXZ0Z_2;
    wire un5_visiblex_cry_1;
    wire beamXZ0Z_3;
    wire un5_visiblex_cry_2;
    wire beamXZ0Z_4;
    wire un5_visiblex_cry_3;
    wire beamXZ0Z_5;
    wire un5_visiblex_cry_4;
    wire beamXZ0Z_6;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire beamXZ0Z_8;
    wire bfn_5_10_0_;
    wire beamXZ0Z_9;
    wire un5_visiblex_cry_8;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_;
    wire g0_0_2_0;
    wire bfn_5_11_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_0;
    wire bfn_5_12_0_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_1;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_;
    wire bfn_5_13_0_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_i_8;
    wire beamY_fast_RNIM4P7_0Z0Z_2_cascade_;
    wire beamY_fast_RNIO71DZ0Z_3;
    wire beamY_fastZ0Z_2;
    wire beamY_fast_RNIM4P7Z0Z_2_cascade_;
    wire beamY_fastZ0Z_3;
    wire bfn_6_5_0_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire beamY_fast_RNIG57D_0Z0Z_4;
    wire beamY_fast_RNI45FMZ0Z_7;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_;
    wire beamY_RNIK0NV_0Z0Z_9;
    wire un5_visibley_ac0_11_d;
    wire un5_visibley_c7_cascade_;
    wire un21_beamy_cry_8_c_RNIOAFZ0Z3;
    wire un21_beamy_cry_6_c_RNIK4DZ0Z3;
    wire un21_beamy_cry_7_c_RNIM7EZ0Z3;
    wire un5_visibley_c5;
    wire beamY_fastZ0Z_9;
    wire font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux;
    wire font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i;
    wire beamY_RNI779U3Z0Z_5;
    wire beamY_RNIUBM4FZ0Z_7;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_c4;
    wire beamY_RNI9N7M7Z0Z_5;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_c5;
    wire beamY_RNI5F8A81Z0Z_3_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_;
    wire beamY_RNIKUC181_0Z0Z_5;
    wire beamY_RNIKPNA02Z0Z_5;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_c4;
    wire font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0;
    wire font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i;
    wire bfn_6_9_0_;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7;
    wire bfn_6_10_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO;
    wire font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_;
    wire un22_visibleylt9_0_0_0;
    wire bfn_6_11_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_i;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_;
    wire un5_visiblex_cry_7_c_RNIVZ0Z952;
    wire un5_visiblex_i_24;
    wire bfn_6_12_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_;
    wire font_un19_pixel_if_generate_plus_mult1_un40_sum_i;
    wire bfn_6_13_0_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i;
    wire bfn_7_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_0;
    wire bfn_7_4_0_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_7;
    wire bfn_7_5_0_;
    wire beamY_RNI9KEQ_0Z0Z_8;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_axb_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_7;
    wire beamY_fastZ0Z_7;
    wire un5_visibley_c6_0_0_0;
    wire un11_visibleylto9_1_cascade_;
    wire un11_visibleylto9_4_cascade_;
    wire un21_beamy_cry_5_c_RNII1CZ0Z3;
    wire beamY_fastZ0Z_6;
    wire un5_visibley_c6_0_0;
    wire un21_beamy_cry_4_c_RNIGUAZ0Z3;
    wire beamY_fastZ0Z_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_axb_3;
    wire beamY_RNIECTA3Z0Z_8_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1;
    wire un1_beamylto9_2;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0;
    wire beamY_RNIECTA3Z0Z_8;
    wire font_un42_pixel_if_generate_plus_mult1_un47_sum_c5;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_;
    wire font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2;
    wire un1_beamylto9_1;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5;
    wire Pixel_1_esr_RNOZ0Z_60;
    wire g1_0_cascade_;
    wire un1_beamxlt10_0;
    wire beamXZ0Z_7;
    wire font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0;
    wire beamY_RNIAJLT9AZ0Z_3;
    wire r_i1_mux_cascade_;
    wire font_un78_pixellto3;
    wire Pixel_3_sqmuxa_1_1_cascade_;
    wire G_25_i_a8_0_0;
    wire Pixel_7_sqmuxa_1_cascade_;
    wire g0_0_0_1;
    wire g1;
    wire g0_0_4_0_cascade_;
    wire N_11;
    wire g0_0_2;
    wire Pixel_3_sqmuxa_1_1;
    wire N_7_0;
    wire G_25_i_a8_1_1;
    wire G_25_i_o8_0_2;
    wire Pixel_7_sqmuxa_1;
    wire bfn_7_11_0_;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5;
    wire g0_10_0_cascade_;
    wire bfn_7_12_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_i;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72;
    wire font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i_8;
    wire Pixel_9_sn_N_7_mux_1_tz;
    wire un16_visibleylt9_0_cascade_;
    wire un16_visibley_4;
    wire un28_visibleylt9_0;
    wire Pixel_7_sqmuxa_3_0_1;
    wire un22_visibley_3;
    wire un22_visibleylt9_0_cascade_;
    wire un22_visibley_2;
    wire un22_visibley;
    wire un1_beamY_if_generate_plus_mult1_un54_sum;
    wire bfn_8_4_0_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6;
    wire bfn_8_5_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_7;
    wire beamY_fast_RNI1QVSZ0Z_9;
    wire un1_beamY_if_generate_plus_mult1_un47_sum;
    wire un1_beamY_if_generate_plus_mult1_un40_sum;
    wire font_un42_pixel_if_generate_plus_mult1_un47_sum_c4;
    wire un5_visibley_c2;
    wire beamX_RNI5457Z0Z_5;
    wire un5_beamx;
    wire un1_beamY_if_generate_plus_mult1_un68_sum;
    wire beamYZ0Z_3;
    wire un4_beamylt6;
    wire un4_beamylt6_cascade_;
    wire beamYZ0Z_4;
    wire beamYZ0Z_8;
    wire un4_beamylt8_0_cascade_;
    wire beamYZ0Z_9;
    wire CONSTANT_ONE_NET;
    wire beamYZ0Z_2;
    wire beamYZ0Z_5;
    wire un8_beamylto9_1;
    wire beamYZ0Z_6;
    wire beamYZ0Z_7;
    wire Pixel_1_sqmuxa_i_cascade_;
    wire un1_beamx;
    wire HSync_c;
    wire un4_beamy_0;
    wire un18_beamylt10_0;
    wire beamXZ0Z_10;
    wire un8_beamy;
    wire un15_beamy_2;
    wire un1_beamx_2;
    wire un13_beamylt10_0;
    wire un15_beamy_2_cascade_;
    wire un11_visibley;
    wire un27lt10;
    wire un1_visiblex_27;
    wire Pixel_9_sqmuxa_0_cascade_;
    wire Pixel_9_sqmuxa;
    wire g0_i_o4_3;
    wire Pixel_9_u_ns_sn;
    wire N_163_cascade_;
    wire Pixel_c;
    wire Pixel_1_sqmuxa_i_0;
    wire g1_0_0;
    wire g0_0_4;
    wire G_25_i_a8_2_0;
    wire g0_0_5_cascade_;
    wire G_25_i_3_0;
    wire N_20;
    wire G_25_i_2_0_cascade_;
    wire G_25_i_0;
    wire Pixel_9_u_ns_rn_0;
    wire g2_1;
    wire bfn_8_10_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_i;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_;
    wire g1_0_1_1;
    wire font_un19_pixel_0_0_0_23_cascade_;
    wire g2_0;
    wire g1_0_2;
    wire font_un237_pixel_6_ns_1_0_0_cascade_;
    wire g1_2_0;
    wire font_un237_pixel_0_0;
    wire g2_cascade_;
    wire font_un83_pixel_0_0;
    wire font_un19_pixel_23;
    wire font_un19_pixel_23_cascade_;
    wire font_un160_pixel_6_1;
    wire g0_1_0_cascade_;
    wire g3_0_0;
    wire bfn_8_12_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum;
    wire font_un19_pixel_if_generate_plus_mult1_un54_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6;
    wire g0_i_o4_2;
    wire bfn_9_6_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6;
    wire un28lto4_1_cascade_;
    wire Pixel_1_esr_RNOZ0Z_62;
    wire un28lt10_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0;
    wire un28_0_1;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0;
    wire beamY_i_2;
    wire un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5;
    wire beamY_RNIJ0DBZ0Z_9;
    wire VSync_c;
    wire PixelClock_g;
    wire g1_1_cascade_;
    wire Pixel_1_esr_RNOZ0Z_39;
    wire N_1304_0_cascade_;
    wire g1_0_1;
    wire N_17_cascade_;
    wire G_25_i_a8_1;
    wire g1_3_cascade_;
    wire N_1302_0_0_0_cascade_;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9;
    wire beamXZ0Z_0;
    wire N_159_0_0_cascade_;
    wire N_156_0;
    wire font_un314_pixel_0;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1;
    wire g1_3_0_0;
    wire un28lto1;
    wire beamYZ0Z_0;
    wire font_un42_pixel_23;
    wire N_1303_0_0;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum;
    wire bfn_9_11_0_;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5;
    wire font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i;
    wire un1_visiblex_24;
    wire font_un19_pixel_if_generate_plus_mult1_un61_sum_i;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__4687),
            .RESETB(N__9094),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__11180),
            .DIN(N__11179),
            .DOUT(N__11178),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__11180),
            .PADOUT(N__11179),
            .PADIN(N__11178),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9223),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__11171),
            .DIN(N__11170),
            .DOUT(N__11169),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__11171),
            .PADOUT(N__11170),
            .PADIN(N__11169),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9855),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__11162),
            .DIN(N__11161),
            .DOUT(N__11160),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__11162),
            .PADOUT(N__11161),
            .PADIN(N__11160),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8676),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__11153),
            .DIN(N__11152),
            .DOUT(N__11151),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__11153),
            .PADOUT(N__11152),
            .PADIN(N__11151),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8683),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__11144),
            .DIN(N__11143),
            .DOUT(N__11142),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__11144),
            .PADOUT(N__11143),
            .PADIN(N__11142),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__11135),
            .DIN(N__11134),
            .DOUT(N__11133),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__11135),
            .PADOUT(N__11134),
            .PADIN(N__11133),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9859),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__11126),
            .DIN(N__11125),
            .DOUT(N__11124),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__11126),
            .PADOUT(N__11125),
            .PADIN(N__11124),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2546 (
            .O(N__11107),
            .I(N__11100));
    InMux I__2545 (
            .O(N__11106),
            .I(N__11097));
    InMux I__2544 (
            .O(N__11105),
            .I(N__11092));
    InMux I__2543 (
            .O(N__11104),
            .I(N__11089));
    InMux I__2542 (
            .O(N__11103),
            .I(N__11086));
    LocalMux I__2541 (
            .O(N__11100),
            .I(N__11081));
    LocalMux I__2540 (
            .O(N__11097),
            .I(N__11081));
    InMux I__2539 (
            .O(N__11096),
            .I(N__11078));
    InMux I__2538 (
            .O(N__11095),
            .I(N__11075));
    LocalMux I__2537 (
            .O(N__11092),
            .I(N__11067));
    LocalMux I__2536 (
            .O(N__11089),
            .I(N__11067));
    LocalMux I__2535 (
            .O(N__11086),
            .I(N__11067));
    Span4Mux_h I__2534 (
            .O(N__11081),
            .I(N__11062));
    LocalMux I__2533 (
            .O(N__11078),
            .I(N__11062));
    LocalMux I__2532 (
            .O(N__11075),
            .I(N__11059));
    InMux I__2531 (
            .O(N__11074),
            .I(N__11056));
    Span4Mux_h I__2530 (
            .O(N__11067),
            .I(N__11053));
    Span4Mux_v I__2529 (
            .O(N__11062),
            .I(N__11048));
    Span4Mux_v I__2528 (
            .O(N__11059),
            .I(N__11048));
    LocalMux I__2527 (
            .O(N__11056),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2526 (
            .O(N__11053),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2525 (
            .O(N__11048),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum));
    InMux I__2524 (
            .O(N__11041),
            .I(N__11038));
    LocalMux I__2523 (
            .O(N__11038),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0));
    InMux I__2522 (
            .O(N__11035),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__2521 (
            .O(N__11032),
            .I(N__11028));
    InMux I__2520 (
            .O(N__11031),
            .I(N__11025));
    LocalMux I__2519 (
            .O(N__11028),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0));
    LocalMux I__2518 (
            .O(N__11025),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0));
    CascadeMux I__2517 (
            .O(N__11020),
            .I(N__11017));
    InMux I__2516 (
            .O(N__11017),
            .I(N__11014));
    LocalMux I__2515 (
            .O(N__11014),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96));
    InMux I__2514 (
            .O(N__11011),
            .I(N__11008));
    LocalMux I__2513 (
            .O(N__11008),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0));
    InMux I__2512 (
            .O(N__11005),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__2511 (
            .O(N__11002),
            .I(N__10999));
    LocalMux I__2510 (
            .O(N__10999),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9));
    CascadeMux I__2509 (
            .O(N__10996),
            .I(N__10992));
    CascadeMux I__2508 (
            .O(N__10995),
            .I(N__10989));
    InMux I__2507 (
            .O(N__10992),
            .I(N__10984));
    InMux I__2506 (
            .O(N__10989),
            .I(N__10984));
    LocalMux I__2505 (
            .O(N__10984),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5));
    InMux I__2504 (
            .O(N__10981),
            .I(N__10978));
    LocalMux I__2503 (
            .O(N__10978),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__2502 (
            .O(N__10975),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__2501 (
            .O(N__10972),
            .I(N__10969));
    LocalMux I__2500 (
            .O(N__10969),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__2499 (
            .O(N__10966),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__2498 (
            .O(N__10963),
            .I(N__10959));
    InMux I__2497 (
            .O(N__10962),
            .I(N__10955));
    InMux I__2496 (
            .O(N__10959),
            .I(N__10950));
    InMux I__2495 (
            .O(N__10958),
            .I(N__10950));
    LocalMux I__2494 (
            .O(N__10955),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0));
    LocalMux I__2493 (
            .O(N__10950),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0));
    InMux I__2492 (
            .O(N__10945),
            .I(N__10938));
    InMux I__2491 (
            .O(N__10944),
            .I(N__10935));
    InMux I__2490 (
            .O(N__10943),
            .I(N__10929));
    InMux I__2489 (
            .O(N__10942),
            .I(N__10926));
    CascadeMux I__2488 (
            .O(N__10941),
            .I(N__10921));
    LocalMux I__2487 (
            .O(N__10938),
            .I(N__10916));
    LocalMux I__2486 (
            .O(N__10935),
            .I(N__10916));
    CascadeMux I__2485 (
            .O(N__10934),
            .I(N__10913));
    CascadeMux I__2484 (
            .O(N__10933),
            .I(N__10910));
    CascadeMux I__2483 (
            .O(N__10932),
            .I(N__10907));
    LocalMux I__2482 (
            .O(N__10929),
            .I(N__10904));
    LocalMux I__2481 (
            .O(N__10926),
            .I(N__10901));
    InMux I__2480 (
            .O(N__10925),
            .I(N__10896));
    InMux I__2479 (
            .O(N__10924),
            .I(N__10896));
    InMux I__2478 (
            .O(N__10921),
            .I(N__10893));
    Span4Mux_v I__2477 (
            .O(N__10916),
            .I(N__10890));
    InMux I__2476 (
            .O(N__10913),
            .I(N__10887));
    InMux I__2475 (
            .O(N__10910),
            .I(N__10882));
    InMux I__2474 (
            .O(N__10907),
            .I(N__10882));
    Span4Mux_h I__2473 (
            .O(N__10904),
            .I(N__10879));
    Span4Mux_v I__2472 (
            .O(N__10901),
            .I(N__10872));
    LocalMux I__2471 (
            .O(N__10896),
            .I(N__10872));
    LocalMux I__2470 (
            .O(N__10893),
            .I(N__10872));
    Odrv4 I__2469 (
            .O(N__10890),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    LocalMux I__2468 (
            .O(N__10887),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    LocalMux I__2467 (
            .O(N__10882),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    Odrv4 I__2466 (
            .O(N__10879),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    Odrv4 I__2465 (
            .O(N__10872),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    CascadeMux I__2464 (
            .O(N__10861),
            .I(N__10858));
    InMux I__2463 (
            .O(N__10858),
            .I(N__10855));
    LocalMux I__2462 (
            .O(N__10855),
            .I(N__10852));
    Odrv12 I__2461 (
            .O(N__10852),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i));
    CascadeMux I__2460 (
            .O(N__10849),
            .I(N__10840));
    InMux I__2459 (
            .O(N__10848),
            .I(N__10837));
    InMux I__2458 (
            .O(N__10847),
            .I(N__10833));
    InMux I__2457 (
            .O(N__10846),
            .I(N__10830));
    InMux I__2456 (
            .O(N__10845),
            .I(N__10824));
    InMux I__2455 (
            .O(N__10844),
            .I(N__10824));
    InMux I__2454 (
            .O(N__10843),
            .I(N__10821));
    InMux I__2453 (
            .O(N__10840),
            .I(N__10817));
    LocalMux I__2452 (
            .O(N__10837),
            .I(N__10814));
    InMux I__2451 (
            .O(N__10836),
            .I(N__10811));
    LocalMux I__2450 (
            .O(N__10833),
            .I(N__10805));
    LocalMux I__2449 (
            .O(N__10830),
            .I(N__10805));
    InMux I__2448 (
            .O(N__10829),
            .I(N__10802));
    LocalMux I__2447 (
            .O(N__10824),
            .I(N__10799));
    LocalMux I__2446 (
            .O(N__10821),
            .I(N__10796));
    InMux I__2445 (
            .O(N__10820),
            .I(N__10793));
    LocalMux I__2444 (
            .O(N__10817),
            .I(N__10790));
    Span4Mux_v I__2443 (
            .O(N__10814),
            .I(N__10785));
    LocalMux I__2442 (
            .O(N__10811),
            .I(N__10785));
    InMux I__2441 (
            .O(N__10810),
            .I(N__10782));
    Span4Mux_h I__2440 (
            .O(N__10805),
            .I(N__10779));
    LocalMux I__2439 (
            .O(N__10802),
            .I(N__10772));
    Span4Mux_v I__2438 (
            .O(N__10799),
            .I(N__10772));
    Span4Mux_v I__2437 (
            .O(N__10796),
            .I(N__10772));
    LocalMux I__2436 (
            .O(N__10793),
            .I(N__10765));
    Span4Mux_h I__2435 (
            .O(N__10790),
            .I(N__10765));
    Span4Mux_h I__2434 (
            .O(N__10785),
            .I(N__10765));
    LocalMux I__2433 (
            .O(N__10782),
            .I(un1_visiblex_24));
    Odrv4 I__2432 (
            .O(N__10779),
            .I(un1_visiblex_24));
    Odrv4 I__2431 (
            .O(N__10772),
            .I(un1_visiblex_24));
    Odrv4 I__2430 (
            .O(N__10765),
            .I(un1_visiblex_24));
    InMux I__2429 (
            .O(N__10756),
            .I(N__10753));
    LocalMux I__2428 (
            .O(N__10753),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_i));
    InMux I__2427 (
            .O(N__10750),
            .I(N__10747));
    LocalMux I__2426 (
            .O(N__10747),
            .I(g1_0_1));
    CascadeMux I__2425 (
            .O(N__10744),
            .I(N_17_cascade_));
    InMux I__2424 (
            .O(N__10741),
            .I(N__10738));
    LocalMux I__2423 (
            .O(N__10738),
            .I(G_25_i_a8_1));
    CascadeMux I__2422 (
            .O(N__10735),
            .I(g1_3_cascade_));
    CascadeMux I__2421 (
            .O(N__10732),
            .I(N_1302_0_0_0_cascade_));
    CascadeMux I__2420 (
            .O(N__10729),
            .I(N__10719));
    InMux I__2419 (
            .O(N__10728),
            .I(N__10716));
    InMux I__2418 (
            .O(N__10727),
            .I(N__10713));
    InMux I__2417 (
            .O(N__10726),
            .I(N__10710));
    InMux I__2416 (
            .O(N__10725),
            .I(N__10705));
    InMux I__2415 (
            .O(N__10724),
            .I(N__10705));
    InMux I__2414 (
            .O(N__10723),
            .I(N__10700));
    InMux I__2413 (
            .O(N__10722),
            .I(N__10700));
    InMux I__2412 (
            .O(N__10719),
            .I(N__10697));
    LocalMux I__2411 (
            .O(N__10716),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    LocalMux I__2410 (
            .O(N__10713),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    LocalMux I__2409 (
            .O(N__10710),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    LocalMux I__2408 (
            .O(N__10705),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    LocalMux I__2407 (
            .O(N__10700),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    LocalMux I__2406 (
            .O(N__10697),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9));
    InMux I__2405 (
            .O(N__10684),
            .I(N__10678));
    InMux I__2404 (
            .O(N__10683),
            .I(N__10670));
    InMux I__2403 (
            .O(N__10682),
            .I(N__10670));
    InMux I__2402 (
            .O(N__10681),
            .I(N__10667));
    LocalMux I__2401 (
            .O(N__10678),
            .I(N__10664));
    InMux I__2400 (
            .O(N__10677),
            .I(N__10659));
    InMux I__2399 (
            .O(N__10676),
            .I(N__10659));
    InMux I__2398 (
            .O(N__10675),
            .I(N__10656));
    LocalMux I__2397 (
            .O(N__10670),
            .I(N__10651));
    LocalMux I__2396 (
            .O(N__10667),
            .I(N__10651));
    Span4Mux_s3_h I__2395 (
            .O(N__10664),
            .I(N__10645));
    LocalMux I__2394 (
            .O(N__10659),
            .I(N__10640));
    LocalMux I__2393 (
            .O(N__10656),
            .I(N__10640));
    Span4Mux_v I__2392 (
            .O(N__10651),
            .I(N__10637));
    CascadeMux I__2391 (
            .O(N__10650),
            .I(N__10631));
    InMux I__2390 (
            .O(N__10649),
            .I(N__10628));
    InMux I__2389 (
            .O(N__10648),
            .I(N__10625));
    Span4Mux_h I__2388 (
            .O(N__10645),
            .I(N__10622));
    Span4Mux_v I__2387 (
            .O(N__10640),
            .I(N__10617));
    Span4Mux_h I__2386 (
            .O(N__10637),
            .I(N__10617));
    InMux I__2385 (
            .O(N__10636),
            .I(N__10610));
    InMux I__2384 (
            .O(N__10635),
            .I(N__10610));
    InMux I__2383 (
            .O(N__10634),
            .I(N__10610));
    InMux I__2382 (
            .O(N__10631),
            .I(N__10607));
    LocalMux I__2381 (
            .O(N__10628),
            .I(beamXZ0Z_0));
    LocalMux I__2380 (
            .O(N__10625),
            .I(beamXZ0Z_0));
    Odrv4 I__2379 (
            .O(N__10622),
            .I(beamXZ0Z_0));
    Odrv4 I__2378 (
            .O(N__10617),
            .I(beamXZ0Z_0));
    LocalMux I__2377 (
            .O(N__10610),
            .I(beamXZ0Z_0));
    LocalMux I__2376 (
            .O(N__10607),
            .I(beamXZ0Z_0));
    CascadeMux I__2375 (
            .O(N__10594),
            .I(N_159_0_0_cascade_));
    InMux I__2374 (
            .O(N__10591),
            .I(N__10588));
    LocalMux I__2373 (
            .O(N__10588),
            .I(N_156_0));
    InMux I__2372 (
            .O(N__10585),
            .I(N__10582));
    LocalMux I__2371 (
            .O(N__10582),
            .I(font_un314_pixel_0));
    CascadeMux I__2370 (
            .O(N__10579),
            .I(N__10568));
    CascadeMux I__2369 (
            .O(N__10578),
            .I(N__10565));
    InMux I__2368 (
            .O(N__10577),
            .I(N__10558));
    InMux I__2367 (
            .O(N__10576),
            .I(N__10558));
    InMux I__2366 (
            .O(N__10575),
            .I(N__10551));
    InMux I__2365 (
            .O(N__10574),
            .I(N__10551));
    InMux I__2364 (
            .O(N__10573),
            .I(N__10551));
    InMux I__2363 (
            .O(N__10572),
            .I(N__10540));
    InMux I__2362 (
            .O(N__10571),
            .I(N__10537));
    InMux I__2361 (
            .O(N__10568),
            .I(N__10534));
    InMux I__2360 (
            .O(N__10565),
            .I(N__10527));
    InMux I__2359 (
            .O(N__10564),
            .I(N__10527));
    InMux I__2358 (
            .O(N__10563),
            .I(N__10527));
    LocalMux I__2357 (
            .O(N__10558),
            .I(N__10524));
    LocalMux I__2356 (
            .O(N__10551),
            .I(N__10521));
    InMux I__2355 (
            .O(N__10550),
            .I(N__10516));
    InMux I__2354 (
            .O(N__10549),
            .I(N__10516));
    CascadeMux I__2353 (
            .O(N__10548),
            .I(N__10513));
    InMux I__2352 (
            .O(N__10547),
            .I(N__10506));
    InMux I__2351 (
            .O(N__10546),
            .I(N__10506));
    InMux I__2350 (
            .O(N__10545),
            .I(N__10506));
    InMux I__2349 (
            .O(N__10544),
            .I(N__10501));
    InMux I__2348 (
            .O(N__10543),
            .I(N__10501));
    LocalMux I__2347 (
            .O(N__10540),
            .I(N__10498));
    LocalMux I__2346 (
            .O(N__10537),
            .I(N__10493));
    LocalMux I__2345 (
            .O(N__10534),
            .I(N__10493));
    LocalMux I__2344 (
            .O(N__10527),
            .I(N__10489));
    Span4Mux_s3_h I__2343 (
            .O(N__10524),
            .I(N__10482));
    Span4Mux_v I__2342 (
            .O(N__10521),
            .I(N__10482));
    LocalMux I__2341 (
            .O(N__10516),
            .I(N__10482));
    InMux I__2340 (
            .O(N__10513),
            .I(N__10479));
    LocalMux I__2339 (
            .O(N__10506),
            .I(N__10474));
    LocalMux I__2338 (
            .O(N__10501),
            .I(N__10474));
    Span4Mux_v I__2337 (
            .O(N__10498),
            .I(N__10469));
    Span4Mux_v I__2336 (
            .O(N__10493),
            .I(N__10469));
    InMux I__2335 (
            .O(N__10492),
            .I(N__10466));
    Span4Mux_h I__2334 (
            .O(N__10489),
            .I(N__10461));
    Span4Mux_h I__2333 (
            .O(N__10482),
            .I(N__10461));
    LocalMux I__2332 (
            .O(N__10479),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum));
    Odrv12 I__2331 (
            .O(N__10474),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum));
    Odrv4 I__2330 (
            .O(N__10469),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum));
    LocalMux I__2329 (
            .O(N__10466),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum));
    Odrv4 I__2328 (
            .O(N__10461),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum));
    CascadeMux I__2327 (
            .O(N__10450),
            .I(N__10439));
    CascadeMux I__2326 (
            .O(N__10449),
            .I(N__10435));
    CascadeMux I__2325 (
            .O(N__10448),
            .I(N__10432));
    CascadeMux I__2324 (
            .O(N__10447),
            .I(N__10426));
    CascadeMux I__2323 (
            .O(N__10446),
            .I(N__10423));
    InMux I__2322 (
            .O(N__10445),
            .I(N__10419));
    InMux I__2321 (
            .O(N__10444),
            .I(N__10412));
    InMux I__2320 (
            .O(N__10443),
            .I(N__10412));
    InMux I__2319 (
            .O(N__10442),
            .I(N__10412));
    InMux I__2318 (
            .O(N__10439),
            .I(N__10407));
    InMux I__2317 (
            .O(N__10438),
            .I(N__10407));
    InMux I__2316 (
            .O(N__10435),
            .I(N__10400));
    InMux I__2315 (
            .O(N__10432),
            .I(N__10400));
    InMux I__2314 (
            .O(N__10431),
            .I(N__10400));
    InMux I__2313 (
            .O(N__10430),
            .I(N__10395));
    InMux I__2312 (
            .O(N__10429),
            .I(N__10395));
    InMux I__2311 (
            .O(N__10426),
            .I(N__10388));
    InMux I__2310 (
            .O(N__10423),
            .I(N__10388));
    InMux I__2309 (
            .O(N__10422),
            .I(N__10388));
    LocalMux I__2308 (
            .O(N__10419),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    LocalMux I__2307 (
            .O(N__10412),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    LocalMux I__2306 (
            .O(N__10407),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    LocalMux I__2305 (
            .O(N__10400),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    LocalMux I__2304 (
            .O(N__10395),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    LocalMux I__2303 (
            .O(N__10388),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1));
    InMux I__2302 (
            .O(N__10375),
            .I(N__10372));
    LocalMux I__2301 (
            .O(N__10372),
            .I(g1_3_0_0));
    CascadeMux I__2300 (
            .O(N__10369),
            .I(N__10364));
    InMux I__2299 (
            .O(N__10368),
            .I(N__10360));
    InMux I__2298 (
            .O(N__10367),
            .I(N__10347));
    InMux I__2297 (
            .O(N__10364),
            .I(N__10342));
    InMux I__2296 (
            .O(N__10363),
            .I(N__10339));
    LocalMux I__2295 (
            .O(N__10360),
            .I(N__10336));
    InMux I__2294 (
            .O(N__10359),
            .I(N__10333));
    InMux I__2293 (
            .O(N__10358),
            .I(N__10330));
    InMux I__2292 (
            .O(N__10357),
            .I(N__10327));
    InMux I__2291 (
            .O(N__10356),
            .I(N__10324));
    CascadeMux I__2290 (
            .O(N__10355),
            .I(N__10321));
    InMux I__2289 (
            .O(N__10354),
            .I(N__10316));
    InMux I__2288 (
            .O(N__10353),
            .I(N__10311));
    InMux I__2287 (
            .O(N__10352),
            .I(N__10311));
    InMux I__2286 (
            .O(N__10351),
            .I(N__10306));
    InMux I__2285 (
            .O(N__10350),
            .I(N__10306));
    LocalMux I__2284 (
            .O(N__10347),
            .I(N__10302));
    CascadeMux I__2283 (
            .O(N__10346),
            .I(N__10299));
    CascadeMux I__2282 (
            .O(N__10345),
            .I(N__10296));
    LocalMux I__2281 (
            .O(N__10342),
            .I(N__10293));
    LocalMux I__2280 (
            .O(N__10339),
            .I(N__10280));
    Span4Mux_v I__2279 (
            .O(N__10336),
            .I(N__10280));
    LocalMux I__2278 (
            .O(N__10333),
            .I(N__10280));
    LocalMux I__2277 (
            .O(N__10330),
            .I(N__10280));
    LocalMux I__2276 (
            .O(N__10327),
            .I(N__10280));
    LocalMux I__2275 (
            .O(N__10324),
            .I(N__10280));
    InMux I__2274 (
            .O(N__10321),
            .I(N__10277));
    InMux I__2273 (
            .O(N__10320),
            .I(N__10272));
    InMux I__2272 (
            .O(N__10319),
            .I(N__10272));
    LocalMux I__2271 (
            .O(N__10316),
            .I(N__10265));
    LocalMux I__2270 (
            .O(N__10311),
            .I(N__10265));
    LocalMux I__2269 (
            .O(N__10306),
            .I(N__10265));
    InMux I__2268 (
            .O(N__10305),
            .I(N__10262));
    Span4Mux_h I__2267 (
            .O(N__10302),
            .I(N__10258));
    InMux I__2266 (
            .O(N__10299),
            .I(N__10255));
    InMux I__2265 (
            .O(N__10296),
            .I(N__10252));
    Span4Mux_h I__2264 (
            .O(N__10293),
            .I(N__10247));
    Span4Mux_v I__2263 (
            .O(N__10280),
            .I(N__10247));
    LocalMux I__2262 (
            .O(N__10277),
            .I(N__10238));
    LocalMux I__2261 (
            .O(N__10272),
            .I(N__10238));
    Span4Mux_v I__2260 (
            .O(N__10265),
            .I(N__10238));
    LocalMux I__2259 (
            .O(N__10262),
            .I(N__10238));
    InMux I__2258 (
            .O(N__10261),
            .I(N__10235));
    Span4Mux_h I__2257 (
            .O(N__10258),
            .I(N__10232));
    LocalMux I__2256 (
            .O(N__10255),
            .I(un28lto1));
    LocalMux I__2255 (
            .O(N__10252),
            .I(un28lto1));
    Odrv4 I__2254 (
            .O(N__10247),
            .I(un28lto1));
    Odrv4 I__2253 (
            .O(N__10238),
            .I(un28lto1));
    LocalMux I__2252 (
            .O(N__10235),
            .I(un28lto1));
    Odrv4 I__2251 (
            .O(N__10232),
            .I(un28lto1));
    CascadeMux I__2250 (
            .O(N__10219),
            .I(N__10206));
    InMux I__2249 (
            .O(N__10218),
            .I(N__10203));
    InMux I__2248 (
            .O(N__10217),
            .I(N__10200));
    InMux I__2247 (
            .O(N__10216),
            .I(N__10193));
    InMux I__2246 (
            .O(N__10215),
            .I(N__10193));
    InMux I__2245 (
            .O(N__10214),
            .I(N__10193));
    InMux I__2244 (
            .O(N__10213),
            .I(N__10187));
    InMux I__2243 (
            .O(N__10212),
            .I(N__10184));
    InMux I__2242 (
            .O(N__10211),
            .I(N__10181));
    InMux I__2241 (
            .O(N__10210),
            .I(N__10176));
    InMux I__2240 (
            .O(N__10209),
            .I(N__10176));
    InMux I__2239 (
            .O(N__10206),
            .I(N__10172));
    LocalMux I__2238 (
            .O(N__10203),
            .I(N__10167));
    LocalMux I__2237 (
            .O(N__10200),
            .I(N__10167));
    LocalMux I__2236 (
            .O(N__10193),
            .I(N__10164));
    InMux I__2235 (
            .O(N__10192),
            .I(N__10161));
    InMux I__2234 (
            .O(N__10191),
            .I(N__10158));
    CascadeMux I__2233 (
            .O(N__10190),
            .I(N__10155));
    LocalMux I__2232 (
            .O(N__10187),
            .I(N__10152));
    LocalMux I__2231 (
            .O(N__10184),
            .I(N__10145));
    LocalMux I__2230 (
            .O(N__10181),
            .I(N__10145));
    LocalMux I__2229 (
            .O(N__10176),
            .I(N__10145));
    CascadeMux I__2228 (
            .O(N__10175),
            .I(N__10142));
    LocalMux I__2227 (
            .O(N__10172),
            .I(N__10139));
    Span4Mux_v I__2226 (
            .O(N__10167),
            .I(N__10134));
    Span4Mux_v I__2225 (
            .O(N__10164),
            .I(N__10134));
    LocalMux I__2224 (
            .O(N__10161),
            .I(N__10130));
    LocalMux I__2223 (
            .O(N__10158),
            .I(N__10127));
    InMux I__2222 (
            .O(N__10155),
            .I(N__10124));
    Span4Mux_v I__2221 (
            .O(N__10152),
            .I(N__10119));
    Span4Mux_v I__2220 (
            .O(N__10145),
            .I(N__10119));
    InMux I__2219 (
            .O(N__10142),
            .I(N__10116));
    Span4Mux_h I__2218 (
            .O(N__10139),
            .I(N__10111));
    Span4Mux_h I__2217 (
            .O(N__10134),
            .I(N__10111));
    InMux I__2216 (
            .O(N__10133),
            .I(N__10108));
    Span4Mux_v I__2215 (
            .O(N__10130),
            .I(N__10103));
    Span4Mux_h I__2214 (
            .O(N__10127),
            .I(N__10103));
    LocalMux I__2213 (
            .O(N__10124),
            .I(N__10100));
    Span4Mux_h I__2212 (
            .O(N__10119),
            .I(N__10097));
    LocalMux I__2211 (
            .O(N__10116),
            .I(N__10092));
    Span4Mux_v I__2210 (
            .O(N__10111),
            .I(N__10092));
    LocalMux I__2209 (
            .O(N__10108),
            .I(N__10087));
    Span4Mux_v I__2208 (
            .O(N__10103),
            .I(N__10087));
    Odrv4 I__2207 (
            .O(N__10100),
            .I(beamYZ0Z_0));
    Odrv4 I__2206 (
            .O(N__10097),
            .I(beamYZ0Z_0));
    Odrv4 I__2205 (
            .O(N__10092),
            .I(beamYZ0Z_0));
    Odrv4 I__2204 (
            .O(N__10087),
            .I(beamYZ0Z_0));
    InMux I__2203 (
            .O(N__10078),
            .I(N__10065));
    InMux I__2202 (
            .O(N__10077),
            .I(N__10065));
    InMux I__2201 (
            .O(N__10076),
            .I(N__10060));
    InMux I__2200 (
            .O(N__10075),
            .I(N__10057));
    InMux I__2199 (
            .O(N__10074),
            .I(N__10054));
    InMux I__2198 (
            .O(N__10073),
            .I(N__10047));
    InMux I__2197 (
            .O(N__10072),
            .I(N__10047));
    InMux I__2196 (
            .O(N__10071),
            .I(N__10047));
    InMux I__2195 (
            .O(N__10070),
            .I(N__10043));
    LocalMux I__2194 (
            .O(N__10065),
            .I(N__10040));
    InMux I__2193 (
            .O(N__10064),
            .I(N__10035));
    InMux I__2192 (
            .O(N__10063),
            .I(N__10035));
    LocalMux I__2191 (
            .O(N__10060),
            .I(N__10027));
    LocalMux I__2190 (
            .O(N__10057),
            .I(N__10027));
    LocalMux I__2189 (
            .O(N__10054),
            .I(N__10022));
    LocalMux I__2188 (
            .O(N__10047),
            .I(N__10022));
    InMux I__2187 (
            .O(N__10046),
            .I(N__10019));
    LocalMux I__2186 (
            .O(N__10043),
            .I(N__10012));
    Span4Mux_v I__2185 (
            .O(N__10040),
            .I(N__10012));
    LocalMux I__2184 (
            .O(N__10035),
            .I(N__10012));
    InMux I__2183 (
            .O(N__10034),
            .I(N__10009));
    InMux I__2182 (
            .O(N__10033),
            .I(N__10004));
    InMux I__2181 (
            .O(N__10032),
            .I(N__10004));
    Span4Mux_h I__2180 (
            .O(N__10027),
            .I(N__10001));
    Span4Mux_h I__2179 (
            .O(N__10022),
            .I(N__9998));
    LocalMux I__2178 (
            .O(N__10019),
            .I(N__9995));
    Span4Mux_h I__2177 (
            .O(N__10012),
            .I(N__9992));
    LocalMux I__2176 (
            .O(N__10009),
            .I(font_un42_pixel_23));
    LocalMux I__2175 (
            .O(N__10004),
            .I(font_un42_pixel_23));
    Odrv4 I__2174 (
            .O(N__10001),
            .I(font_un42_pixel_23));
    Odrv4 I__2173 (
            .O(N__9998),
            .I(font_un42_pixel_23));
    Odrv12 I__2172 (
            .O(N__9995),
            .I(font_un42_pixel_23));
    Odrv4 I__2171 (
            .O(N__9992),
            .I(font_un42_pixel_23));
    InMux I__2170 (
            .O(N__9979),
            .I(N__9976));
    LocalMux I__2169 (
            .O(N__9976),
            .I(N_1303_0_0));
    CascadeMux I__2168 (
            .O(N__9973),
            .I(un28lto4_1_cascade_));
    InMux I__2167 (
            .O(N__9970),
            .I(N__9967));
    LocalMux I__2166 (
            .O(N__9967),
            .I(Pixel_1_esr_RNOZ0Z_62));
    CascadeMux I__2165 (
            .O(N__9964),
            .I(un28lt10_cascade_));
    InMux I__2164 (
            .O(N__9961),
            .I(N__9952));
    InMux I__2163 (
            .O(N__9960),
            .I(N__9952));
    InMux I__2162 (
            .O(N__9959),
            .I(N__9952));
    LocalMux I__2161 (
            .O(N__9952),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0));
    InMux I__2160 (
            .O(N__9949),
            .I(N__9946));
    LocalMux I__2159 (
            .O(N__9946),
            .I(un28_0_1));
    InMux I__2158 (
            .O(N__9943),
            .I(N__9937));
    InMux I__2157 (
            .O(N__9942),
            .I(N__9937));
    LocalMux I__2156 (
            .O(N__9937),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0));
    InMux I__2155 (
            .O(N__9934),
            .I(N__9928));
    InMux I__2154 (
            .O(N__9933),
            .I(N__9928));
    LocalMux I__2153 (
            .O(N__9928),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0));
    CascadeMux I__2152 (
            .O(N__9925),
            .I(N__9918));
    CascadeMux I__2151 (
            .O(N__9924),
            .I(N__9915));
    InMux I__2150 (
            .O(N__9923),
            .I(N__9912));
    InMux I__2149 (
            .O(N__9922),
            .I(N__9905));
    InMux I__2148 (
            .O(N__9921),
            .I(N__9905));
    InMux I__2147 (
            .O(N__9918),
            .I(N__9905));
    InMux I__2146 (
            .O(N__9915),
            .I(N__9902));
    LocalMux I__2145 (
            .O(N__9912),
            .I(beamY_i_2));
    LocalMux I__2144 (
            .O(N__9905),
            .I(beamY_i_2));
    LocalMux I__2143 (
            .O(N__9902),
            .I(beamY_i_2));
    InMux I__2142 (
            .O(N__9895),
            .I(N__9892));
    LocalMux I__2141 (
            .O(N__9892),
            .I(un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5));
    SRMux I__2140 (
            .O(N__9889),
            .I(N__9885));
    InMux I__2139 (
            .O(N__9888),
            .I(N__9882));
    LocalMux I__2138 (
            .O(N__9885),
            .I(N__9879));
    LocalMux I__2137 (
            .O(N__9882),
            .I(N__9876));
    Span4Mux_h I__2136 (
            .O(N__9879),
            .I(N__9872));
    Span4Mux_h I__2135 (
            .O(N__9876),
            .I(N__9869));
    InMux I__2134 (
            .O(N__9875),
            .I(N__9866));
    Odrv4 I__2133 (
            .O(N__9872),
            .I(beamY_RNIJ0DBZ0Z_9));
    Odrv4 I__2132 (
            .O(N__9869),
            .I(beamY_RNIJ0DBZ0Z_9));
    LocalMux I__2131 (
            .O(N__9866),
            .I(beamY_RNIJ0DBZ0Z_9));
    IoInMux I__2130 (
            .O(N__9859),
            .I(N__9856));
    LocalMux I__2129 (
            .O(N__9856),
            .I(N__9852));
    IoInMux I__2128 (
            .O(N__9855),
            .I(N__9849));
    Span4Mux_s0_v I__2127 (
            .O(N__9852),
            .I(N__9846));
    LocalMux I__2126 (
            .O(N__9849),
            .I(N__9843));
    Span4Mux_v I__2125 (
            .O(N__9846),
            .I(N__9840));
    IoSpan4Mux I__2124 (
            .O(N__9843),
            .I(N__9837));
    Span4Mux_v I__2123 (
            .O(N__9840),
            .I(N__9834));
    Span4Mux_s3_v I__2122 (
            .O(N__9837),
            .I(N__9831));
    Odrv4 I__2121 (
            .O(N__9834),
            .I(VSync_c));
    Odrv4 I__2120 (
            .O(N__9831),
            .I(VSync_c));
    ClkMux I__2119 (
            .O(N__9826),
            .I(N__9781));
    ClkMux I__2118 (
            .O(N__9825),
            .I(N__9781));
    ClkMux I__2117 (
            .O(N__9824),
            .I(N__9781));
    ClkMux I__2116 (
            .O(N__9823),
            .I(N__9781));
    ClkMux I__2115 (
            .O(N__9822),
            .I(N__9781));
    ClkMux I__2114 (
            .O(N__9821),
            .I(N__9781));
    ClkMux I__2113 (
            .O(N__9820),
            .I(N__9781));
    ClkMux I__2112 (
            .O(N__9819),
            .I(N__9781));
    ClkMux I__2111 (
            .O(N__9818),
            .I(N__9781));
    ClkMux I__2110 (
            .O(N__9817),
            .I(N__9781));
    ClkMux I__2109 (
            .O(N__9816),
            .I(N__9781));
    ClkMux I__2108 (
            .O(N__9815),
            .I(N__9781));
    ClkMux I__2107 (
            .O(N__9814),
            .I(N__9781));
    ClkMux I__2106 (
            .O(N__9813),
            .I(N__9781));
    ClkMux I__2105 (
            .O(N__9812),
            .I(N__9781));
    GlobalMux I__2104 (
            .O(N__9781),
            .I(N__9778));
    gio2CtrlBuf I__2103 (
            .O(N__9778),
            .I(PixelClock_g));
    CascadeMux I__2102 (
            .O(N__9775),
            .I(g1_1_cascade_));
    InMux I__2101 (
            .O(N__9772),
            .I(N__9769));
    LocalMux I__2100 (
            .O(N__9769),
            .I(Pixel_1_esr_RNOZ0Z_39));
    CascadeMux I__2099 (
            .O(N__9766),
            .I(N_1304_0_cascade_));
    CascadeMux I__2098 (
            .O(N__9763),
            .I(N__9755));
    InMux I__2097 (
            .O(N__9762),
            .I(N__9749));
    InMux I__2096 (
            .O(N__9761),
            .I(N__9744));
    InMux I__2095 (
            .O(N__9760),
            .I(N__9744));
    InMux I__2094 (
            .O(N__9759),
            .I(N__9741));
    InMux I__2093 (
            .O(N__9758),
            .I(N__9738));
    InMux I__2092 (
            .O(N__9755),
            .I(N__9733));
    InMux I__2091 (
            .O(N__9754),
            .I(N__9733));
    InMux I__2090 (
            .O(N__9753),
            .I(N__9730));
    InMux I__2089 (
            .O(N__9752),
            .I(N__9727));
    LocalMux I__2088 (
            .O(N__9749),
            .I(N__9720));
    LocalMux I__2087 (
            .O(N__9744),
            .I(N__9720));
    LocalMux I__2086 (
            .O(N__9741),
            .I(N__9715));
    LocalMux I__2085 (
            .O(N__9738),
            .I(N__9712));
    LocalMux I__2084 (
            .O(N__9733),
            .I(N__9709));
    LocalMux I__2083 (
            .O(N__9730),
            .I(N__9704));
    LocalMux I__2082 (
            .O(N__9727),
            .I(N__9704));
    InMux I__2081 (
            .O(N__9726),
            .I(N__9701));
    InMux I__2080 (
            .O(N__9725),
            .I(N__9698));
    Span4Mux_v I__2079 (
            .O(N__9720),
            .I(N__9695));
    InMux I__2078 (
            .O(N__9719),
            .I(N__9690));
    InMux I__2077 (
            .O(N__9718),
            .I(N__9690));
    Span4Mux_h I__2076 (
            .O(N__9715),
            .I(N__9685));
    Span4Mux_h I__2075 (
            .O(N__9712),
            .I(N__9685));
    Span4Mux_h I__2074 (
            .O(N__9709),
            .I(N__9680));
    Span4Mux_h I__2073 (
            .O(N__9704),
            .I(N__9680));
    LocalMux I__2072 (
            .O(N__9701),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    LocalMux I__2071 (
            .O(N__9698),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__2070 (
            .O(N__9695),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    LocalMux I__2069 (
            .O(N__9690),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__2068 (
            .O(N__9685),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__2067 (
            .O(N__9680),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    InMux I__2066 (
            .O(N__9667),
            .I(N__9664));
    LocalMux I__2065 (
            .O(N__9664),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__2064 (
            .O(N__9661),
            .I(N__9658));
    LocalMux I__2063 (
            .O(N__9658),
            .I(N__9652));
    InMux I__2062 (
            .O(N__9657),
            .I(N__9649));
    InMux I__2061 (
            .O(N__9656),
            .I(N__9642));
    InMux I__2060 (
            .O(N__9655),
            .I(N__9642));
    Span4Mux_h I__2059 (
            .O(N__9652),
            .I(N__9633));
    LocalMux I__2058 (
            .O(N__9649),
            .I(N__9633));
    InMux I__2057 (
            .O(N__9648),
            .I(N__9630));
    InMux I__2056 (
            .O(N__9647),
            .I(N__9627));
    LocalMux I__2055 (
            .O(N__9642),
            .I(N__9624));
    InMux I__2054 (
            .O(N__9641),
            .I(N__9619));
    InMux I__2053 (
            .O(N__9640),
            .I(N__9619));
    InMux I__2052 (
            .O(N__9639),
            .I(N__9616));
    InMux I__2051 (
            .O(N__9638),
            .I(N__9613));
    Span4Mux_v I__2050 (
            .O(N__9633),
            .I(N__9610));
    LocalMux I__2049 (
            .O(N__9630),
            .I(N__9605));
    LocalMux I__2048 (
            .O(N__9627),
            .I(N__9605));
    Span4Mux_h I__2047 (
            .O(N__9624),
            .I(N__9602));
    LocalMux I__2046 (
            .O(N__9619),
            .I(N__9599));
    LocalMux I__2045 (
            .O(N__9616),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    LocalMux I__2044 (
            .O(N__9613),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2043 (
            .O(N__9610),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2042 (
            .O(N__9605),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2041 (
            .O(N__9602),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__2040 (
            .O(N__9599),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    CascadeMux I__2039 (
            .O(N__9586),
            .I(N__9581));
    InMux I__2038 (
            .O(N__9585),
            .I(N__9576));
    InMux I__2037 (
            .O(N__9584),
            .I(N__9569));
    InMux I__2036 (
            .O(N__9581),
            .I(N__9569));
    InMux I__2035 (
            .O(N__9580),
            .I(N__9569));
    CascadeMux I__2034 (
            .O(N__9579),
            .I(N__9566));
    LocalMux I__2033 (
            .O(N__9576),
            .I(N__9556));
    LocalMux I__2032 (
            .O(N__9569),
            .I(N__9556));
    InMux I__2031 (
            .O(N__9566),
            .I(N__9553));
    InMux I__2030 (
            .O(N__9565),
            .I(N__9550));
    CascadeMux I__2029 (
            .O(N__9564),
            .I(N__9547));
    CascadeMux I__2028 (
            .O(N__9563),
            .I(N__9541));
    InMux I__2027 (
            .O(N__9562),
            .I(N__9534));
    InMux I__2026 (
            .O(N__9561),
            .I(N__9534));
    Span4Mux_v I__2025 (
            .O(N__9556),
            .I(N__9531));
    LocalMux I__2024 (
            .O(N__9553),
            .I(N__9528));
    LocalMux I__2023 (
            .O(N__9550),
            .I(N__9525));
    InMux I__2022 (
            .O(N__9547),
            .I(N__9522));
    InMux I__2021 (
            .O(N__9546),
            .I(N__9513));
    InMux I__2020 (
            .O(N__9545),
            .I(N__9513));
    InMux I__2019 (
            .O(N__9544),
            .I(N__9513));
    InMux I__2018 (
            .O(N__9541),
            .I(N__9513));
    InMux I__2017 (
            .O(N__9540),
            .I(N__9508));
    InMux I__2016 (
            .O(N__9539),
            .I(N__9508));
    LocalMux I__2015 (
            .O(N__9534),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    Odrv4 I__2014 (
            .O(N__9531),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    Odrv12 I__2013 (
            .O(N__9528),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    Odrv4 I__2012 (
            .O(N__9525),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    LocalMux I__2011 (
            .O(N__9522),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    LocalMux I__2010 (
            .O(N__9513),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    LocalMux I__2009 (
            .O(N__9508),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6));
    InMux I__2008 (
            .O(N__9493),
            .I(N__9490));
    LocalMux I__2007 (
            .O(N__9490),
            .I(N__9487));
    Odrv12 I__2006 (
            .O(N__9487),
            .I(g0_i_o4_2));
    InMux I__2005 (
            .O(N__9484),
            .I(N__9481));
    LocalMux I__2004 (
            .O(N__9481),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__2003 (
            .O(N__9478),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__2002 (
            .O(N__9475),
            .I(N__9472));
    InMux I__2001 (
            .O(N__9472),
            .I(N__9469));
    LocalMux I__2000 (
            .O(N__9469),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5));
    InMux I__1999 (
            .O(N__9466),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__1998 (
            .O(N__9463),
            .I(N__9460));
    LocalMux I__1997 (
            .O(N__9460),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399));
    InMux I__1996 (
            .O(N__9457),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1995 (
            .O(N__9454),
            .I(N__9451));
    InMux I__1994 (
            .O(N__9451),
            .I(N__9448));
    LocalMux I__1993 (
            .O(N__9448),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9));
    CascadeMux I__1992 (
            .O(N__9445),
            .I(N__9440));
    CascadeMux I__1991 (
            .O(N__9444),
            .I(N__9436));
    InMux I__1990 (
            .O(N__9443),
            .I(N__9432));
    InMux I__1989 (
            .O(N__9440),
            .I(N__9423));
    InMux I__1988 (
            .O(N__9439),
            .I(N__9423));
    InMux I__1987 (
            .O(N__9436),
            .I(N__9423));
    InMux I__1986 (
            .O(N__9435),
            .I(N__9423));
    LocalMux I__1985 (
            .O(N__9432),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0));
    LocalMux I__1984 (
            .O(N__9423),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0));
    InMux I__1983 (
            .O(N__9418),
            .I(N__9415));
    LocalMux I__1982 (
            .O(N__9415),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__1981 (
            .O(N__9412),
            .I(N__9409));
    LocalMux I__1980 (
            .O(N__9409),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__1979 (
            .O(N__9406),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6));
    CascadeMux I__1978 (
            .O(N__9403),
            .I(g0_1_0_cascade_));
    InMux I__1977 (
            .O(N__9400),
            .I(N__9397));
    LocalMux I__1976 (
            .O(N__9397),
            .I(g3_0_0));
    InMux I__1975 (
            .O(N__9394),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__1974 (
            .O(N__9391),
            .I(N__9387));
    InMux I__1973 (
            .O(N__9390),
            .I(N__9384));
    LocalMux I__1972 (
            .O(N__9387),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5));
    LocalMux I__1971 (
            .O(N__9384),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5));
    CascadeMux I__1970 (
            .O(N__9379),
            .I(N__9376));
    InMux I__1969 (
            .O(N__9376),
            .I(N__9373));
    LocalMux I__1968 (
            .O(N__9373),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43));
    InMux I__1967 (
            .O(N__9370),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__1966 (
            .O(N__9367),
            .I(N__9364));
    LocalMux I__1965 (
            .O(N__9364),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4));
    CascadeMux I__1964 (
            .O(N__9361),
            .I(N__9357));
    CascadeMux I__1963 (
            .O(N__9360),
            .I(N__9354));
    InMux I__1962 (
            .O(N__9357),
            .I(N__9349));
    InMux I__1961 (
            .O(N__9354),
            .I(N__9349));
    LocalMux I__1960 (
            .O(N__9349),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__1959 (
            .O(N__9346),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__1958 (
            .O(N__9343),
            .I(N__9340));
    LocalMux I__1957 (
            .O(N__9340),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__1956 (
            .O(N__9337),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__1955 (
            .O(N__9334),
            .I(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_));
    CascadeMux I__1954 (
            .O(N__9331),
            .I(N__9327));
    CascadeMux I__1953 (
            .O(N__9330),
            .I(N__9324));
    InMux I__1952 (
            .O(N__9327),
            .I(N__9319));
    InMux I__1951 (
            .O(N__9324),
            .I(N__9319));
    LocalMux I__1950 (
            .O(N__9319),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5));
    InMux I__1949 (
            .O(N__9316),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1948 (
            .O(N__9313),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_));
    InMux I__1947 (
            .O(N__9310),
            .I(N__9307));
    LocalMux I__1946 (
            .O(N__9307),
            .I(g1_0_1_1));
    CascadeMux I__1945 (
            .O(N__9304),
            .I(font_un19_pixel_0_0_0_23_cascade_));
    InMux I__1944 (
            .O(N__9301),
            .I(N__9298));
    LocalMux I__1943 (
            .O(N__9298),
            .I(g2_0));
    InMux I__1942 (
            .O(N__9295),
            .I(N__9292));
    LocalMux I__1941 (
            .O(N__9292),
            .I(g1_0_2));
    CascadeMux I__1940 (
            .O(N__9289),
            .I(font_un237_pixel_6_ns_1_0_0_cascade_));
    InMux I__1939 (
            .O(N__9286),
            .I(N__9283));
    LocalMux I__1938 (
            .O(N__9283),
            .I(g1_2_0));
    CascadeMux I__1937 (
            .O(N__9280),
            .I(N__9277));
    InMux I__1936 (
            .O(N__9277),
            .I(N__9274));
    LocalMux I__1935 (
            .O(N__9274),
            .I(font_un237_pixel_0_0));
    CascadeMux I__1934 (
            .O(N__9271),
            .I(g2_cascade_));
    InMux I__1933 (
            .O(N__9268),
            .I(N__9265));
    LocalMux I__1932 (
            .O(N__9265),
            .I(font_un83_pixel_0_0));
    InMux I__1931 (
            .O(N__9262),
            .I(N__9259));
    LocalMux I__1930 (
            .O(N__9259),
            .I(font_un19_pixel_23));
    CascadeMux I__1929 (
            .O(N__9256),
            .I(font_un19_pixel_23_cascade_));
    InMux I__1928 (
            .O(N__9253),
            .I(N__9250));
    LocalMux I__1927 (
            .O(N__9250),
            .I(N__9247));
    Odrv4 I__1926 (
            .O(N__9247),
            .I(font_un160_pixel_6_1));
    InMux I__1925 (
            .O(N__9244),
            .I(N__9241));
    LocalMux I__1924 (
            .O(N__9241),
            .I(N__9238));
    Span4Mux_h I__1923 (
            .O(N__9238),
            .I(N__9235));
    Odrv4 I__1922 (
            .O(N__9235),
            .I(g0_i_o4_3));
    InMux I__1921 (
            .O(N__9232),
            .I(N__9229));
    LocalMux I__1920 (
            .O(N__9229),
            .I(Pixel_9_u_ns_sn));
    CascadeMux I__1919 (
            .O(N__9226),
            .I(N_163_cascade_));
    IoInMux I__1918 (
            .O(N__9223),
            .I(N__9219));
    IoInMux I__1917 (
            .O(N__9222),
            .I(N__9216));
    LocalMux I__1916 (
            .O(N__9219),
            .I(N__9213));
    LocalMux I__1915 (
            .O(N__9216),
            .I(N__9210));
    Span4Mux_s3_v I__1914 (
            .O(N__9213),
            .I(N__9207));
    Span4Mux_s3_v I__1913 (
            .O(N__9210),
            .I(N__9204));
    Span4Mux_v I__1912 (
            .O(N__9207),
            .I(N__9201));
    Span4Mux_v I__1911 (
            .O(N__9204),
            .I(N__9198));
    Odrv4 I__1910 (
            .O(N__9201),
            .I(Pixel_c));
    Odrv4 I__1909 (
            .O(N__9198),
            .I(Pixel_c));
    CEMux I__1908 (
            .O(N__9193),
            .I(N__9190));
    LocalMux I__1907 (
            .O(N__9190),
            .I(Pixel_1_sqmuxa_i_0));
    InMux I__1906 (
            .O(N__9187),
            .I(N__9184));
    LocalMux I__1905 (
            .O(N__9184),
            .I(g1_0_0));
    InMux I__1904 (
            .O(N__9181),
            .I(N__9178));
    LocalMux I__1903 (
            .O(N__9178),
            .I(g0_0_4));
    InMux I__1902 (
            .O(N__9175),
            .I(N__9172));
    LocalMux I__1901 (
            .O(N__9172),
            .I(G_25_i_a8_2_0));
    CascadeMux I__1900 (
            .O(N__9169),
            .I(g0_0_5_cascade_));
    InMux I__1899 (
            .O(N__9166),
            .I(N__9163));
    LocalMux I__1898 (
            .O(N__9163),
            .I(G_25_i_3_0));
    InMux I__1897 (
            .O(N__9160),
            .I(N__9157));
    LocalMux I__1896 (
            .O(N__9157),
            .I(N_20));
    CascadeMux I__1895 (
            .O(N__9154),
            .I(G_25_i_2_0_cascade_));
    InMux I__1894 (
            .O(N__9151),
            .I(N__9148));
    LocalMux I__1893 (
            .O(N__9148),
            .I(G_25_i_0));
    InMux I__1892 (
            .O(N__9145),
            .I(N__9142));
    LocalMux I__1891 (
            .O(N__9142),
            .I(Pixel_9_u_ns_rn_0));
    CascadeMux I__1890 (
            .O(N__9139),
            .I(N__9136));
    InMux I__1889 (
            .O(N__9136),
            .I(N__9133));
    LocalMux I__1888 (
            .O(N__9133),
            .I(g2_1));
    InMux I__1887 (
            .O(N__9130),
            .I(N__9127));
    LocalMux I__1886 (
            .O(N__9127),
            .I(font_un19_pixel_if_generate_plus_mult1_un68_sum_i));
    InMux I__1885 (
            .O(N__9124),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__1884 (
            .O(N__9121),
            .I(N__9118));
    LocalMux I__1883 (
            .O(N__9118),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21));
    InMux I__1882 (
            .O(N__9115),
            .I(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__1881 (
            .O(N__9112),
            .I(N__9106));
    CascadeMux I__1880 (
            .O(N__9111),
            .I(N__9103));
    CascadeMux I__1879 (
            .O(N__9110),
            .I(N__9099));
    CascadeMux I__1878 (
            .O(N__9109),
            .I(N__9096));
    InMux I__1877 (
            .O(N__9106),
            .I(N__9091));
    InMux I__1876 (
            .O(N__9103),
            .I(N__9086));
    InMux I__1875 (
            .O(N__9102),
            .I(N__9086));
    InMux I__1874 (
            .O(N__9099),
            .I(N__9083));
    InMux I__1873 (
            .O(N__9096),
            .I(N__9080));
    InMux I__1872 (
            .O(N__9095),
            .I(N__9077));
    IoInMux I__1871 (
            .O(N__9094),
            .I(N__9072));
    LocalMux I__1870 (
            .O(N__9091),
            .I(N__9063));
    LocalMux I__1869 (
            .O(N__9086),
            .I(N__9063));
    LocalMux I__1868 (
            .O(N__9083),
            .I(N__9063));
    LocalMux I__1867 (
            .O(N__9080),
            .I(N__9063));
    LocalMux I__1866 (
            .O(N__9077),
            .I(N__9060));
    InMux I__1865 (
            .O(N__9076),
            .I(N__9057));
    InMux I__1864 (
            .O(N__9075),
            .I(N__9054));
    LocalMux I__1863 (
            .O(N__9072),
            .I(N__9049));
    Span4Mux_h I__1862 (
            .O(N__9063),
            .I(N__9046));
    Span4Mux_v I__1861 (
            .O(N__9060),
            .I(N__9039));
    LocalMux I__1860 (
            .O(N__9057),
            .I(N__9039));
    LocalMux I__1859 (
            .O(N__9054),
            .I(N__9039));
    InMux I__1858 (
            .O(N__9053),
            .I(N__9036));
    CascadeMux I__1857 (
            .O(N__9052),
            .I(N__9032));
    Span12Mux_s11_v I__1856 (
            .O(N__9049),
            .I(N__9029));
    Span4Mux_v I__1855 (
            .O(N__9046),
            .I(N__9022));
    Span4Mux_h I__1854 (
            .O(N__9039),
            .I(N__9022));
    LocalMux I__1853 (
            .O(N__9036),
            .I(N__9022));
    InMux I__1852 (
            .O(N__9035),
            .I(N__9019));
    InMux I__1851 (
            .O(N__9032),
            .I(N__9016));
    Odrv12 I__1850 (
            .O(N__9029),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1849 (
            .O(N__9022),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1848 (
            .O(N__9019),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1847 (
            .O(N__9016),
            .I(CONSTANT_ONE_NET));
    InMux I__1846 (
            .O(N__9007),
            .I(N__8997));
    InMux I__1845 (
            .O(N__9006),
            .I(N__8997));
    InMux I__1844 (
            .O(N__9005),
            .I(N__8997));
    InMux I__1843 (
            .O(N__9004),
            .I(N__8987));
    LocalMux I__1842 (
            .O(N__8997),
            .I(N__8984));
    InMux I__1841 (
            .O(N__8996),
            .I(N__8981));
    InMux I__1840 (
            .O(N__8995),
            .I(N__8976));
    InMux I__1839 (
            .O(N__8994),
            .I(N__8976));
    InMux I__1838 (
            .O(N__8993),
            .I(N__8973));
    InMux I__1837 (
            .O(N__8992),
            .I(N__8970));
    InMux I__1836 (
            .O(N__8991),
            .I(N__8966));
    InMux I__1835 (
            .O(N__8990),
            .I(N__8963));
    LocalMux I__1834 (
            .O(N__8987),
            .I(N__8954));
    Span4Mux_v I__1833 (
            .O(N__8984),
            .I(N__8954));
    LocalMux I__1832 (
            .O(N__8981),
            .I(N__8954));
    LocalMux I__1831 (
            .O(N__8976),
            .I(N__8954));
    LocalMux I__1830 (
            .O(N__8973),
            .I(N__8949));
    LocalMux I__1829 (
            .O(N__8970),
            .I(N__8949));
    InMux I__1828 (
            .O(N__8969),
            .I(N__8946));
    LocalMux I__1827 (
            .O(N__8966),
            .I(N__8942));
    LocalMux I__1826 (
            .O(N__8963),
            .I(N__8933));
    Span4Mux_v I__1825 (
            .O(N__8954),
            .I(N__8933));
    Span4Mux_v I__1824 (
            .O(N__8949),
            .I(N__8933));
    LocalMux I__1823 (
            .O(N__8946),
            .I(N__8933));
    InMux I__1822 (
            .O(N__8945),
            .I(N__8930));
    Odrv12 I__1821 (
            .O(N__8942),
            .I(beamYZ0Z_2));
    Odrv4 I__1820 (
            .O(N__8933),
            .I(beamYZ0Z_2));
    LocalMux I__1819 (
            .O(N__8930),
            .I(beamYZ0Z_2));
    InMux I__1818 (
            .O(N__8923),
            .I(N__8915));
    InMux I__1817 (
            .O(N__8922),
            .I(N__8915));
    InMux I__1816 (
            .O(N__8921),
            .I(N__8911));
    InMux I__1815 (
            .O(N__8920),
            .I(N__8908));
    LocalMux I__1814 (
            .O(N__8915),
            .I(N__8905));
    InMux I__1813 (
            .O(N__8914),
            .I(N__8902));
    LocalMux I__1812 (
            .O(N__8911),
            .I(N__8898));
    LocalMux I__1811 (
            .O(N__8908),
            .I(N__8895));
    Span4Mux_v I__1810 (
            .O(N__8905),
            .I(N__8890));
    LocalMux I__1809 (
            .O(N__8902),
            .I(N__8890));
    InMux I__1808 (
            .O(N__8901),
            .I(N__8883));
    Span4Mux_v I__1807 (
            .O(N__8898),
            .I(N__8880));
    Span4Mux_h I__1806 (
            .O(N__8895),
            .I(N__8875));
    Span4Mux_h I__1805 (
            .O(N__8890),
            .I(N__8875));
    InMux I__1804 (
            .O(N__8889),
            .I(N__8872));
    InMux I__1803 (
            .O(N__8888),
            .I(N__8865));
    InMux I__1802 (
            .O(N__8887),
            .I(N__8865));
    InMux I__1801 (
            .O(N__8886),
            .I(N__8865));
    LocalMux I__1800 (
            .O(N__8883),
            .I(beamYZ0Z_5));
    Odrv4 I__1799 (
            .O(N__8880),
            .I(beamYZ0Z_5));
    Odrv4 I__1798 (
            .O(N__8875),
            .I(beamYZ0Z_5));
    LocalMux I__1797 (
            .O(N__8872),
            .I(beamYZ0Z_5));
    LocalMux I__1796 (
            .O(N__8865),
            .I(beamYZ0Z_5));
    InMux I__1795 (
            .O(N__8854),
            .I(N__8851));
    LocalMux I__1794 (
            .O(N__8851),
            .I(un8_beamylto9_1));
    CascadeMux I__1793 (
            .O(N__8848),
            .I(N__8843));
    InMux I__1792 (
            .O(N__8847),
            .I(N__8839));
    InMux I__1791 (
            .O(N__8846),
            .I(N__8835));
    InMux I__1790 (
            .O(N__8843),
            .I(N__8832));
    InMux I__1789 (
            .O(N__8842),
            .I(N__8829));
    LocalMux I__1788 (
            .O(N__8839),
            .I(N__8823));
    InMux I__1787 (
            .O(N__8838),
            .I(N__8820));
    LocalMux I__1786 (
            .O(N__8835),
            .I(N__8813));
    LocalMux I__1785 (
            .O(N__8832),
            .I(N__8813));
    LocalMux I__1784 (
            .O(N__8829),
            .I(N__8813));
    CascadeMux I__1783 (
            .O(N__8828),
            .I(N__8809));
    CascadeMux I__1782 (
            .O(N__8827),
            .I(N__8804));
    CascadeMux I__1781 (
            .O(N__8826),
            .I(N__8801));
    Span4Mux_v I__1780 (
            .O(N__8823),
            .I(N__8794));
    LocalMux I__1779 (
            .O(N__8820),
            .I(N__8794));
    Span4Mux_v I__1778 (
            .O(N__8813),
            .I(N__8794));
    InMux I__1777 (
            .O(N__8812),
            .I(N__8791));
    InMux I__1776 (
            .O(N__8809),
            .I(N__8788));
    InMux I__1775 (
            .O(N__8808),
            .I(N__8785));
    InMux I__1774 (
            .O(N__8807),
            .I(N__8778));
    InMux I__1773 (
            .O(N__8804),
            .I(N__8778));
    InMux I__1772 (
            .O(N__8801),
            .I(N__8778));
    Odrv4 I__1771 (
            .O(N__8794),
            .I(beamYZ0Z_6));
    LocalMux I__1770 (
            .O(N__8791),
            .I(beamYZ0Z_6));
    LocalMux I__1769 (
            .O(N__8788),
            .I(beamYZ0Z_6));
    LocalMux I__1768 (
            .O(N__8785),
            .I(beamYZ0Z_6));
    LocalMux I__1767 (
            .O(N__8778),
            .I(beamYZ0Z_6));
    InMux I__1766 (
            .O(N__8767),
            .I(N__8760));
    InMux I__1765 (
            .O(N__8766),
            .I(N__8755));
    InMux I__1764 (
            .O(N__8765),
            .I(N__8755));
    InMux I__1763 (
            .O(N__8764),
            .I(N__8752));
    InMux I__1762 (
            .O(N__8763),
            .I(N__8747));
    LocalMux I__1761 (
            .O(N__8760),
            .I(N__8742));
    LocalMux I__1760 (
            .O(N__8755),
            .I(N__8742));
    LocalMux I__1759 (
            .O(N__8752),
            .I(N__8738));
    CascadeMux I__1758 (
            .O(N__8751),
            .I(N__8734));
    InMux I__1757 (
            .O(N__8750),
            .I(N__8731));
    LocalMux I__1756 (
            .O(N__8747),
            .I(N__8728));
    Span4Mux_h I__1755 (
            .O(N__8742),
            .I(N__8725));
    InMux I__1754 (
            .O(N__8741),
            .I(N__8722));
    Span4Mux_v I__1753 (
            .O(N__8738),
            .I(N__8719));
    InMux I__1752 (
            .O(N__8737),
            .I(N__8714));
    InMux I__1751 (
            .O(N__8734),
            .I(N__8714));
    LocalMux I__1750 (
            .O(N__8731),
            .I(beamYZ0Z_7));
    Odrv4 I__1749 (
            .O(N__8728),
            .I(beamYZ0Z_7));
    Odrv4 I__1748 (
            .O(N__8725),
            .I(beamYZ0Z_7));
    LocalMux I__1747 (
            .O(N__8722),
            .I(beamYZ0Z_7));
    Odrv4 I__1746 (
            .O(N__8719),
            .I(beamYZ0Z_7));
    LocalMux I__1745 (
            .O(N__8714),
            .I(beamYZ0Z_7));
    CascadeMux I__1744 (
            .O(N__8701),
            .I(Pixel_1_sqmuxa_i_cascade_));
    CascadeMux I__1743 (
            .O(N__8698),
            .I(N__8694));
    InMux I__1742 (
            .O(N__8697),
            .I(N__8689));
    InMux I__1741 (
            .O(N__8694),
            .I(N__8689));
    LocalMux I__1740 (
            .O(N__8689),
            .I(N__8686));
    Odrv4 I__1739 (
            .O(N__8686),
            .I(un1_beamx));
    IoInMux I__1738 (
            .O(N__8683),
            .I(N__8680));
    LocalMux I__1737 (
            .O(N__8680),
            .I(N__8677));
    Span4Mux_s2_v I__1736 (
            .O(N__8677),
            .I(N__8673));
    IoInMux I__1735 (
            .O(N__8676),
            .I(N__8670));
    Span4Mux_h I__1734 (
            .O(N__8673),
            .I(N__8667));
    LocalMux I__1733 (
            .O(N__8670),
            .I(N__8664));
    Sp12to4 I__1732 (
            .O(N__8667),
            .I(N__8661));
    Span4Mux_s3_v I__1731 (
            .O(N__8664),
            .I(N__8658));
    Odrv12 I__1730 (
            .O(N__8661),
            .I(HSync_c));
    Odrv4 I__1729 (
            .O(N__8658),
            .I(HSync_c));
    InMux I__1728 (
            .O(N__8653),
            .I(N__8650));
    LocalMux I__1727 (
            .O(N__8650),
            .I(un4_beamy_0));
    InMux I__1726 (
            .O(N__8647),
            .I(N__8644));
    LocalMux I__1725 (
            .O(N__8644),
            .I(N__8641));
    Odrv4 I__1724 (
            .O(N__8641),
            .I(un18_beamylt10_0));
    CascadeMux I__1723 (
            .O(N__8638),
            .I(N__8633));
    CascadeMux I__1722 (
            .O(N__8637),
            .I(N__8630));
    InMux I__1721 (
            .O(N__8636),
            .I(N__8627));
    InMux I__1720 (
            .O(N__8633),
            .I(N__8624));
    InMux I__1719 (
            .O(N__8630),
            .I(N__8620));
    LocalMux I__1718 (
            .O(N__8627),
            .I(N__8617));
    LocalMux I__1717 (
            .O(N__8624),
            .I(N__8614));
    InMux I__1716 (
            .O(N__8623),
            .I(N__8611));
    LocalMux I__1715 (
            .O(N__8620),
            .I(N__8608));
    Span4Mux_h I__1714 (
            .O(N__8617),
            .I(N__8603));
    Span4Mux_h I__1713 (
            .O(N__8614),
            .I(N__8603));
    LocalMux I__1712 (
            .O(N__8611),
            .I(beamXZ0Z_10));
    Odrv4 I__1711 (
            .O(N__8608),
            .I(beamXZ0Z_10));
    Odrv4 I__1710 (
            .O(N__8603),
            .I(beamXZ0Z_10));
    InMux I__1709 (
            .O(N__8596),
            .I(N__8593));
    LocalMux I__1708 (
            .O(N__8593),
            .I(un8_beamy));
    InMux I__1707 (
            .O(N__8590),
            .I(N__8587));
    LocalMux I__1706 (
            .O(N__8587),
            .I(un15_beamy_2));
    InMux I__1705 (
            .O(N__8584),
            .I(N__8578));
    InMux I__1704 (
            .O(N__8583),
            .I(N__8573));
    InMux I__1703 (
            .O(N__8582),
            .I(N__8573));
    InMux I__1702 (
            .O(N__8581),
            .I(N__8570));
    LocalMux I__1701 (
            .O(N__8578),
            .I(N__8565));
    LocalMux I__1700 (
            .O(N__8573),
            .I(N__8565));
    LocalMux I__1699 (
            .O(N__8570),
            .I(un1_beamx_2));
    Odrv12 I__1698 (
            .O(N__8565),
            .I(un1_beamx_2));
    InMux I__1697 (
            .O(N__8560),
            .I(N__8554));
    InMux I__1696 (
            .O(N__8559),
            .I(N__8554));
    LocalMux I__1695 (
            .O(N__8554),
            .I(N__8551));
    Odrv4 I__1694 (
            .O(N__8551),
            .I(un13_beamylt10_0));
    CascadeMux I__1693 (
            .O(N__8548),
            .I(un15_beamy_2_cascade_));
    InMux I__1692 (
            .O(N__8545),
            .I(N__8541));
    InMux I__1691 (
            .O(N__8544),
            .I(N__8538));
    LocalMux I__1690 (
            .O(N__8541),
            .I(N__8535));
    LocalMux I__1689 (
            .O(N__8538),
            .I(N__8532));
    Odrv4 I__1688 (
            .O(N__8535),
            .I(un11_visibley));
    Odrv4 I__1687 (
            .O(N__8532),
            .I(un11_visibley));
    InMux I__1686 (
            .O(N__8527),
            .I(N__8524));
    LocalMux I__1685 (
            .O(N__8524),
            .I(un27lt10));
    InMux I__1684 (
            .O(N__8521),
            .I(N__8518));
    LocalMux I__1683 (
            .O(N__8518),
            .I(un1_visiblex_27));
    CascadeMux I__1682 (
            .O(N__8515),
            .I(Pixel_9_sqmuxa_0_cascade_));
    InMux I__1681 (
            .O(N__8512),
            .I(N__8509));
    LocalMux I__1680 (
            .O(N__8509),
            .I(Pixel_9_sqmuxa));
    CascadeMux I__1679 (
            .O(N__8506),
            .I(N__8501));
    InMux I__1678 (
            .O(N__8505),
            .I(N__8496));
    InMux I__1677 (
            .O(N__8504),
            .I(N__8487));
    InMux I__1676 (
            .O(N__8501),
            .I(N__8487));
    InMux I__1675 (
            .O(N__8500),
            .I(N__8487));
    InMux I__1674 (
            .O(N__8499),
            .I(N__8487));
    LocalMux I__1673 (
            .O(N__8496),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5));
    LocalMux I__1672 (
            .O(N__8487),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5));
    InMux I__1671 (
            .O(N__8482),
            .I(N__8479));
    LocalMux I__1670 (
            .O(N__8479),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_7));
    CascadeMux I__1669 (
            .O(N__8476),
            .I(N__8471));
    InMux I__1668 (
            .O(N__8475),
            .I(N__8466));
    CascadeMux I__1667 (
            .O(N__8474),
            .I(N__8462));
    InMux I__1666 (
            .O(N__8471),
            .I(N__8458));
    CascadeMux I__1665 (
            .O(N__8470),
            .I(N__8455));
    CascadeMux I__1664 (
            .O(N__8469),
            .I(N__8451));
    LocalMux I__1663 (
            .O(N__8466),
            .I(N__8448));
    InMux I__1662 (
            .O(N__8465),
            .I(N__8445));
    InMux I__1661 (
            .O(N__8462),
            .I(N__8440));
    InMux I__1660 (
            .O(N__8461),
            .I(N__8440));
    LocalMux I__1659 (
            .O(N__8458),
            .I(N__8437));
    InMux I__1658 (
            .O(N__8455),
            .I(N__8434));
    InMux I__1657 (
            .O(N__8454),
            .I(N__8429));
    InMux I__1656 (
            .O(N__8451),
            .I(N__8429));
    Odrv4 I__1655 (
            .O(N__8448),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    LocalMux I__1654 (
            .O(N__8445),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    LocalMux I__1653 (
            .O(N__8440),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    Odrv4 I__1652 (
            .O(N__8437),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    LocalMux I__1651 (
            .O(N__8434),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    LocalMux I__1650 (
            .O(N__8429),
            .I(beamY_fast_RNI1QVSZ0Z_9));
    InMux I__1649 (
            .O(N__8416),
            .I(N__8403));
    InMux I__1648 (
            .O(N__8415),
            .I(N__8399));
    InMux I__1647 (
            .O(N__8414),
            .I(N__8394));
    InMux I__1646 (
            .O(N__8413),
            .I(N__8394));
    InMux I__1645 (
            .O(N__8412),
            .I(N__8385));
    InMux I__1644 (
            .O(N__8411),
            .I(N__8385));
    InMux I__1643 (
            .O(N__8410),
            .I(N__8385));
    InMux I__1642 (
            .O(N__8409),
            .I(N__8385));
    InMux I__1641 (
            .O(N__8408),
            .I(N__8378));
    InMux I__1640 (
            .O(N__8407),
            .I(N__8378));
    InMux I__1639 (
            .O(N__8406),
            .I(N__8378));
    LocalMux I__1638 (
            .O(N__8403),
            .I(N__8374));
    InMux I__1637 (
            .O(N__8402),
            .I(N__8371));
    LocalMux I__1636 (
            .O(N__8399),
            .I(N__8366));
    LocalMux I__1635 (
            .O(N__8394),
            .I(N__8366));
    LocalMux I__1634 (
            .O(N__8385),
            .I(N__8361));
    LocalMux I__1633 (
            .O(N__8378),
            .I(N__8361));
    InMux I__1632 (
            .O(N__8377),
            .I(N__8358));
    Span4Mux_v I__1631 (
            .O(N__8374),
            .I(N__8353));
    LocalMux I__1630 (
            .O(N__8371),
            .I(N__8353));
    Odrv4 I__1629 (
            .O(N__8366),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1628 (
            .O(N__8361),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    LocalMux I__1627 (
            .O(N__8358),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1626 (
            .O(N__8353),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    InMux I__1625 (
            .O(N__8344),
            .I(N__8334));
    InMux I__1624 (
            .O(N__8343),
            .I(N__8334));
    InMux I__1623 (
            .O(N__8342),
            .I(N__8328));
    InMux I__1622 (
            .O(N__8341),
            .I(N__8325));
    InMux I__1621 (
            .O(N__8340),
            .I(N__8321));
    InMux I__1620 (
            .O(N__8339),
            .I(N__8318));
    LocalMux I__1619 (
            .O(N__8334),
            .I(N__8315));
    InMux I__1618 (
            .O(N__8333),
            .I(N__8308));
    InMux I__1617 (
            .O(N__8332),
            .I(N__8308));
    InMux I__1616 (
            .O(N__8331),
            .I(N__8308));
    LocalMux I__1615 (
            .O(N__8328),
            .I(N__8303));
    LocalMux I__1614 (
            .O(N__8325),
            .I(N__8303));
    InMux I__1613 (
            .O(N__8324),
            .I(N__8300));
    LocalMux I__1612 (
            .O(N__8321),
            .I(N__8297));
    LocalMux I__1611 (
            .O(N__8318),
            .I(N__8288));
    Span4Mux_v I__1610 (
            .O(N__8315),
            .I(N__8288));
    LocalMux I__1609 (
            .O(N__8308),
            .I(N__8288));
    Span4Mux_v I__1608 (
            .O(N__8303),
            .I(N__8288));
    LocalMux I__1607 (
            .O(N__8300),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    Odrv4 I__1606 (
            .O(N__8297),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    Odrv4 I__1605 (
            .O(N__8288),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    InMux I__1604 (
            .O(N__8281),
            .I(N__8278));
    LocalMux I__1603 (
            .O(N__8278),
            .I(N__8275));
    Span4Mux_h I__1602 (
            .O(N__8275),
            .I(N__8272));
    Odrv4 I__1601 (
            .O(N__8272),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c4));
    CascadeMux I__1600 (
            .O(N__8269),
            .I(N__8266));
    InMux I__1599 (
            .O(N__8266),
            .I(N__8263));
    LocalMux I__1598 (
            .O(N__8263),
            .I(N__8260));
    Span4Mux_h I__1597 (
            .O(N__8260),
            .I(N__8257));
    Odrv4 I__1596 (
            .O(N__8257),
            .I(un5_visibley_c2));
    InMux I__1595 (
            .O(N__8254),
            .I(N__8251));
    LocalMux I__1594 (
            .O(N__8251),
            .I(N__8245));
    CEMux I__1593 (
            .O(N__8250),
            .I(N__8242));
    InMux I__1592 (
            .O(N__8249),
            .I(N__8238));
    CEMux I__1591 (
            .O(N__8248),
            .I(N__8235));
    Span4Mux_h I__1590 (
            .O(N__8245),
            .I(N__8230));
    LocalMux I__1589 (
            .O(N__8242),
            .I(N__8230));
    CEMux I__1588 (
            .O(N__8241),
            .I(N__8225));
    LocalMux I__1587 (
            .O(N__8238),
            .I(N__8219));
    LocalMux I__1586 (
            .O(N__8235),
            .I(N__8219));
    Span4Mux_h I__1585 (
            .O(N__8230),
            .I(N__8216));
    CEMux I__1584 (
            .O(N__8229),
            .I(N__8213));
    CEMux I__1583 (
            .O(N__8228),
            .I(N__8210));
    LocalMux I__1582 (
            .O(N__8225),
            .I(N__8207));
    CEMux I__1581 (
            .O(N__8224),
            .I(N__8204));
    Span4Mux_v I__1580 (
            .O(N__8219),
            .I(N__8196));
    Span4Mux_s3_h I__1579 (
            .O(N__8216),
            .I(N__8196));
    LocalMux I__1578 (
            .O(N__8213),
            .I(N__8196));
    LocalMux I__1577 (
            .O(N__8210),
            .I(N__8192));
    Span4Mux_s3_v I__1576 (
            .O(N__8207),
            .I(N__8187));
    LocalMux I__1575 (
            .O(N__8204),
            .I(N__8187));
    InMux I__1574 (
            .O(N__8203),
            .I(N__8184));
    Span4Mux_h I__1573 (
            .O(N__8196),
            .I(N__8181));
    InMux I__1572 (
            .O(N__8195),
            .I(N__8178));
    Span4Mux_v I__1571 (
            .O(N__8192),
            .I(N__8175));
    Span4Mux_h I__1570 (
            .O(N__8187),
            .I(N__8172));
    LocalMux I__1569 (
            .O(N__8184),
            .I(N__8167));
    Span4Mux_s3_h I__1568 (
            .O(N__8181),
            .I(N__8167));
    LocalMux I__1567 (
            .O(N__8178),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__1566 (
            .O(N__8175),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__1565 (
            .O(N__8172),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__1564 (
            .O(N__8167),
            .I(beamX_RNI5457Z0Z_5));
    InMux I__1563 (
            .O(N__8158),
            .I(N__8149));
    InMux I__1562 (
            .O(N__8157),
            .I(N__8146));
    InMux I__1561 (
            .O(N__8156),
            .I(N__8139));
    InMux I__1560 (
            .O(N__8155),
            .I(N__8139));
    InMux I__1559 (
            .O(N__8154),
            .I(N__8139));
    InMux I__1558 (
            .O(N__8153),
            .I(N__8134));
    InMux I__1557 (
            .O(N__8152),
            .I(N__8134));
    LocalMux I__1556 (
            .O(N__8149),
            .I(N__8128));
    LocalMux I__1555 (
            .O(N__8146),
            .I(N__8123));
    LocalMux I__1554 (
            .O(N__8139),
            .I(N__8123));
    LocalMux I__1553 (
            .O(N__8134),
            .I(N__8120));
    InMux I__1552 (
            .O(N__8133),
            .I(N__8113));
    InMux I__1551 (
            .O(N__8132),
            .I(N__8113));
    InMux I__1550 (
            .O(N__8131),
            .I(N__8113));
    Odrv12 I__1549 (
            .O(N__8128),
            .I(un5_beamx));
    Odrv4 I__1548 (
            .O(N__8123),
            .I(un5_beamx));
    Odrv4 I__1547 (
            .O(N__8120),
            .I(un5_beamx));
    LocalMux I__1546 (
            .O(N__8113),
            .I(un5_beamx));
    InMux I__1545 (
            .O(N__8104),
            .I(N__8099));
    InMux I__1544 (
            .O(N__8103),
            .I(N__8096));
    InMux I__1543 (
            .O(N__8102),
            .I(N__8093));
    LocalMux I__1542 (
            .O(N__8099),
            .I(N__8087));
    LocalMux I__1541 (
            .O(N__8096),
            .I(N__8087));
    LocalMux I__1540 (
            .O(N__8093),
            .I(N__8084));
    InMux I__1539 (
            .O(N__8092),
            .I(N__8081));
    Span4Mux_h I__1538 (
            .O(N__8087),
            .I(N__8078));
    Span4Mux_h I__1537 (
            .O(N__8084),
            .I(N__8075));
    LocalMux I__1536 (
            .O(N__8081),
            .I(N__8072));
    Odrv4 I__1535 (
            .O(N__8078),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1534 (
            .O(N__8075),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    Odrv12 I__1533 (
            .O(N__8072),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    InMux I__1532 (
            .O(N__8065),
            .I(N__8062));
    LocalMux I__1531 (
            .O(N__8062),
            .I(N__8056));
    InMux I__1530 (
            .O(N__8061),
            .I(N__8049));
    InMux I__1529 (
            .O(N__8060),
            .I(N__8049));
    InMux I__1528 (
            .O(N__8059),
            .I(N__8049));
    Span4Mux_v I__1527 (
            .O(N__8056),
            .I(N__8041));
    LocalMux I__1526 (
            .O(N__8049),
            .I(N__8041));
    InMux I__1525 (
            .O(N__8048),
            .I(N__8038));
    InMux I__1524 (
            .O(N__8047),
            .I(N__8035));
    InMux I__1523 (
            .O(N__8046),
            .I(N__8030));
    Span4Mux_v I__1522 (
            .O(N__8041),
            .I(N__8023));
    LocalMux I__1521 (
            .O(N__8038),
            .I(N__8023));
    LocalMux I__1520 (
            .O(N__8035),
            .I(N__8023));
    InMux I__1519 (
            .O(N__8034),
            .I(N__8020));
    InMux I__1518 (
            .O(N__8033),
            .I(N__8014));
    LocalMux I__1517 (
            .O(N__8030),
            .I(N__8007));
    Span4Mux_v I__1516 (
            .O(N__8023),
            .I(N__8007));
    LocalMux I__1515 (
            .O(N__8020),
            .I(N__8007));
    CascadeMux I__1514 (
            .O(N__8019),
            .I(N__8004));
    InMux I__1513 (
            .O(N__8018),
            .I(N__8001));
    InMux I__1512 (
            .O(N__8017),
            .I(N__7998));
    LocalMux I__1511 (
            .O(N__8014),
            .I(N__7993));
    Span4Mux_h I__1510 (
            .O(N__8007),
            .I(N__7993));
    InMux I__1509 (
            .O(N__8004),
            .I(N__7990));
    LocalMux I__1508 (
            .O(N__8001),
            .I(beamYZ0Z_3));
    LocalMux I__1507 (
            .O(N__7998),
            .I(beamYZ0Z_3));
    Odrv4 I__1506 (
            .O(N__7993),
            .I(beamYZ0Z_3));
    LocalMux I__1505 (
            .O(N__7990),
            .I(beamYZ0Z_3));
    InMux I__1504 (
            .O(N__7981),
            .I(N__7978));
    LocalMux I__1503 (
            .O(N__7978),
            .I(N__7975));
    Span4Mux_h I__1502 (
            .O(N__7975),
            .I(N__7972));
    Odrv4 I__1501 (
            .O(N__7972),
            .I(un4_beamylt6));
    CascadeMux I__1500 (
            .O(N__7969),
            .I(un4_beamylt6_cascade_));
    CascadeMux I__1499 (
            .O(N__7966),
            .I(N__7962));
    InMux I__1498 (
            .O(N__7965),
            .I(N__7955));
    InMux I__1497 (
            .O(N__7962),
            .I(N__7952));
    InMux I__1496 (
            .O(N__7961),
            .I(N__7948));
    InMux I__1495 (
            .O(N__7960),
            .I(N__7943));
    InMux I__1494 (
            .O(N__7959),
            .I(N__7943));
    InMux I__1493 (
            .O(N__7958),
            .I(N__7940));
    LocalMux I__1492 (
            .O(N__7955),
            .I(N__7933));
    LocalMux I__1491 (
            .O(N__7952),
            .I(N__7933));
    InMux I__1490 (
            .O(N__7951),
            .I(N__7927));
    LocalMux I__1489 (
            .O(N__7948),
            .I(N__7922));
    LocalMux I__1488 (
            .O(N__7943),
            .I(N__7922));
    LocalMux I__1487 (
            .O(N__7940),
            .I(N__7919));
    InMux I__1486 (
            .O(N__7939),
            .I(N__7916));
    InMux I__1485 (
            .O(N__7938),
            .I(N__7913));
    Span4Mux_h I__1484 (
            .O(N__7933),
            .I(N__7910));
    InMux I__1483 (
            .O(N__7932),
            .I(N__7907));
    InMux I__1482 (
            .O(N__7931),
            .I(N__7902));
    InMux I__1481 (
            .O(N__7930),
            .I(N__7902));
    LocalMux I__1480 (
            .O(N__7927),
            .I(N__7893));
    Span4Mux_h I__1479 (
            .O(N__7922),
            .I(N__7893));
    Span4Mux_h I__1478 (
            .O(N__7919),
            .I(N__7893));
    LocalMux I__1477 (
            .O(N__7916),
            .I(N__7893));
    LocalMux I__1476 (
            .O(N__7913),
            .I(beamYZ0Z_4));
    Odrv4 I__1475 (
            .O(N__7910),
            .I(beamYZ0Z_4));
    LocalMux I__1474 (
            .O(N__7907),
            .I(beamYZ0Z_4));
    LocalMux I__1473 (
            .O(N__7902),
            .I(beamYZ0Z_4));
    Odrv4 I__1472 (
            .O(N__7893),
            .I(beamYZ0Z_4));
    InMux I__1471 (
            .O(N__7882),
            .I(N__7877));
    InMux I__1470 (
            .O(N__7881),
            .I(N__7874));
    InMux I__1469 (
            .O(N__7880),
            .I(N__7871));
    LocalMux I__1468 (
            .O(N__7877),
            .I(N__7865));
    LocalMux I__1467 (
            .O(N__7874),
            .I(N__7862));
    LocalMux I__1466 (
            .O(N__7871),
            .I(N__7859));
    InMux I__1465 (
            .O(N__7870),
            .I(N__7856));
    CascadeMux I__1464 (
            .O(N__7869),
            .I(N__7850));
    InMux I__1463 (
            .O(N__7868),
            .I(N__7846));
    Span4Mux_h I__1462 (
            .O(N__7865),
            .I(N__7837));
    Span4Mux_v I__1461 (
            .O(N__7862),
            .I(N__7837));
    Span4Mux_v I__1460 (
            .O(N__7859),
            .I(N__7837));
    LocalMux I__1459 (
            .O(N__7856),
            .I(N__7837));
    InMux I__1458 (
            .O(N__7855),
            .I(N__7832));
    InMux I__1457 (
            .O(N__7854),
            .I(N__7832));
    InMux I__1456 (
            .O(N__7853),
            .I(N__7829));
    InMux I__1455 (
            .O(N__7850),
            .I(N__7824));
    InMux I__1454 (
            .O(N__7849),
            .I(N__7824));
    LocalMux I__1453 (
            .O(N__7846),
            .I(beamYZ0Z_8));
    Odrv4 I__1452 (
            .O(N__7837),
            .I(beamYZ0Z_8));
    LocalMux I__1451 (
            .O(N__7832),
            .I(beamYZ0Z_8));
    LocalMux I__1450 (
            .O(N__7829),
            .I(beamYZ0Z_8));
    LocalMux I__1449 (
            .O(N__7824),
            .I(beamYZ0Z_8));
    CascadeMux I__1448 (
            .O(N__7813),
            .I(un4_beamylt8_0_cascade_));
    InMux I__1447 (
            .O(N__7810),
            .I(N__7806));
    InMux I__1446 (
            .O(N__7809),
            .I(N__7802));
    LocalMux I__1445 (
            .O(N__7806),
            .I(N__7797));
    InMux I__1444 (
            .O(N__7805),
            .I(N__7794));
    LocalMux I__1443 (
            .O(N__7802),
            .I(N__7791));
    InMux I__1442 (
            .O(N__7801),
            .I(N__7788));
    InMux I__1441 (
            .O(N__7800),
            .I(N__7782));
    Span4Mux_v I__1440 (
            .O(N__7797),
            .I(N__7775));
    LocalMux I__1439 (
            .O(N__7794),
            .I(N__7775));
    Span4Mux_v I__1438 (
            .O(N__7791),
            .I(N__7775));
    LocalMux I__1437 (
            .O(N__7788),
            .I(N__7772));
    InMux I__1436 (
            .O(N__7787),
            .I(N__7769));
    InMux I__1435 (
            .O(N__7786),
            .I(N__7766));
    InMux I__1434 (
            .O(N__7785),
            .I(N__7763));
    LocalMux I__1433 (
            .O(N__7782),
            .I(beamYZ0Z_9));
    Odrv4 I__1432 (
            .O(N__7775),
            .I(beamYZ0Z_9));
    Odrv4 I__1431 (
            .O(N__7772),
            .I(beamYZ0Z_9));
    LocalMux I__1430 (
            .O(N__7769),
            .I(beamYZ0Z_9));
    LocalMux I__1429 (
            .O(N__7766),
            .I(beamYZ0Z_9));
    LocalMux I__1428 (
            .O(N__7763),
            .I(beamYZ0Z_9));
    InMux I__1427 (
            .O(N__7750),
            .I(N__7747));
    LocalMux I__1426 (
            .O(N__7747),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_7));
    CascadeMux I__1425 (
            .O(N__7744),
            .I(N__7741));
    InMux I__1424 (
            .O(N__7741),
            .I(N__7738));
    LocalMux I__1423 (
            .O(N__7738),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32));
    InMux I__1422 (
            .O(N__7735),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1421 (
            .O(N__7732),
            .I(N__7729));
    LocalMux I__1420 (
            .O(N__7729),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__1419 (
            .O(N__7726),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1418 (
            .O(N__7723),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1417 (
            .O(N__7720),
            .I(N__7717));
    LocalMux I__1416 (
            .O(N__7717),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3));
    InMux I__1415 (
            .O(N__7714),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__1414 (
            .O(N__7711),
            .I(N__7708));
    InMux I__1413 (
            .O(N__7708),
            .I(N__7705));
    LocalMux I__1412 (
            .O(N__7705),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3));
    InMux I__1411 (
            .O(N__7702),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1410 (
            .O(N__7699),
            .I(N__7696));
    InMux I__1409 (
            .O(N__7696),
            .I(N__7693));
    LocalMux I__1408 (
            .O(N__7693),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4));
    InMux I__1407 (
            .O(N__7690),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1406 (
            .O(N__7687),
            .I(N__7684));
    LocalMux I__1405 (
            .O(N__7684),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__1404 (
            .O(N__7681),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__1403 (
            .O(N__7678),
            .I(N__7674));
    CascadeMux I__1402 (
            .O(N__7677),
            .I(N__7669));
    InMux I__1401 (
            .O(N__7674),
            .I(N__7659));
    InMux I__1400 (
            .O(N__7673),
            .I(N__7659));
    InMux I__1399 (
            .O(N__7672),
            .I(N__7659));
    InMux I__1398 (
            .O(N__7669),
            .I(N__7654));
    InMux I__1397 (
            .O(N__7668),
            .I(N__7654));
    CascadeMux I__1396 (
            .O(N__7667),
            .I(N__7650));
    InMux I__1395 (
            .O(N__7666),
            .I(N__7647));
    LocalMux I__1394 (
            .O(N__7659),
            .I(N__7644));
    LocalMux I__1393 (
            .O(N__7654),
            .I(N__7641));
    InMux I__1392 (
            .O(N__7653),
            .I(N__7636));
    InMux I__1391 (
            .O(N__7650),
            .I(N__7636));
    LocalMux I__1390 (
            .O(N__7647),
            .I(N__7626));
    Span4Mux_v I__1389 (
            .O(N__7644),
            .I(N__7626));
    Span4Mux_v I__1388 (
            .O(N__7641),
            .I(N__7626));
    LocalMux I__1387 (
            .O(N__7636),
            .I(N__7626));
    InMux I__1386 (
            .O(N__7635),
            .I(N__7623));
    Span4Mux_v I__1385 (
            .O(N__7626),
            .I(N__7619));
    LocalMux I__1384 (
            .O(N__7623),
            .I(N__7616));
    InMux I__1383 (
            .O(N__7622),
            .I(N__7613));
    Odrv4 I__1382 (
            .O(N__7619),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1381 (
            .O(N__7616),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    LocalMux I__1380 (
            .O(N__7613),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1379 (
            .O(N__7606),
            .I(N__7603));
    InMux I__1378 (
            .O(N__7603),
            .I(N__7600));
    LocalMux I__1377 (
            .O(N__7600),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__1376 (
            .O(N__7597),
            .I(N__7594));
    LocalMux I__1375 (
            .O(N__7594),
            .I(N__7591));
    Odrv4 I__1374 (
            .O(N__7591),
            .I(un28_visibleylt9_0));
    InMux I__1373 (
            .O(N__7588),
            .I(N__7585));
    LocalMux I__1372 (
            .O(N__7585),
            .I(Pixel_7_sqmuxa_3_0_1));
    CascadeMux I__1371 (
            .O(N__7582),
            .I(N__7579));
    InMux I__1370 (
            .O(N__7579),
            .I(N__7576));
    LocalMux I__1369 (
            .O(N__7576),
            .I(N__7573));
    Span4Mux_h I__1368 (
            .O(N__7573),
            .I(N__7568));
    InMux I__1367 (
            .O(N__7572),
            .I(N__7565));
    InMux I__1366 (
            .O(N__7571),
            .I(N__7562));
    Odrv4 I__1365 (
            .O(N__7568),
            .I(un22_visibley_3));
    LocalMux I__1364 (
            .O(N__7565),
            .I(un22_visibley_3));
    LocalMux I__1363 (
            .O(N__7562),
            .I(un22_visibley_3));
    CascadeMux I__1362 (
            .O(N__7555),
            .I(un22_visibleylt9_0_cascade_));
    InMux I__1361 (
            .O(N__7552),
            .I(N__7545));
    InMux I__1360 (
            .O(N__7551),
            .I(N__7545));
    InMux I__1359 (
            .O(N__7550),
            .I(N__7542));
    LocalMux I__1358 (
            .O(N__7545),
            .I(N__7537));
    LocalMux I__1357 (
            .O(N__7542),
            .I(N__7537));
    Span4Mux_v I__1356 (
            .O(N__7537),
            .I(N__7534));
    Odrv4 I__1355 (
            .O(N__7534),
            .I(un22_visibley_2));
    CascadeMux I__1354 (
            .O(N__7531),
            .I(N__7528));
    InMux I__1353 (
            .O(N__7528),
            .I(N__7525));
    LocalMux I__1352 (
            .O(N__7525),
            .I(un22_visibley));
    InMux I__1351 (
            .O(N__7522),
            .I(N__7511));
    InMux I__1350 (
            .O(N__7521),
            .I(N__7511));
    InMux I__1349 (
            .O(N__7520),
            .I(N__7499));
    InMux I__1348 (
            .O(N__7519),
            .I(N__7499));
    InMux I__1347 (
            .O(N__7518),
            .I(N__7499));
    InMux I__1346 (
            .O(N__7517),
            .I(N__7495));
    InMux I__1345 (
            .O(N__7516),
            .I(N__7492));
    LocalMux I__1344 (
            .O(N__7511),
            .I(N__7489));
    InMux I__1343 (
            .O(N__7510),
            .I(N__7484));
    InMux I__1342 (
            .O(N__7509),
            .I(N__7484));
    InMux I__1341 (
            .O(N__7508),
            .I(N__7477));
    InMux I__1340 (
            .O(N__7507),
            .I(N__7477));
    InMux I__1339 (
            .O(N__7506),
            .I(N__7477));
    LocalMux I__1338 (
            .O(N__7499),
            .I(N__7474));
    InMux I__1337 (
            .O(N__7498),
            .I(N__7471));
    LocalMux I__1336 (
            .O(N__7495),
            .I(N__7466));
    LocalMux I__1335 (
            .O(N__7492),
            .I(N__7466));
    Span4Mux_v I__1334 (
            .O(N__7489),
            .I(N__7463));
    LocalMux I__1333 (
            .O(N__7484),
            .I(N__7452));
    LocalMux I__1332 (
            .O(N__7477),
            .I(N__7452));
    Span4Mux_h I__1331 (
            .O(N__7474),
            .I(N__7452));
    LocalMux I__1330 (
            .O(N__7471),
            .I(N__7452));
    Span4Mux_h I__1329 (
            .O(N__7466),
            .I(N__7452));
    Odrv4 I__1328 (
            .O(N__7463),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1327 (
            .O(N__7452),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    CascadeMux I__1326 (
            .O(N__7447),
            .I(N__7444));
    InMux I__1325 (
            .O(N__7444),
            .I(N__7441));
    LocalMux I__1324 (
            .O(N__7441),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__1323 (
            .O(N__7438),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__1322 (
            .O(N__7435),
            .I(N__7432));
    LocalMux I__1321 (
            .O(N__7432),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0));
    InMux I__1320 (
            .O(N__7429),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__1319 (
            .O(N__7426),
            .I(N__7422));
    InMux I__1318 (
            .O(N__7425),
            .I(N__7412));
    InMux I__1317 (
            .O(N__7422),
            .I(N__7412));
    InMux I__1316 (
            .O(N__7421),
            .I(N__7412));
    InMux I__1315 (
            .O(N__7420),
            .I(N__7409));
    InMux I__1314 (
            .O(N__7419),
            .I(N__7406));
    LocalMux I__1313 (
            .O(N__7412),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2));
    LocalMux I__1312 (
            .O(N__7409),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2));
    LocalMux I__1311 (
            .O(N__7406),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2));
    CascadeMux I__1310 (
            .O(N__7399),
            .I(N__7396));
    InMux I__1309 (
            .O(N__7396),
            .I(N__7393));
    LocalMux I__1308 (
            .O(N__7393),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1));
    InMux I__1307 (
            .O(N__7390),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__1306 (
            .O(N__7387),
            .I(N__7384));
    LocalMux I__1305 (
            .O(N__7384),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72));
    CascadeMux I__1304 (
            .O(N__7381),
            .I(N__7377));
    CascadeMux I__1303 (
            .O(N__7380),
            .I(N__7374));
    InMux I__1302 (
            .O(N__7377),
            .I(N__7369));
    InMux I__1301 (
            .O(N__7374),
            .I(N__7369));
    LocalMux I__1300 (
            .O(N__7369),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__1299 (
            .O(N__7366),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__1298 (
            .O(N__7363),
            .I(N__7360));
    LocalMux I__1297 (
            .O(N__7360),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__1296 (
            .O(N__7357),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__1295 (
            .O(N__7354),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_));
    CascadeMux I__1294 (
            .O(N__7351),
            .I(N__7348));
    InMux I__1293 (
            .O(N__7348),
            .I(N__7344));
    InMux I__1292 (
            .O(N__7347),
            .I(N__7341));
    LocalMux I__1291 (
            .O(N__7344),
            .I(N__7338));
    LocalMux I__1290 (
            .O(N__7341),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332));
    Odrv4 I__1289 (
            .O(N__7338),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332));
    InMux I__1288 (
            .O(N__7333),
            .I(N__7330));
    LocalMux I__1287 (
            .O(N__7330),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4));
    InMux I__1286 (
            .O(N__7327),
            .I(N__7323));
    CascadeMux I__1285 (
            .O(N__7326),
            .I(N__7319));
    LocalMux I__1284 (
            .O(N__7323),
            .I(N__7315));
    InMux I__1283 (
            .O(N__7322),
            .I(N__7312));
    InMux I__1282 (
            .O(N__7319),
            .I(N__7307));
    InMux I__1281 (
            .O(N__7318),
            .I(N__7307));
    Odrv4 I__1280 (
            .O(N__7315),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2));
    LocalMux I__1279 (
            .O(N__7312),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2));
    LocalMux I__1278 (
            .O(N__7307),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2));
    InMux I__1277 (
            .O(N__7300),
            .I(N__7297));
    LocalMux I__1276 (
            .O(N__7297),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__1275 (
            .O(N__7294),
            .I(N__7291));
    LocalMux I__1274 (
            .O(N__7291),
            .I(N__7288));
    Span4Mux_h I__1273 (
            .O(N__7288),
            .I(N__7285));
    Odrv4 I__1272 (
            .O(N__7285),
            .I(Pixel_9_sn_N_7_mux_1_tz));
    CascadeMux I__1271 (
            .O(N__7282),
            .I(un16_visibleylt9_0_cascade_));
    InMux I__1270 (
            .O(N__7279),
            .I(N__7276));
    LocalMux I__1269 (
            .O(N__7276),
            .I(N__7272));
    InMux I__1268 (
            .O(N__7275),
            .I(N__7269));
    Odrv4 I__1267 (
            .O(N__7272),
            .I(un16_visibley_4));
    LocalMux I__1266 (
            .O(N__7269),
            .I(un16_visibley_4));
    CascadeMux I__1265 (
            .O(N__7264),
            .I(N__7261));
    InMux I__1264 (
            .O(N__7261),
            .I(N__7258));
    LocalMux I__1263 (
            .O(N__7258),
            .I(N__7255));
    Odrv4 I__1262 (
            .O(N__7255),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1));
    CascadeMux I__1261 (
            .O(N__7252),
            .I(N__7249));
    InMux I__1260 (
            .O(N__7249),
            .I(N__7246));
    LocalMux I__1259 (
            .O(N__7246),
            .I(N__7243));
    Odrv4 I__1258 (
            .O(N__7243),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4));
    InMux I__1257 (
            .O(N__7240),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1256 (
            .O(N__7237),
            .I(N__7234));
    LocalMux I__1255 (
            .O(N__7234),
            .I(N__7231));
    Odrv4 I__1254 (
            .O(N__7231),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__1253 (
            .O(N__7228),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__1252 (
            .O(N__7225),
            .I(N__7222));
    LocalMux I__1251 (
            .O(N__7222),
            .I(N__7219));
    Odrv4 I__1250 (
            .O(N__7219),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__1249 (
            .O(N__7216),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__1248 (
            .O(N__7213),
            .I(N__7206));
    InMux I__1247 (
            .O(N__7212),
            .I(N__7206));
    InMux I__1246 (
            .O(N__7211),
            .I(N__7203));
    LocalMux I__1245 (
            .O(N__7206),
            .I(N__7200));
    LocalMux I__1244 (
            .O(N__7203),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5));
    Odrv4 I__1243 (
            .O(N__7200),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5));
    CascadeMux I__1242 (
            .O(N__7195),
            .I(g0_10_0_cascade_));
    InMux I__1241 (
            .O(N__7192),
            .I(N__7189));
    LocalMux I__1240 (
            .O(N__7189),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__1239 (
            .O(N__7186),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__1238 (
            .O(N__7183),
            .I(N__7179));
    InMux I__1237 (
            .O(N__7182),
            .I(N__7176));
    LocalMux I__1236 (
            .O(N__7179),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2));
    LocalMux I__1235 (
            .O(N__7176),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2));
    CascadeMux I__1234 (
            .O(N__7171),
            .I(N__7168));
    InMux I__1233 (
            .O(N__7168),
            .I(N__7165));
    LocalMux I__1232 (
            .O(N__7165),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1));
    InMux I__1231 (
            .O(N__7162),
            .I(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__1230 (
            .O(N__7159),
            .I(N__7156));
    LocalMux I__1229 (
            .O(N__7156),
            .I(N__7153));
    Odrv4 I__1228 (
            .O(N__7153),
            .I(N_7_0));
    InMux I__1227 (
            .O(N__7150),
            .I(N__7147));
    LocalMux I__1226 (
            .O(N__7147),
            .I(N__7144));
    Span4Mux_v I__1225 (
            .O(N__7144),
            .I(N__7141));
    Odrv4 I__1224 (
            .O(N__7141),
            .I(G_25_i_a8_1_1));
    CascadeMux I__1223 (
            .O(N__7138),
            .I(N__7135));
    InMux I__1222 (
            .O(N__7135),
            .I(N__7132));
    LocalMux I__1221 (
            .O(N__7132),
            .I(N__7128));
    InMux I__1220 (
            .O(N__7131),
            .I(N__7125));
    Odrv4 I__1219 (
            .O(N__7128),
            .I(G_25_i_o8_0_2));
    LocalMux I__1218 (
            .O(N__7125),
            .I(G_25_i_o8_0_2));
    InMux I__1217 (
            .O(N__7120),
            .I(N__7114));
    InMux I__1216 (
            .O(N__7119),
            .I(N__7114));
    LocalMux I__1215 (
            .O(N__7114),
            .I(Pixel_7_sqmuxa_1));
    CascadeMux I__1214 (
            .O(N__7111),
            .I(N__7108));
    InMux I__1213 (
            .O(N__7108),
            .I(N__7105));
    LocalMux I__1212 (
            .O(N__7105),
            .I(N__7102));
    Odrv4 I__1211 (
            .O(N__7102),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03));
    InMux I__1210 (
            .O(N__7099),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1209 (
            .O(N__7096),
            .I(r_i1_mux_cascade_));
    InMux I__1208 (
            .O(N__7093),
            .I(N__7090));
    LocalMux I__1207 (
            .O(N__7090),
            .I(font_un78_pixellto3));
    CascadeMux I__1206 (
            .O(N__7087),
            .I(Pixel_3_sqmuxa_1_1_cascade_));
    InMux I__1205 (
            .O(N__7084),
            .I(N__7081));
    LocalMux I__1204 (
            .O(N__7081),
            .I(N__7078));
    Odrv4 I__1203 (
            .O(N__7078),
            .I(G_25_i_a8_0_0));
    CascadeMux I__1202 (
            .O(N__7075),
            .I(Pixel_7_sqmuxa_1_cascade_));
    CascadeMux I__1201 (
            .O(N__7072),
            .I(N__7069));
    InMux I__1200 (
            .O(N__7069),
            .I(N__7066));
    LocalMux I__1199 (
            .O(N__7066),
            .I(N__7063));
    Span4Mux_h I__1198 (
            .O(N__7063),
            .I(N__7060));
    Odrv4 I__1197 (
            .O(N__7060),
            .I(g0_0_0_1));
    InMux I__1196 (
            .O(N__7057),
            .I(N__7054));
    LocalMux I__1195 (
            .O(N__7054),
            .I(g1));
    CascadeMux I__1194 (
            .O(N__7051),
            .I(g0_0_4_0_cascade_));
    InMux I__1193 (
            .O(N__7048),
            .I(N__7045));
    LocalMux I__1192 (
            .O(N__7045),
            .I(N_11));
    InMux I__1191 (
            .O(N__7042),
            .I(N__7039));
    LocalMux I__1190 (
            .O(N__7039),
            .I(g0_0_2));
    InMux I__1189 (
            .O(N__7036),
            .I(N__7030));
    InMux I__1188 (
            .O(N__7035),
            .I(N__7030));
    LocalMux I__1187 (
            .O(N__7030),
            .I(Pixel_3_sqmuxa_1_1));
    InMux I__1186 (
            .O(N__7027),
            .I(N__7016));
    InMux I__1185 (
            .O(N__7026),
            .I(N__7016));
    InMux I__1184 (
            .O(N__7025),
            .I(N__7016));
    InMux I__1183 (
            .O(N__7024),
            .I(N__7011));
    InMux I__1182 (
            .O(N__7023),
            .I(N__7011));
    LocalMux I__1181 (
            .O(N__7016),
            .I(N__7008));
    LocalMux I__1180 (
            .O(N__7011),
            .I(beamY_RNIECTA3Z0Z_8));
    Odrv4 I__1179 (
            .O(N__7008),
            .I(beamY_RNIECTA3Z0Z_8));
    CascadeMux I__1178 (
            .O(N__7003),
            .I(N__6996));
    InMux I__1177 (
            .O(N__7002),
            .I(N__6985));
    InMux I__1176 (
            .O(N__7001),
            .I(N__6985));
    InMux I__1175 (
            .O(N__7000),
            .I(N__6985));
    InMux I__1174 (
            .O(N__6999),
            .I(N__6985));
    InMux I__1173 (
            .O(N__6996),
            .I(N__6982));
    InMux I__1172 (
            .O(N__6995),
            .I(N__6977));
    InMux I__1171 (
            .O(N__6994),
            .I(N__6977));
    LocalMux I__1170 (
            .O(N__6985),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5));
    LocalMux I__1169 (
            .O(N__6982),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5));
    LocalMux I__1168 (
            .O(N__6977),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5));
    CascadeMux I__1167 (
            .O(N__6970),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_));
    InMux I__1166 (
            .O(N__6967),
            .I(N__6964));
    LocalMux I__1165 (
            .O(N__6964),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2));
    InMux I__1164 (
            .O(N__6961),
            .I(N__6958));
    LocalMux I__1163 (
            .O(N__6958),
            .I(un1_beamylto9_1));
    InMux I__1162 (
            .O(N__6955),
            .I(N__6949));
    InMux I__1161 (
            .O(N__6954),
            .I(N__6949));
    LocalMux I__1160 (
            .O(N__6949),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0));
    InMux I__1159 (
            .O(N__6946),
            .I(N__6940));
    InMux I__1158 (
            .O(N__6945),
            .I(N__6940));
    LocalMux I__1157 (
            .O(N__6940),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5));
    InMux I__1156 (
            .O(N__6937),
            .I(N__6934));
    LocalMux I__1155 (
            .O(N__6934),
            .I(Pixel_1_esr_RNOZ0Z_60));
    CascadeMux I__1154 (
            .O(N__6931),
            .I(g1_0_cascade_));
    CascadeMux I__1153 (
            .O(N__6928),
            .I(N__6925));
    InMux I__1152 (
            .O(N__6925),
            .I(N__6922));
    LocalMux I__1151 (
            .O(N__6922),
            .I(N__6919));
    Odrv12 I__1150 (
            .O(N__6919),
            .I(un1_beamxlt10_0));
    InMux I__1149 (
            .O(N__6916),
            .I(N__6913));
    LocalMux I__1148 (
            .O(N__6913),
            .I(N__6907));
    CascadeMux I__1147 (
            .O(N__6912),
            .I(N__6904));
    InMux I__1146 (
            .O(N__6911),
            .I(N__6899));
    InMux I__1145 (
            .O(N__6910),
            .I(N__6896));
    Span4Mux_h I__1144 (
            .O(N__6907),
            .I(N__6893));
    InMux I__1143 (
            .O(N__6904),
            .I(N__6888));
    InMux I__1142 (
            .O(N__6903),
            .I(N__6888));
    InMux I__1141 (
            .O(N__6902),
            .I(N__6885));
    LocalMux I__1140 (
            .O(N__6899),
            .I(beamXZ0Z_7));
    LocalMux I__1139 (
            .O(N__6896),
            .I(beamXZ0Z_7));
    Odrv4 I__1138 (
            .O(N__6893),
            .I(beamXZ0Z_7));
    LocalMux I__1137 (
            .O(N__6888),
            .I(beamXZ0Z_7));
    LocalMux I__1136 (
            .O(N__6885),
            .I(beamXZ0Z_7));
    CascadeMux I__1135 (
            .O(N__6874),
            .I(N__6869));
    InMux I__1134 (
            .O(N__6873),
            .I(N__6862));
    InMux I__1133 (
            .O(N__6872),
            .I(N__6862));
    InMux I__1132 (
            .O(N__6869),
            .I(N__6862));
    LocalMux I__1131 (
            .O(N__6862),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0));
    CascadeMux I__1130 (
            .O(N__6859),
            .I(N__6856));
    InMux I__1129 (
            .O(N__6856),
            .I(N__6846));
    InMux I__1128 (
            .O(N__6855),
            .I(N__6846));
    InMux I__1127 (
            .O(N__6854),
            .I(N__6846));
    InMux I__1126 (
            .O(N__6853),
            .I(N__6843));
    LocalMux I__1125 (
            .O(N__6846),
            .I(beamY_RNIAJLT9AZ0Z_3));
    LocalMux I__1124 (
            .O(N__6843),
            .I(beamY_RNIAJLT9AZ0Z_3));
    InMux I__1123 (
            .O(N__6838),
            .I(N__6835));
    LocalMux I__1122 (
            .O(N__6835),
            .I(N__6832));
    Span4Mux_h I__1121 (
            .O(N__6832),
            .I(N__6828));
    InMux I__1120 (
            .O(N__6831),
            .I(N__6825));
    Odrv4 I__1119 (
            .O(N__6828),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    LocalMux I__1118 (
            .O(N__6825),
            .I(un21_beamy_cry_5_c_RNII1CZ0Z3));
    InMux I__1117 (
            .O(N__6820),
            .I(N__6815));
    InMux I__1116 (
            .O(N__6819),
            .I(N__6812));
    InMux I__1115 (
            .O(N__6818),
            .I(N__6809));
    LocalMux I__1114 (
            .O(N__6815),
            .I(beamY_fastZ0Z_6));
    LocalMux I__1113 (
            .O(N__6812),
            .I(beamY_fastZ0Z_6));
    LocalMux I__1112 (
            .O(N__6809),
            .I(beamY_fastZ0Z_6));
    InMux I__1111 (
            .O(N__6802),
            .I(N__6799));
    LocalMux I__1110 (
            .O(N__6799),
            .I(N__6795));
    InMux I__1109 (
            .O(N__6798),
            .I(N__6792));
    Odrv4 I__1108 (
            .O(N__6795),
            .I(un5_visibley_c6_0_0));
    LocalMux I__1107 (
            .O(N__6792),
            .I(un5_visibley_c6_0_0));
    InMux I__1106 (
            .O(N__6787),
            .I(N__6784));
    LocalMux I__1105 (
            .O(N__6784),
            .I(N__6781));
    Span4Mux_h I__1104 (
            .O(N__6781),
            .I(N__6777));
    InMux I__1103 (
            .O(N__6780),
            .I(N__6774));
    Odrv4 I__1102 (
            .O(N__6777),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    LocalMux I__1101 (
            .O(N__6774),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    InMux I__1100 (
            .O(N__6769),
            .I(N__6763));
    InMux I__1099 (
            .O(N__6768),
            .I(N__6763));
    LocalMux I__1098 (
            .O(N__6763),
            .I(N__6759));
    InMux I__1097 (
            .O(N__6762),
            .I(N__6754));
    Span4Mux_h I__1096 (
            .O(N__6759),
            .I(N__6751));
    InMux I__1095 (
            .O(N__6758),
            .I(N__6748));
    InMux I__1094 (
            .O(N__6757),
            .I(N__6745));
    LocalMux I__1093 (
            .O(N__6754),
            .I(beamY_fastZ0Z_5));
    Odrv4 I__1092 (
            .O(N__6751),
            .I(beamY_fastZ0Z_5));
    LocalMux I__1091 (
            .O(N__6748),
            .I(beamY_fastZ0Z_5));
    LocalMux I__1090 (
            .O(N__6745),
            .I(beamY_fastZ0Z_5));
    InMux I__1089 (
            .O(N__6736),
            .I(N__6730));
    InMux I__1088 (
            .O(N__6735),
            .I(N__6724));
    InMux I__1087 (
            .O(N__6734),
            .I(N__6721));
    InMux I__1086 (
            .O(N__6733),
            .I(N__6718));
    LocalMux I__1085 (
            .O(N__6730),
            .I(N__6715));
    InMux I__1084 (
            .O(N__6729),
            .I(N__6712));
    InMux I__1083 (
            .O(N__6728),
            .I(N__6709));
    InMux I__1082 (
            .O(N__6727),
            .I(N__6706));
    LocalMux I__1081 (
            .O(N__6724),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__1080 (
            .O(N__6721),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__1079 (
            .O(N__6718),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    Odrv4 I__1078 (
            .O(N__6715),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__1077 (
            .O(N__6712),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__1076 (
            .O(N__6709),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    LocalMux I__1075 (
            .O(N__6706),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum));
    InMux I__1074 (
            .O(N__6691),
            .I(N__6686));
    InMux I__1073 (
            .O(N__6690),
            .I(N__6681));
    InMux I__1072 (
            .O(N__6689),
            .I(N__6677));
    LocalMux I__1071 (
            .O(N__6686),
            .I(N__6674));
    InMux I__1070 (
            .O(N__6685),
            .I(N__6671));
    InMux I__1069 (
            .O(N__6684),
            .I(N__6668));
    LocalMux I__1068 (
            .O(N__6681),
            .I(N__6665));
    InMux I__1067 (
            .O(N__6680),
            .I(N__6662));
    LocalMux I__1066 (
            .O(N__6677),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    Odrv4 I__1065 (
            .O(N__6674),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    LocalMux I__1064 (
            .O(N__6671),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    LocalMux I__1063 (
            .O(N__6668),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    Odrv4 I__1062 (
            .O(N__6665),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    LocalMux I__1061 (
            .O(N__6662),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    CascadeMux I__1060 (
            .O(N__6649),
            .I(beamY_RNIECTA3Z0Z_8_cascade_));
    InMux I__1059 (
            .O(N__6646),
            .I(N__6642));
    InMux I__1058 (
            .O(N__6645),
            .I(N__6639));
    LocalMux I__1057 (
            .O(N__6642),
            .I(N__6632));
    LocalMux I__1056 (
            .O(N__6639),
            .I(N__6632));
    InMux I__1055 (
            .O(N__6638),
            .I(N__6627));
    InMux I__1054 (
            .O(N__6637),
            .I(N__6627));
    Odrv4 I__1053 (
            .O(N__6632),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3));
    LocalMux I__1052 (
            .O(N__6627),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3));
    CascadeMux I__1051 (
            .O(N__6622),
            .I(N__6619));
    InMux I__1050 (
            .O(N__6619),
            .I(N__6616));
    LocalMux I__1049 (
            .O(N__6616),
            .I(N__6613));
    Odrv12 I__1048 (
            .O(N__6613),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1));
    CascadeMux I__1047 (
            .O(N__6610),
            .I(N__6607));
    InMux I__1046 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__1045 (
            .O(N__6604),
            .I(un1_beamylto9_2));
    InMux I__1044 (
            .O(N__6601),
            .I(N__6598));
    LocalMux I__1043 (
            .O(N__6598),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0));
    InMux I__1042 (
            .O(N__6595),
            .I(N__6592));
    LocalMux I__1041 (
            .O(N__6592),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1));
    CascadeMux I__1040 (
            .O(N__6589),
            .I(N__6586));
    InMux I__1039 (
            .O(N__6586),
            .I(N__6583));
    LocalMux I__1038 (
            .O(N__6583),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1));
    InMux I__1037 (
            .O(N__6580),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__1036 (
            .O(N__6577),
            .I(N__6574));
    LocalMux I__1035 (
            .O(N__6574),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1));
    CascadeMux I__1034 (
            .O(N__6571),
            .I(N__6568));
    InMux I__1033 (
            .O(N__6568),
            .I(N__6565));
    LocalMux I__1032 (
            .O(N__6565),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1));
    InMux I__1031 (
            .O(N__6562),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__1030 (
            .O(N__6559),
            .I(N__6555));
    InMux I__1029 (
            .O(N__6558),
            .I(N__6551));
    InMux I__1028 (
            .O(N__6555),
            .I(N__6548));
    InMux I__1027 (
            .O(N__6554),
            .I(N__6545));
    LocalMux I__1026 (
            .O(N__6551),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__1025 (
            .O(N__6548),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__1024 (
            .O(N__6545),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    InMux I__1023 (
            .O(N__6538),
            .I(N__6535));
    LocalMux I__1022 (
            .O(N__6535),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__1021 (
            .O(N__6532),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__1020 (
            .O(N__6529),
            .I(N__6526));
    LocalMux I__1019 (
            .O(N__6526),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__1018 (
            .O(N__6523),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__1017 (
            .O(N__6520),
            .I(N__6515));
    InMux I__1016 (
            .O(N__6519),
            .I(N__6505));
    InMux I__1015 (
            .O(N__6518),
            .I(N__6505));
    InMux I__1014 (
            .O(N__6515),
            .I(N__6505));
    InMux I__1013 (
            .O(N__6514),
            .I(N__6505));
    LocalMux I__1012 (
            .O(N__6505),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0));
    CascadeMux I__1011 (
            .O(N__6502),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_));
    InMux I__1010 (
            .O(N__6499),
            .I(N__6496));
    LocalMux I__1009 (
            .O(N__6496),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_7));
    CascadeMux I__1008 (
            .O(N__6493),
            .I(N__6490));
    InMux I__1007 (
            .O(N__6490),
            .I(N__6485));
    InMux I__1006 (
            .O(N__6489),
            .I(N__6482));
    InMux I__1005 (
            .O(N__6488),
            .I(N__6479));
    LocalMux I__1004 (
            .O(N__6485),
            .I(beamY_fastZ0Z_7));
    LocalMux I__1003 (
            .O(N__6482),
            .I(beamY_fastZ0Z_7));
    LocalMux I__1002 (
            .O(N__6479),
            .I(beamY_fastZ0Z_7));
    InMux I__1001 (
            .O(N__6472),
            .I(N__6469));
    LocalMux I__1000 (
            .O(N__6469),
            .I(un5_visibley_c6_0_0_0));
    CascadeMux I__999 (
            .O(N__6466),
            .I(un11_visibleylto9_1_cascade_));
    CascadeMux I__998 (
            .O(N__6463),
            .I(un11_visibleylto9_4_cascade_));
    CascadeMux I__997 (
            .O(N__6460),
            .I(N__6457));
    InMux I__996 (
            .O(N__6457),
            .I(N__6454));
    LocalMux I__995 (
            .O(N__6454),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1));
    InMux I__994 (
            .O(N__6451),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3));
    CascadeMux I__993 (
            .O(N__6448),
            .I(N__6445));
    InMux I__992 (
            .O(N__6445),
            .I(N__6442));
    LocalMux I__991 (
            .O(N__6442),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1));
    InMux I__990 (
            .O(N__6439),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__989 (
            .O(N__6436),
            .I(N__6433));
    LocalMux I__988 (
            .O(N__6433),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__987 (
            .O(N__6430),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__986 (
            .O(N__6427),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__985 (
            .O(N__6424),
            .I(N__6420));
    InMux I__984 (
            .O(N__6423),
            .I(N__6411));
    InMux I__983 (
            .O(N__6420),
            .I(N__6411));
    InMux I__982 (
            .O(N__6419),
            .I(N__6411));
    InMux I__981 (
            .O(N__6418),
            .I(N__6408));
    LocalMux I__980 (
            .O(N__6411),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    LocalMux I__979 (
            .O(N__6408),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    CascadeMux I__978 (
            .O(N__6403),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_));
    InMux I__977 (
            .O(N__6400),
            .I(N__6397));
    LocalMux I__976 (
            .O(N__6397),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__975 (
            .O(N__6394),
            .I(N__6391));
    InMux I__974 (
            .O(N__6391),
            .I(N__6388));
    LocalMux I__973 (
            .O(N__6388),
            .I(beamY_RNI9KEQ_0Z0Z_8));
    InMux I__972 (
            .O(N__6385),
            .I(N__6382));
    LocalMux I__971 (
            .O(N__6382),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0));
    InMux I__970 (
            .O(N__6379),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__969 (
            .O(N__6376),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__968 (
            .O(N__6373),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__967 (
            .O(N__6370),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__966 (
            .O(N__6367),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__965 (
            .O(N__6364),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__964 (
            .O(N__6361),
            .I(N__6358));
    InMux I__963 (
            .O(N__6358),
            .I(N__6355));
    LocalMux I__962 (
            .O(N__6355),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_0));
    CascadeMux I__961 (
            .O(N__6352),
            .I(N__6349));
    InMux I__960 (
            .O(N__6349),
            .I(N__6346));
    LocalMux I__959 (
            .O(N__6346),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__958 (
            .O(N__6343),
            .I(N__6340));
    LocalMux I__957 (
            .O(N__6340),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0));
    InMux I__956 (
            .O(N__6337),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__955 (
            .O(N__6334),
            .I(N__6331));
    LocalMux I__954 (
            .O(N__6331),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_i));
    InMux I__953 (
            .O(N__6328),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__952 (
            .O(N__6325),
            .I(N__6321));
    InMux I__951 (
            .O(N__6324),
            .I(N__6318));
    LocalMux I__950 (
            .O(N__6321),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31));
    LocalMux I__949 (
            .O(N__6318),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31));
    CascadeMux I__948 (
            .O(N__6313),
            .I(N__6310));
    InMux I__947 (
            .O(N__6310),
            .I(N__6307));
    LocalMux I__946 (
            .O(N__6307),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0));
    InMux I__945 (
            .O(N__6304),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__944 (
            .O(N__6301),
            .I(N__6295));
    InMux I__943 (
            .O(N__6300),
            .I(N__6295));
    LocalMux I__942 (
            .O(N__6295),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__941 (
            .O(N__6292),
            .I(N__6289));
    InMux I__940 (
            .O(N__6289),
            .I(N__6286));
    LocalMux I__939 (
            .O(N__6286),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831));
    InMux I__938 (
            .O(N__6283),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__937 (
            .O(N__6280),
            .I(N__6277));
    LocalMux I__936 (
            .O(N__6277),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__935 (
            .O(N__6274),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__934 (
            .O(N__6271),
            .I(N__6267));
    CascadeMux I__933 (
            .O(N__6270),
            .I(N__6264));
    LocalMux I__932 (
            .O(N__6267),
            .I(N__6258));
    InMux I__931 (
            .O(N__6264),
            .I(N__6255));
    InMux I__930 (
            .O(N__6263),
            .I(N__6249));
    InMux I__929 (
            .O(N__6262),
            .I(N__6244));
    InMux I__928 (
            .O(N__6261),
            .I(N__6244));
    Span4Mux_v I__927 (
            .O(N__6258),
            .I(N__6241));
    LocalMux I__926 (
            .O(N__6255),
            .I(N__6238));
    InMux I__925 (
            .O(N__6254),
            .I(N__6235));
    InMux I__924 (
            .O(N__6253),
            .I(N__6230));
    InMux I__923 (
            .O(N__6252),
            .I(N__6230));
    LocalMux I__922 (
            .O(N__6249),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__921 (
            .O(N__6244),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    Odrv4 I__920 (
            .O(N__6241),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    Odrv12 I__919 (
            .O(N__6238),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__918 (
            .O(N__6235),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    LocalMux I__917 (
            .O(N__6230),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    CascadeMux I__916 (
            .O(N__6217),
            .I(N__6214));
    InMux I__915 (
            .O(N__6214),
            .I(N__6211));
    LocalMux I__914 (
            .O(N__6211),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i));
    InMux I__913 (
            .O(N__6208),
            .I(N__6205));
    LocalMux I__912 (
            .O(N__6205),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__911 (
            .O(N__6202),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__910 (
            .O(N__6199),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_));
    InMux I__909 (
            .O(N__6196),
            .I(N__6188));
    InMux I__908 (
            .O(N__6195),
            .I(N__6181));
    InMux I__907 (
            .O(N__6194),
            .I(N__6181));
    InMux I__906 (
            .O(N__6193),
            .I(N__6176));
    InMux I__905 (
            .O(N__6192),
            .I(N__6176));
    InMux I__904 (
            .O(N__6191),
            .I(N__6173));
    LocalMux I__903 (
            .O(N__6188),
            .I(N__6170));
    InMux I__902 (
            .O(N__6187),
            .I(N__6167));
    InMux I__901 (
            .O(N__6186),
            .I(N__6164));
    LocalMux I__900 (
            .O(N__6181),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__899 (
            .O(N__6176),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__898 (
            .O(N__6173),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    Odrv4 I__897 (
            .O(N__6170),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__896 (
            .O(N__6167),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    LocalMux I__895 (
            .O(N__6164),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    CascadeMux I__894 (
            .O(N__6151),
            .I(N__6148));
    InMux I__893 (
            .O(N__6148),
            .I(N__6144));
    CascadeMux I__892 (
            .O(N__6147),
            .I(N__6141));
    LocalMux I__891 (
            .O(N__6144),
            .I(N__6138));
    InMux I__890 (
            .O(N__6141),
            .I(N__6135));
    Odrv4 I__889 (
            .O(N__6138),
            .I(un5_visiblex_i_24));
    LocalMux I__888 (
            .O(N__6135),
            .I(un5_visiblex_i_24));
    InMux I__887 (
            .O(N__6130),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1));
    InMux I__886 (
            .O(N__6127),
            .I(N__6123));
    InMux I__885 (
            .O(N__6126),
            .I(N__6120));
    LocalMux I__884 (
            .O(N__6123),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1));
    LocalMux I__883 (
            .O(N__6120),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1));
    CascadeMux I__882 (
            .O(N__6115),
            .I(N__6112));
    InMux I__881 (
            .O(N__6112),
            .I(N__6109));
    LocalMux I__880 (
            .O(N__6109),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0));
    InMux I__879 (
            .O(N__6106),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__878 (
            .O(N__6103),
            .I(N__6100));
    LocalMux I__877 (
            .O(N__6100),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41));
    CascadeMux I__876 (
            .O(N__6097),
            .I(N__6093));
    CascadeMux I__875 (
            .O(N__6096),
            .I(N__6090));
    InMux I__874 (
            .O(N__6093),
            .I(N__6085));
    InMux I__873 (
            .O(N__6090),
            .I(N__6085));
    LocalMux I__872 (
            .O(N__6085),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5));
    InMux I__871 (
            .O(N__6082),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__870 (
            .O(N__6079),
            .I(N__6076));
    LocalMux I__869 (
            .O(N__6076),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__868 (
            .O(N__6073),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__867 (
            .O(N__6070),
            .I(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_));
    InMux I__866 (
            .O(N__6067),
            .I(N__6064));
    LocalMux I__865 (
            .O(N__6064),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO));
    InMux I__864 (
            .O(N__6061),
            .I(N__6055));
    InMux I__863 (
            .O(N__6060),
            .I(N__6055));
    LocalMux I__862 (
            .O(N__6055),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3));
    InMux I__861 (
            .O(N__6052),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__860 (
            .O(N__6049),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_));
    InMux I__859 (
            .O(N__6046),
            .I(N__6043));
    LocalMux I__858 (
            .O(N__6043),
            .I(un22_visibleylt9_0_0_0));
    InMux I__857 (
            .O(N__6040),
            .I(N__6037));
    LocalMux I__856 (
            .O(N__6037),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_i));
    InMux I__855 (
            .O(N__6034),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1));
    InMux I__854 (
            .O(N__6031),
            .I(N__6027));
    InMux I__853 (
            .O(N__6030),
            .I(N__6024));
    LocalMux I__852 (
            .O(N__6027),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0));
    LocalMux I__851 (
            .O(N__6024),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0));
    CascadeMux I__850 (
            .O(N__6019),
            .I(N__6016));
    InMux I__849 (
            .O(N__6016),
            .I(N__6013));
    LocalMux I__848 (
            .O(N__6013),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0));
    InMux I__847 (
            .O(N__6010),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__846 (
            .O(N__6007),
            .I(N__6004));
    LocalMux I__845 (
            .O(N__6004),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0));
    CascadeMux I__844 (
            .O(N__6001),
            .I(N__5997));
    CascadeMux I__843 (
            .O(N__6000),
            .I(N__5994));
    InMux I__842 (
            .O(N__5997),
            .I(N__5989));
    InMux I__841 (
            .O(N__5994),
            .I(N__5989));
    LocalMux I__840 (
            .O(N__5989),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5));
    InMux I__839 (
            .O(N__5986),
            .I(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__838 (
            .O(N__5983),
            .I(N__5977));
    InMux I__837 (
            .O(N__5982),
            .I(N__5977));
    LocalMux I__836 (
            .O(N__5977),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__835 (
            .O(N__5974),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__834 (
            .O(N__5971),
            .I(N__5967));
    InMux I__833 (
            .O(N__5970),
            .I(N__5964));
    LocalMux I__832 (
            .O(N__5967),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    LocalMux I__831 (
            .O(N__5964),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO));
    InMux I__830 (
            .O(N__5959),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1));
    CascadeMux I__829 (
            .O(N__5956),
            .I(N__5953));
    InMux I__828 (
            .O(N__5953),
            .I(N__5950));
    LocalMux I__827 (
            .O(N__5950),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5));
    InMux I__826 (
            .O(N__5947),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__825 (
            .O(N__5944),
            .I(N__5940));
    InMux I__824 (
            .O(N__5943),
            .I(N__5937));
    LocalMux I__823 (
            .O(N__5940),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06));
    LocalMux I__822 (
            .O(N__5937),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06));
    CascadeMux I__821 (
            .O(N__5932),
            .I(N__5929));
    InMux I__820 (
            .O(N__5929),
            .I(N__5926));
    LocalMux I__819 (
            .O(N__5926),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9));
    InMux I__818 (
            .O(N__5923),
            .I(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__817 (
            .O(N__5920),
            .I(N__5914));
    InMux I__816 (
            .O(N__5919),
            .I(N__5911));
    InMux I__815 (
            .O(N__5918),
            .I(N__5906));
    InMux I__814 (
            .O(N__5917),
            .I(N__5906));
    LocalMux I__813 (
            .O(N__5914),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__812 (
            .O(N__5911),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c5));
    LocalMux I__811 (
            .O(N__5906),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c5));
    CascadeMux I__810 (
            .O(N__5899),
            .I(beamY_RNI5F8A81Z0Z_3_cascade_));
    InMux I__809 (
            .O(N__5896),
            .I(N__5887));
    InMux I__808 (
            .O(N__5895),
            .I(N__5887));
    InMux I__807 (
            .O(N__5894),
            .I(N__5884));
    InMux I__806 (
            .O(N__5893),
            .I(N__5879));
    InMux I__805 (
            .O(N__5892),
            .I(N__5879));
    LocalMux I__804 (
            .O(N__5887),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i));
    LocalMux I__803 (
            .O(N__5884),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i));
    LocalMux I__802 (
            .O(N__5879),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i));
    InMux I__801 (
            .O(N__5872),
            .I(N__5869));
    LocalMux I__800 (
            .O(N__5869),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0));
    CascadeMux I__799 (
            .O(N__5866),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_));
    InMux I__798 (
            .O(N__5863),
            .I(N__5860));
    LocalMux I__797 (
            .O(N__5860),
            .I(beamY_RNIKUC181_0Z0Z_5));
    CascadeMux I__796 (
            .O(N__5857),
            .I(N__5854));
    InMux I__795 (
            .O(N__5854),
            .I(N__5848));
    InMux I__794 (
            .O(N__5853),
            .I(N__5848));
    LocalMux I__793 (
            .O(N__5848),
            .I(beamY_RNIKPNA02Z0Z_5));
    InMux I__792 (
            .O(N__5845),
            .I(N__5839));
    InMux I__791 (
            .O(N__5844),
            .I(N__5839));
    LocalMux I__790 (
            .O(N__5839),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3));
    InMux I__789 (
            .O(N__5836),
            .I(N__5832));
    InMux I__788 (
            .O(N__5835),
            .I(N__5829));
    LocalMux I__787 (
            .O(N__5832),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11));
    LocalMux I__786 (
            .O(N__5829),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11));
    CascadeMux I__785 (
            .O(N__5824),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_));
    InMux I__784 (
            .O(N__5821),
            .I(N__5818));
    LocalMux I__783 (
            .O(N__5818),
            .I(N__5815));
    Span4Mux_h I__782 (
            .O(N__5815),
            .I(N__5811));
    InMux I__781 (
            .O(N__5814),
            .I(N__5808));
    Odrv4 I__780 (
            .O(N__5811),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10));
    LocalMux I__779 (
            .O(N__5808),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10));
    InMux I__778 (
            .O(N__5803),
            .I(N__5800));
    LocalMux I__777 (
            .O(N__5800),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_c4));
    InMux I__776 (
            .O(N__5797),
            .I(N__5794));
    LocalMux I__775 (
            .O(N__5794),
            .I(font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0));
    CascadeMux I__774 (
            .O(N__5791),
            .I(N__5787));
    InMux I__773 (
            .O(N__5790),
            .I(N__5782));
    InMux I__772 (
            .O(N__5787),
            .I(N__5782));
    LocalMux I__771 (
            .O(N__5782),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i));
    CascadeMux I__770 (
            .O(N__5779),
            .I(N__5776));
    InMux I__769 (
            .O(N__5776),
            .I(N__5773));
    LocalMux I__768 (
            .O(N__5773),
            .I(N__5770));
    Span4Mux_h I__767 (
            .O(N__5770),
            .I(N__5767));
    Odrv4 I__766 (
            .O(N__5767),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i));
    InMux I__765 (
            .O(N__5764),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__764 (
            .O(N__5761),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__763 (
            .O(N__5758),
            .I(N__5751));
    InMux I__762 (
            .O(N__5757),
            .I(N__5751));
    InMux I__761 (
            .O(N__5756),
            .I(N__5748));
    LocalMux I__760 (
            .O(N__5751),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux));
    LocalMux I__759 (
            .O(N__5748),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux));
    CascadeMux I__758 (
            .O(N__5743),
            .I(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_));
    CascadeMux I__757 (
            .O(N__5740),
            .I(N__5737));
    InMux I__756 (
            .O(N__5737),
            .I(N__5734));
    LocalMux I__755 (
            .O(N__5734),
            .I(N__5730));
    InMux I__754 (
            .O(N__5733),
            .I(N__5727));
    Odrv4 I__753 (
            .O(N__5730),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6));
    LocalMux I__752 (
            .O(N__5727),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6));
    CascadeMux I__751 (
            .O(N__5722),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_));
    CascadeMux I__750 (
            .O(N__5719),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_));
    InMux I__749 (
            .O(N__5716),
            .I(N__5713));
    LocalMux I__748 (
            .O(N__5713),
            .I(N__5710));
    Odrv4 I__747 (
            .O(N__5710),
            .I(font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i));
    InMux I__746 (
            .O(N__5707),
            .I(N__5701));
    InMux I__745 (
            .O(N__5706),
            .I(N__5701));
    LocalMux I__744 (
            .O(N__5701),
            .I(beamY_RNI779U3Z0Z_5));
    InMux I__743 (
            .O(N__5698),
            .I(N__5694));
    InMux I__742 (
            .O(N__5697),
            .I(N__5691));
    LocalMux I__741 (
            .O(N__5694),
            .I(N__5683));
    LocalMux I__740 (
            .O(N__5691),
            .I(N__5683));
    InMux I__739 (
            .O(N__5690),
            .I(N__5680));
    InMux I__738 (
            .O(N__5689),
            .I(N__5675));
    InMux I__737 (
            .O(N__5688),
            .I(N__5675));
    Odrv4 I__736 (
            .O(N__5683),
            .I(beamY_RNIUBM4FZ0Z_7));
    LocalMux I__735 (
            .O(N__5680),
            .I(beamY_RNIUBM4FZ0Z_7));
    LocalMux I__734 (
            .O(N__5675),
            .I(beamY_RNIUBM4FZ0Z_7));
    InMux I__733 (
            .O(N__5668),
            .I(N__5662));
    InMux I__732 (
            .O(N__5667),
            .I(N__5662));
    LocalMux I__731 (
            .O(N__5662),
            .I(N__5656));
    InMux I__730 (
            .O(N__5661),
            .I(N__5653));
    InMux I__729 (
            .O(N__5660),
            .I(N__5650));
    InMux I__728 (
            .O(N__5659),
            .I(N__5647));
    Odrv4 I__727 (
            .O(N__5656),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c4));
    LocalMux I__726 (
            .O(N__5653),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c4));
    LocalMux I__725 (
            .O(N__5650),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c4));
    LocalMux I__724 (
            .O(N__5647),
            .I(font_un42_pixel_if_generate_plus_mult1_un61_sum_c4));
    CascadeMux I__723 (
            .O(N__5638),
            .I(N__5634));
    CascadeMux I__722 (
            .O(N__5637),
            .I(N__5629));
    InMux I__721 (
            .O(N__5634),
            .I(N__5624));
    InMux I__720 (
            .O(N__5633),
            .I(N__5624));
    InMux I__719 (
            .O(N__5632),
            .I(N__5619));
    InMux I__718 (
            .O(N__5629),
            .I(N__5619));
    LocalMux I__717 (
            .O(N__5624),
            .I(beamY_RNI9N7M7Z0Z_5));
    LocalMux I__716 (
            .O(N__5619),
            .I(beamY_RNI9N7M7Z0Z_5));
    InMux I__715 (
            .O(N__5614),
            .I(N__5611));
    LocalMux I__714 (
            .O(N__5611),
            .I(beamY_fast_RNIG57D_0Z0Z_4));
    InMux I__713 (
            .O(N__5608),
            .I(N__5605));
    LocalMux I__712 (
            .O(N__5605),
            .I(beamY_fast_RNI45FMZ0Z_7));
    CascadeMux I__711 (
            .O(N__5602),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_));
    InMux I__710 (
            .O(N__5599),
            .I(N__5596));
    LocalMux I__709 (
            .O(N__5596),
            .I(beamY_RNIK0NV_0Z0Z_9));
    InMux I__708 (
            .O(N__5593),
            .I(N__5590));
    LocalMux I__707 (
            .O(N__5590),
            .I(un5_visibley_ac0_11_d));
    CascadeMux I__706 (
            .O(N__5587),
            .I(un5_visibley_c7_cascade_));
    InMux I__705 (
            .O(N__5584),
            .I(N__5581));
    LocalMux I__704 (
            .O(N__5581),
            .I(N__5578));
    Span4Mux_h I__703 (
            .O(N__5578),
            .I(N__5574));
    InMux I__702 (
            .O(N__5577),
            .I(N__5571));
    Odrv4 I__701 (
            .O(N__5574),
            .I(un21_beamy_cry_8_c_RNIOAFZ0Z3));
    LocalMux I__700 (
            .O(N__5571),
            .I(un21_beamy_cry_8_c_RNIOAFZ0Z3));
    InMux I__699 (
            .O(N__5566),
            .I(N__5563));
    LocalMux I__698 (
            .O(N__5563),
            .I(N__5559));
    InMux I__697 (
            .O(N__5562),
            .I(N__5556));
    Span4Mux_h I__696 (
            .O(N__5559),
            .I(N__5551));
    LocalMux I__695 (
            .O(N__5556),
            .I(N__5551));
    Odrv4 I__694 (
            .O(N__5551),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    InMux I__693 (
            .O(N__5548),
            .I(N__5545));
    LocalMux I__692 (
            .O(N__5545),
            .I(N__5541));
    InMux I__691 (
            .O(N__5544),
            .I(N__5538));
    Span4Mux_h I__690 (
            .O(N__5541),
            .I(N__5533));
    LocalMux I__689 (
            .O(N__5538),
            .I(N__5533));
    Odrv4 I__688 (
            .O(N__5533),
            .I(un21_beamy_cry_7_c_RNIM7EZ0Z3));
    InMux I__687 (
            .O(N__5530),
            .I(N__5527));
    LocalMux I__686 (
            .O(N__5527),
            .I(N__5524));
    Odrv4 I__685 (
            .O(N__5524),
            .I(un5_visibley_c5));
    CascadeMux I__684 (
            .O(N__5521),
            .I(N__5518));
    InMux I__683 (
            .O(N__5518),
            .I(N__5515));
    LocalMux I__682 (
            .O(N__5515),
            .I(N__5512));
    Span4Mux_v I__681 (
            .O(N__5512),
            .I(N__5509));
    Odrv4 I__680 (
            .O(N__5509),
            .I(beamY_fastZ0Z_9));
    CascadeMux I__679 (
            .O(N__5506),
            .I(beamY_fast_RNIM4P7_0Z0Z_2_cascade_));
    CascadeMux I__678 (
            .O(N__5503),
            .I(N__5500));
    InMux I__677 (
            .O(N__5500),
            .I(N__5497));
    LocalMux I__676 (
            .O(N__5497),
            .I(N__5494));
    Span4Mux_h I__675 (
            .O(N__5494),
            .I(N__5491));
    Odrv4 I__674 (
            .O(N__5491),
            .I(beamY_fast_RNIO71DZ0Z_3));
    InMux I__673 (
            .O(N__5488),
            .I(N__5479));
    InMux I__672 (
            .O(N__5487),
            .I(N__5474));
    InMux I__671 (
            .O(N__5486),
            .I(N__5474));
    InMux I__670 (
            .O(N__5485),
            .I(N__5471));
    InMux I__669 (
            .O(N__5484),
            .I(N__5464));
    InMux I__668 (
            .O(N__5483),
            .I(N__5464));
    InMux I__667 (
            .O(N__5482),
            .I(N__5464));
    LocalMux I__666 (
            .O(N__5479),
            .I(beamY_fastZ0Z_2));
    LocalMux I__665 (
            .O(N__5474),
            .I(beamY_fastZ0Z_2));
    LocalMux I__664 (
            .O(N__5471),
            .I(beamY_fastZ0Z_2));
    LocalMux I__663 (
            .O(N__5464),
            .I(beamY_fastZ0Z_2));
    CascadeMux I__662 (
            .O(N__5455),
            .I(beamY_fast_RNIM4P7Z0Z_2_cascade_));
    InMux I__661 (
            .O(N__5452),
            .I(N__5446));
    InMux I__660 (
            .O(N__5451),
            .I(N__5440));
    InMux I__659 (
            .O(N__5450),
            .I(N__5435));
    InMux I__658 (
            .O(N__5449),
            .I(N__5435));
    LocalMux I__657 (
            .O(N__5446),
            .I(N__5432));
    InMux I__656 (
            .O(N__5445),
            .I(N__5425));
    InMux I__655 (
            .O(N__5444),
            .I(N__5425));
    InMux I__654 (
            .O(N__5443),
            .I(N__5425));
    LocalMux I__653 (
            .O(N__5440),
            .I(beamY_fastZ0Z_3));
    LocalMux I__652 (
            .O(N__5435),
            .I(beamY_fastZ0Z_3));
    Odrv4 I__651 (
            .O(N__5432),
            .I(beamY_fastZ0Z_3));
    LocalMux I__650 (
            .O(N__5425),
            .I(beamY_fastZ0Z_3));
    InMux I__649 (
            .O(N__5416),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__648 (
            .O(N__5413),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__647 (
            .O(N__5410),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5));
    CascadeMux I__646 (
            .O(N__5407),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    InMux I__645 (
            .O(N__5404),
            .I(N__5401));
    LocalMux I__644 (
            .O(N__5401),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    InMux I__643 (
            .O(N__5398),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__642 (
            .O(N__5395),
            .I(N__5392));
    InMux I__641 (
            .O(N__5392),
            .I(N__5389));
    LocalMux I__640 (
            .O(N__5389),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0));
    InMux I__639 (
            .O(N__5386),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5));
    CascadeMux I__638 (
            .O(N__5383),
            .I(N__5380));
    InMux I__637 (
            .O(N__5380),
            .I(N__5377));
    LocalMux I__636 (
            .O(N__5377),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0));
    InMux I__635 (
            .O(N__5374),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__634 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__633 (
            .O(N__5368),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO));
    InMux I__632 (
            .O(N__5365),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__631 (
            .O(N__5362),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_));
    InMux I__630 (
            .O(N__5359),
            .I(N__5350));
    InMux I__629 (
            .O(N__5358),
            .I(N__5350));
    InMux I__628 (
            .O(N__5357),
            .I(N__5350));
    LocalMux I__627 (
            .O(N__5350),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0));
    InMux I__626 (
            .O(N__5347),
            .I(N__5344));
    LocalMux I__625 (
            .O(N__5344),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8));
    CascadeMux I__624 (
            .O(N__5341),
            .I(N__5338));
    InMux I__623 (
            .O(N__5338),
            .I(N__5335));
    LocalMux I__622 (
            .O(N__5335),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_0));
    InMux I__621 (
            .O(N__5332),
            .I(N__5329));
    LocalMux I__620 (
            .O(N__5329),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf));
    InMux I__619 (
            .O(N__5326),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__618 (
            .O(N__5323),
            .I(N__5320));
    LocalMux I__617 (
            .O(N__5320),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_1));
    InMux I__616 (
            .O(N__5317),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__615 (
            .O(N__5314),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__614 (
            .O(N__5311),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7));
    CascadeMux I__613 (
            .O(N__5308),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_));
    CascadeMux I__612 (
            .O(N__5305),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_));
    InMux I__611 (
            .O(N__5302),
            .I(N__5299));
    LocalMux I__610 (
            .O(N__5299),
            .I(g0_0_2_0));
    CascadeMux I__609 (
            .O(N__5296),
            .I(N__5293));
    InMux I__608 (
            .O(N__5293),
            .I(N__5290));
    LocalMux I__607 (
            .O(N__5290),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf));
    InMux I__606 (
            .O(N__5287),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1));
    InMux I__605 (
            .O(N__5284),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__604 (
            .O(N__5281),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3));
    InMux I__603 (
            .O(N__5278),
            .I(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4));
    CascadeMux I__602 (
            .O(N__5275),
            .I(N__5269));
    InMux I__601 (
            .O(N__5274),
            .I(N__5266));
    InMux I__600 (
            .O(N__5273),
            .I(N__5261));
    InMux I__599 (
            .O(N__5272),
            .I(N__5261));
    InMux I__598 (
            .O(N__5269),
            .I(N__5258));
    LocalMux I__597 (
            .O(N__5266),
            .I(beamXZ0Z_2));
    LocalMux I__596 (
            .O(N__5261),
            .I(beamXZ0Z_2));
    LocalMux I__595 (
            .O(N__5258),
            .I(beamXZ0Z_2));
    InMux I__594 (
            .O(N__5251),
            .I(un5_visiblex_cry_1));
    CascadeMux I__593 (
            .O(N__5248),
            .I(N__5241));
    InMux I__592 (
            .O(N__5247),
            .I(N__5238));
    InMux I__591 (
            .O(N__5246),
            .I(N__5231));
    InMux I__590 (
            .O(N__5245),
            .I(N__5231));
    InMux I__589 (
            .O(N__5244),
            .I(N__5231));
    InMux I__588 (
            .O(N__5241),
            .I(N__5228));
    LocalMux I__587 (
            .O(N__5238),
            .I(beamXZ0Z_3));
    LocalMux I__586 (
            .O(N__5231),
            .I(beamXZ0Z_3));
    LocalMux I__585 (
            .O(N__5228),
            .I(beamXZ0Z_3));
    InMux I__584 (
            .O(N__5221),
            .I(un5_visiblex_cry_2));
    CascadeMux I__583 (
            .O(N__5218),
            .I(N__5211));
    InMux I__582 (
            .O(N__5217),
            .I(N__5208));
    InMux I__581 (
            .O(N__5216),
            .I(N__5205));
    InMux I__580 (
            .O(N__5215),
            .I(N__5200));
    InMux I__579 (
            .O(N__5214),
            .I(N__5200));
    InMux I__578 (
            .O(N__5211),
            .I(N__5197));
    LocalMux I__577 (
            .O(N__5208),
            .I(beamXZ0Z_4));
    LocalMux I__576 (
            .O(N__5205),
            .I(beamXZ0Z_4));
    LocalMux I__575 (
            .O(N__5200),
            .I(beamXZ0Z_4));
    LocalMux I__574 (
            .O(N__5197),
            .I(beamXZ0Z_4));
    InMux I__573 (
            .O(N__5188),
            .I(un5_visiblex_cry_3));
    CascadeMux I__572 (
            .O(N__5185),
            .I(N__5179));
    CascadeMux I__571 (
            .O(N__5184),
            .I(N__5174));
    InMux I__570 (
            .O(N__5183),
            .I(N__5171));
    InMux I__569 (
            .O(N__5182),
            .I(N__5168));
    InMux I__568 (
            .O(N__5179),
            .I(N__5165));
    InMux I__567 (
            .O(N__5178),
            .I(N__5160));
    InMux I__566 (
            .O(N__5177),
            .I(N__5160));
    InMux I__565 (
            .O(N__5174),
            .I(N__5157));
    LocalMux I__564 (
            .O(N__5171),
            .I(beamXZ0Z_5));
    LocalMux I__563 (
            .O(N__5168),
            .I(beamXZ0Z_5));
    LocalMux I__562 (
            .O(N__5165),
            .I(beamXZ0Z_5));
    LocalMux I__561 (
            .O(N__5160),
            .I(beamXZ0Z_5));
    LocalMux I__560 (
            .O(N__5157),
            .I(beamXZ0Z_5));
    InMux I__559 (
            .O(N__5146),
            .I(un5_visiblex_cry_4));
    CascadeMux I__558 (
            .O(N__5143),
            .I(N__5135));
    InMux I__557 (
            .O(N__5142),
            .I(N__5132));
    InMux I__556 (
            .O(N__5141),
            .I(N__5127));
    InMux I__555 (
            .O(N__5140),
            .I(N__5127));
    InMux I__554 (
            .O(N__5139),
            .I(N__5122));
    InMux I__553 (
            .O(N__5138),
            .I(N__5122));
    InMux I__552 (
            .O(N__5135),
            .I(N__5119));
    LocalMux I__551 (
            .O(N__5132),
            .I(beamXZ0Z_6));
    LocalMux I__550 (
            .O(N__5127),
            .I(beamXZ0Z_6));
    LocalMux I__549 (
            .O(N__5122),
            .I(beamXZ0Z_6));
    LocalMux I__548 (
            .O(N__5119),
            .I(beamXZ0Z_6));
    InMux I__547 (
            .O(N__5110),
            .I(un5_visiblex_cry_5));
    InMux I__546 (
            .O(N__5107),
            .I(un5_visiblex_cry_6));
    CascadeMux I__545 (
            .O(N__5104),
            .I(N__5098));
    InMux I__544 (
            .O(N__5103),
            .I(N__5095));
    InMux I__543 (
            .O(N__5102),
            .I(N__5092));
    InMux I__542 (
            .O(N__5101),
            .I(N__5089));
    InMux I__541 (
            .O(N__5098),
            .I(N__5086));
    LocalMux I__540 (
            .O(N__5095),
            .I(beamXZ0Z_8));
    LocalMux I__539 (
            .O(N__5092),
            .I(beamXZ0Z_8));
    LocalMux I__538 (
            .O(N__5089),
            .I(beamXZ0Z_8));
    LocalMux I__537 (
            .O(N__5086),
            .I(beamXZ0Z_8));
    InMux I__536 (
            .O(N__5077),
            .I(bfn_5_10_0_));
    CascadeMux I__535 (
            .O(N__5074),
            .I(N__5070));
    InMux I__534 (
            .O(N__5073),
            .I(N__5066));
    InMux I__533 (
            .O(N__5070),
            .I(N__5063));
    InMux I__532 (
            .O(N__5069),
            .I(N__5059));
    LocalMux I__531 (
            .O(N__5066),
            .I(N__5054));
    LocalMux I__530 (
            .O(N__5063),
            .I(N__5054));
    InMux I__529 (
            .O(N__5062),
            .I(N__5051));
    LocalMux I__528 (
            .O(N__5059),
            .I(beamXZ0Z_9));
    Odrv4 I__527 (
            .O(N__5054),
            .I(beamXZ0Z_9));
    LocalMux I__526 (
            .O(N__5051),
            .I(beamXZ0Z_9));
    InMux I__525 (
            .O(N__5044),
            .I(un5_visiblex_cry_8));
    CascadeMux I__524 (
            .O(N__5041),
            .I(beamY_RNIID28F1_0Z0Z_3_cascade_));
    InMux I__523 (
            .O(N__5038),
            .I(N__5032));
    InMux I__522 (
            .O(N__5037),
            .I(N__5032));
    LocalMux I__521 (
            .O(N__5032),
            .I(un18_beamylt5_0));
    CascadeMux I__520 (
            .O(N__5029),
            .I(un18_beamylto9_2_cascade_));
    InMux I__519 (
            .O(N__5026),
            .I(N__5023));
    LocalMux I__518 (
            .O(N__5023),
            .I(beamY_RNIID28F1Z0Z_3));
    InMux I__517 (
            .O(N__5020),
            .I(N__5015));
    CascadeMux I__516 (
            .O(N__5019),
            .I(N__5012));
    CascadeMux I__515 (
            .O(N__5018),
            .I(N__5007));
    LocalMux I__514 (
            .O(N__5015),
            .I(N__5004));
    InMux I__513 (
            .O(N__5012),
            .I(N__5001));
    InMux I__512 (
            .O(N__5011),
            .I(N__4996));
    InMux I__511 (
            .O(N__5010),
            .I(N__4996));
    InMux I__510 (
            .O(N__5007),
            .I(N__4993));
    Odrv4 I__509 (
            .O(N__5004),
            .I(beamXZ0Z_1));
    LocalMux I__508 (
            .O(N__5001),
            .I(beamXZ0Z_1));
    LocalMux I__507 (
            .O(N__4996),
            .I(beamXZ0Z_1));
    LocalMux I__506 (
            .O(N__4993),
            .I(beamXZ0Z_1));
    InMux I__505 (
            .O(N__4984),
            .I(un5_visiblex_cry_0));
    CascadeMux I__504 (
            .O(N__4981),
            .I(beamY_RNICDD7FZ0Z_5_cascade_));
    InMux I__503 (
            .O(N__4978),
            .I(N__4974));
    InMux I__502 (
            .O(N__4977),
            .I(N__4971));
    LocalMux I__501 (
            .O(N__4974),
            .I(N__4966));
    LocalMux I__500 (
            .O(N__4971),
            .I(N__4966));
    Odrv4 I__499 (
            .O(N__4966),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3));
    CascadeMux I__498 (
            .O(N__4963),
            .I(beamY_RNIUBM4FZ0Z_7_cascade_));
    InMux I__497 (
            .O(N__4960),
            .I(N__4956));
    InMux I__496 (
            .O(N__4959),
            .I(N__4953));
    LocalMux I__495 (
            .O(N__4956),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1));
    LocalMux I__494 (
            .O(N__4953),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1));
    CascadeMux I__493 (
            .O(N__4948),
            .I(N__4945));
    InMux I__492 (
            .O(N__4945),
            .I(N__4942));
    LocalMux I__491 (
            .O(N__4942),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1));
    CascadeMux I__490 (
            .O(N__4939),
            .I(N__4933));
    InMux I__489 (
            .O(N__4938),
            .I(N__4921));
    InMux I__488 (
            .O(N__4937),
            .I(N__4921));
    InMux I__487 (
            .O(N__4936),
            .I(N__4921));
    InMux I__486 (
            .O(N__4933),
            .I(N__4921));
    InMux I__485 (
            .O(N__4932),
            .I(N__4921));
    LocalMux I__484 (
            .O(N__4921),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_c5));
    CascadeMux I__483 (
            .O(N__4918),
            .I(N__4914));
    CascadeMux I__482 (
            .O(N__4917),
            .I(N__4910));
    InMux I__481 (
            .O(N__4914),
            .I(N__4900));
    InMux I__480 (
            .O(N__4913),
            .I(N__4900));
    InMux I__479 (
            .O(N__4910),
            .I(N__4900));
    InMux I__478 (
            .O(N__4909),
            .I(N__4900));
    LocalMux I__477 (
            .O(N__4900),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i));
    CascadeMux I__476 (
            .O(N__4897),
            .I(N__4894));
    InMux I__475 (
            .O(N__4894),
            .I(N__4891));
    LocalMux I__474 (
            .O(N__4891),
            .I(beamY_fastZ0Z_8));
    InMux I__473 (
            .O(N__4888),
            .I(N__4883));
    InMux I__472 (
            .O(N__4887),
            .I(N__4878));
    InMux I__471 (
            .O(N__4886),
            .I(N__4878));
    LocalMux I__470 (
            .O(N__4883),
            .I(beamY_fastZ0Z_4));
    LocalMux I__469 (
            .O(N__4878),
            .I(beamY_fastZ0Z_4));
    CascadeMux I__468 (
            .O(N__4873),
            .I(beamY_fast_RNI24GAZ0Z_2_cascade_));
    CascadeMux I__467 (
            .O(N__4870),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cascade_));
    InMux I__466 (
            .O(N__4867),
            .I(N__4864));
    LocalMux I__465 (
            .O(N__4864),
            .I(beamY_RNI2GUN3Z0Z_9));
    CascadeMux I__464 (
            .O(N__4861),
            .I(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_));
    InMux I__463 (
            .O(N__4858),
            .I(N__4855));
    LocalMux I__462 (
            .O(N__4855),
            .I(beamY_RNI2GUN3_0Z0Z_9));
    InMux I__461 (
            .O(N__4852),
            .I(N__4849));
    LocalMux I__460 (
            .O(N__4849),
            .I(d_i4_mux));
    CascadeMux I__459 (
            .O(N__4846),
            .I(beamY_fast_RNIG57DZ0Z_4_cascade_));
    CascadeMux I__458 (
            .O(N__4843),
            .I(un5_visibley_c5_cascade_));
    InMux I__457 (
            .O(N__4840),
            .I(N__4836));
    InMux I__456 (
            .O(N__4839),
            .I(N__4833));
    LocalMux I__455 (
            .O(N__4836),
            .I(N__4830));
    LocalMux I__454 (
            .O(N__4833),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    Odrv12 I__453 (
            .O(N__4830),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    InMux I__452 (
            .O(N__4825),
            .I(N__4819));
    InMux I__451 (
            .O(N__4824),
            .I(N__4819));
    LocalMux I__450 (
            .O(N__4819),
            .I(un21_beamy_cry_3_c_RNIERZ0Z93));
    InMux I__449 (
            .O(N__4816),
            .I(N__4813));
    LocalMux I__448 (
            .O(N__4813),
            .I(N__4809));
    InMux I__447 (
            .O(N__4812),
            .I(N__4806));
    Odrv4 I__446 (
            .O(N__4809),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    LocalMux I__445 (
            .O(N__4806),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    CascadeMux I__444 (
            .O(N__4801),
            .I(un5_visibley_ac0_11_d_cascade_));
    CascadeMux I__443 (
            .O(N__4798),
            .I(N_7_1_cascade_));
    CascadeMux I__442 (
            .O(N__4795),
            .I(N__4792));
    InMux I__441 (
            .O(N__4792),
            .I(N__4789));
    LocalMux I__440 (
            .O(N__4789),
            .I(g2_1_0));
    CascadeMux I__439 (
            .O(N__4786),
            .I(N_14_cascade_));
    InMux I__438 (
            .O(N__4783),
            .I(un8_beamx_cry_1));
    InMux I__437 (
            .O(N__4780),
            .I(un8_beamx_cry_2));
    InMux I__436 (
            .O(N__4777),
            .I(un8_beamx_cry_3));
    InMux I__435 (
            .O(N__4774),
            .I(un8_beamx_cry_4));
    InMux I__434 (
            .O(N__4771),
            .I(un8_beamx_cry_5));
    InMux I__433 (
            .O(N__4768),
            .I(un8_beamx_cry_6));
    InMux I__432 (
            .O(N__4765),
            .I(un8_beamx_cry_7));
    InMux I__431 (
            .O(N__4762),
            .I(bfn_4_10_0_));
    InMux I__430 (
            .O(N__4759),
            .I(un8_beamx_cry_9));
    CascadeMux I__429 (
            .O(N__4756),
            .I(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_));
    CascadeMux I__428 (
            .O(N__4753),
            .I(un3_beamx_5_cascade_));
    CascadeMux I__427 (
            .O(N__4750),
            .I(un3_beamx_7_cascade_));
    CascadeMux I__426 (
            .O(N__4747),
            .I(beamX_RNI5457Z0Z_5_cascade_));
    CascadeMux I__425 (
            .O(N__4744),
            .I(un13_beamylto2_0_cascade_));
    InMux I__424 (
            .O(N__4741),
            .I(N__4738));
    LocalMux I__423 (
            .O(N__4738),
            .I(un5_beamx_3));
    CascadeMux I__422 (
            .O(N__4735),
            .I(un5_beamx_4_cascade_));
    InMux I__421 (
            .O(N__4732),
            .I(N__4729));
    LocalMux I__420 (
            .O(N__4729),
            .I(beamY_RNIMA24P1Z0Z_5));
    InMux I__419 (
            .O(N__4726),
            .I(un21_beamy_cry_2));
    InMux I__418 (
            .O(N__4723),
            .I(un21_beamy_cry_3));
    InMux I__417 (
            .O(N__4720),
            .I(un21_beamy_cry_4));
    InMux I__416 (
            .O(N__4717),
            .I(un21_beamy_cry_5));
    InMux I__415 (
            .O(N__4714),
            .I(un21_beamy_cry_6));
    InMux I__414 (
            .O(N__4711),
            .I(un21_beamy_cry_7));
    InMux I__413 (
            .O(N__4708),
            .I(bfn_4_4_0_));
    IoInMux I__412 (
            .O(N__4705),
            .I(N__4702));
    LocalMux I__411 (
            .O(N__4702),
            .I(N__4699));
    IoSpan4Mux I__410 (
            .O(N__4699),
            .I(N__4696));
    IoSpan4Mux I__409 (
            .O(N__4696),
            .I(N__4693));
    IoSpan4Mux I__408 (
            .O(N__4693),
            .I(N__4690));
    Odrv4 I__407 (
            .O(N__4690),
            .I(\Clock50MHz.PixelClock ));
    IoInMux I__406 (
            .O(N__4687),
            .I(N__4684));
    LocalMux I__405 (
            .O(N__4684),
            .I(N__4681));
    IoSpan4Mux I__404 (
            .O(N__4681),
            .I(N__4678));
    Odrv4 I__403 (
            .O(N__4678),
            .I(Clock12MHz_c));
    InMux I__402 (
            .O(N__4675),
            .I(un21_beamy_cry_1));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__4705),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_4_3_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_4_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(N__10367),
            .in2(N__10190),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_RNIAL73_LC_4_3_1.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_4_3_1.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_4_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_1_c_RNIAL73_LC_4_3_1 (
            .in0(_gnd_net_),
            .in1(N__8990),
            .in2(_gnd_net_),
            .in3(N__4675),
            .lcout(un21_beamy_cry_1_c_RNIALZ0Z73),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_2_c_RNICO83_LC_4_3_2.C_ON=1'b1;
    defparam un21_beamy_cry_2_c_RNICO83_LC_4_3_2.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_2_c_RNICO83_LC_4_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_2_c_RNICO83_LC_4_3_2 (
            .in0(_gnd_net_),
            .in1(N__8046),
            .in2(_gnd_net_),
            .in3(N__4726),
            .lcout(un21_beamy_cry_2_c_RNICOZ0Z83),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_3_c_RNIER93_LC_4_3_3.C_ON=1'b1;
    defparam un21_beamy_cry_3_c_RNIER93_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_3_c_RNIER93_LC_4_3_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_3_c_RNIER93_LC_4_3_3 (
            .in0(_gnd_net_),
            .in1(N__7938),
            .in2(_gnd_net_),
            .in3(N__4723),
            .lcout(un21_beamy_cry_3_c_RNIERZ0Z93),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_4_3_4.C_ON=1'b1;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_4_3_4.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_4_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_4_c_RNIGUA3_LC_4_3_4 (
            .in0(_gnd_net_),
            .in1(N__8901),
            .in2(_gnd_net_),
            .in3(N__4720),
            .lcout(un21_beamy_cry_4_c_RNIGUAZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_5_c_RNII1C3_LC_4_3_5.C_ON=1'b1;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_4_3_5.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_5_c_RNII1C3_LC_4_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_5_c_RNII1C3_LC_4_3_5 (
            .in0(_gnd_net_),
            .in1(N__8838),
            .in2(_gnd_net_),
            .in3(N__4717),
            .lcout(un21_beamy_cry_5_c_RNII1CZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_4_3_6.C_ON=1'b1;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_4_3_6.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_4_3_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_6_c_RNIK4D3_LC_4_3_6 (
            .in0(_gnd_net_),
            .in1(N__8763),
            .in2(_gnd_net_),
            .in3(N__4714),
            .lcout(un21_beamy_cry_6_c_RNIK4DZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_4_3_7.C_ON=1'b1;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_4_3_7.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_7_c_RNIM7E3_LC_4_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_7_c_RNIM7E3_LC_4_3_7 (
            .in0(_gnd_net_),
            .in1(N__7881),
            .in2(_gnd_net_),
            .in3(N__4711),
            .lcout(un21_beamy_cry_7_c_RNIM7EZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_4_4_0.C_ON=1'b0;
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_4_4_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_8_c_RNIOAF3_LC_4_4_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 un21_beamy_cry_8_c_RNIOAF3_LC_4_4_0 (
            .in0(_gnd_net_),
            .in1(N__7810),
            .in2(_gnd_net_),
            .in3(N__4708),
            .lcout(un21_beamy_cry_8_c_RNIOAFZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_4_4_1.C_ON=1'b0;
    defparam beamY_0_LC_4_4_1.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_4_4_1.LUT_INIT=16'b0011001101000100;
    LogicCell40 beamY_0_LC_4_4_1 (
            .in0(N__8157),
            .in1(N__8249),
            .in2(_gnd_net_),
            .in3(N__10133),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9818),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_5_LC_4_4_3.C_ON=1'b0;
    defparam beamY_RNI6125_5_LC_4_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_5_LC_4_4_3.LUT_INIT=16'b1001001100110011;
    LogicCell40 beamY_RNI6125_5_LC_4_4_3 (
            .in0(N__8945),
            .in1(N__8889),
            .in2(N__8019),
            .in3(N__7932),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_3_LC_4_5_1.C_ON=1'b0;
    defparam beamY_3_LC_4_5_1.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_4_5_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_3_LC_4_5_1 (
            .in0(N__8131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4840),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9817),
            .ce(N__8248),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_4_5_2.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_4_5_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_3_LC_4_5_2 (
            .in0(_gnd_net_),
            .in1(N__8017),
            .in2(_gnd_net_),
            .in3(N__8992),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_9_LC_4_5_4.C_ON=1'b0;
    defparam beamY_fast_9_LC_4_5_4.SEQ_MODE=4'b1000;
    defparam beamY_fast_9_LC_4_5_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 beamY_fast_9_LC_4_5_4 (
            .in0(_gnd_net_),
            .in1(N__8133),
            .in2(_gnd_net_),
            .in3(N__5577),
            .lcout(beamY_fastZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9817),
            .ce(N__8248),
            .sr(_gnd_net_));
    defparam beamY_7_LC_4_5_5.C_ON=1'b0;
    defparam beamY_7_LC_4_5_5.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_4_5_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_7_LC_4_5_5 (
            .in0(N__8132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5562),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9817),
            .ce(N__8248),
            .sr(_gnd_net_));
    defparam beamY_RNIC725_9_LC_4_6_1.C_ON=1'b0;
    defparam beamY_RNIC725_9_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIC725_9_LC_4_6_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamY_RNIC725_9_LC_4_6_1 (
            .in0(N__8018),
            .in1(N__7805),
            .in2(N__10369),
            .in3(N__8750),
            .lcout(un5_beamx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5025_5_LC_4_6_3.C_ON=1'b0;
    defparam beamY_RNI5025_5_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI5025_5_LC_4_6_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamY_RNI5025_5_LC_4_6_3 (
            .in0(N__8993),
            .in1(N__8847),
            .in2(N__10175),
            .in3(N__8920),
            .lcout(),
            .ltout(un5_beamx_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_8_LC_4_6_4.C_ON=1'b0;
    defparam beamY_RNI9DLC_8_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_8_LC_4_6_4.LUT_INIT=16'b0000000010000000;
    LogicCell40 beamY_RNI9DLC_8_LC_4_6_4 (
            .in0(N__4741),
            .in1(N__7951),
            .in2(N__4735),
            .in3(N__7882),
            .lcout(un5_beamx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMA24P1_5_LC_4_7_2.C_ON=1'b0;
    defparam beamY_RNIMA24P1_5_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIMA24P1_5_LC_4_7_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIMA24P1_5_LC_4_7_2 (
            .in0(N__5690),
            .in1(N__5660),
            .in2(N__4948),
            .in3(N__7509),
            .lcout(beamY_RNIMA24P1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMM6891_5_LC_4_7_6.C_ON=1'b0;
    defparam beamY_RNIMM6891_5_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIMM6891_5_LC_4_7_6.LUT_INIT=16'b0101011001011010;
    LogicCell40 beamY_RNIMM6891_5_LC_4_7_6 (
            .in0(N__4959),
            .in1(N__6646),
            .in2(N__5740),
            .in3(N__7510),
            .lcout(),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPFUEA4_3_LC_4_7_7.C_ON=1'b0;
    defparam beamY_RNIPFUEA4_3_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIPFUEA4_3_LC_4_7_7.LUT_INIT=16'b1100001101000001;
    LogicCell40 beamY_RNIPFUEA4_3_LC_4_7_7 (
            .in0(N__4732),
            .in1(N__5919),
            .in2(N__4756),
            .in3(N__8033),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI6PL_3_LC_4_8_0.C_ON=1'b0;
    defparam beamX_RNI6PL_3_LC_4_8_0.SEQ_MODE=4'b0000;
    defparam beamX_RNI6PL_3_LC_4_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNI6PL_3_LC_4_8_0 (
            .in0(N__5245),
            .in1(N__5215),
            .in2(N__5185),
            .in3(N__5140),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_4_8_1.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_4_8_1.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_RNIR4B_9_LC_4_8_1 (
            .in0(_gnd_net_),
            .in1(N__5073),
            .in2(_gnd_net_),
            .in3(N__5102),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_10_LC_4_8_2.C_ON=1'b0;
    defparam beamX_RNICPU5_10_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_10_LC_4_8_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNICPU5_10_LC_4_8_2 (
            .in0(N__5216),
            .in1(N__5273),
            .in2(N__8637),
            .in3(N__5011),
            .lcout(),
            .ltout(un3_beamx_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_3_LC_4_8_3.C_ON=1'b0;
    defparam beamX_RNIKVE6_3_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_3_LC_4_8_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNIKVE6_3_LC_4_8_3 (
            .in0(N__5141),
            .in1(N__5246),
            .in2(N__4753),
            .in3(N__10635),
            .lcout(),
            .ltout(un3_beamx_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_4_8_4.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_4_8_4.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNI5457_5_LC_4_8_4 (
            .in0(N__8581),
            .in1(N__6910),
            .in2(N__4750),
            .in3(N__5182),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(beamX_RNI5457Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_4_8_5.C_ON=1'b0;
    defparam beamX_0_LC_4_8_5.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_4_8_5.LUT_INIT=16'b0000000000001111;
    LogicCell40 beamX_0_LC_4_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4747),
            .in3(N__10636),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9814),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIDMA_1_LC_4_8_6.C_ON=1'b0;
    defparam beamX_RNIDMA_1_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam beamX_RNIDMA_1_LC_4_8_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamX_RNIDMA_1_LC_4_8_6 (
            .in0(_gnd_net_),
            .in1(N__5272),
            .in2(_gnd_net_),
            .in3(N__5010),
            .lcout(),
            .ltout(un13_beamylto2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIJQQ_3_LC_4_8_7.C_ON=1'b0;
    defparam beamX_RNIJQQ_3_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIJQQ_3_LC_4_8_7.LUT_INIT=16'b1010100010001000;
    LogicCell40 beamX_RNIJQQ_3_LC_4_8_7 (
            .in0(N__5214),
            .in1(N__5244),
            .in2(N__4744),
            .in3(N__10634),
            .lcout(un18_beamylt5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_4_9_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_4_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_4_9_0 (
            .in0(_gnd_net_),
            .in1(N__10648),
            .in2(N__5019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_4_9_1.C_ON=1'b1;
    defparam beamX_2_LC_4_9_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_4_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(N__5274),
            .in2(_gnd_net_),
            .in3(N__4783),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_4_9_2.C_ON=1'b1;
    defparam beamX_3_LC_4_9_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_4_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(N__5247),
            .in2(_gnd_net_),
            .in3(N__4780),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_4_9_3.C_ON=1'b1;
    defparam beamX_4_LC_4_9_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_4_9_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_4_9_3 (
            .in0(N__8195),
            .in1(N__5217),
            .in2(_gnd_net_),
            .in3(N__4777),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_4_9_4.C_ON=1'b1;
    defparam beamX_5_LC_4_9_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_4_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_4_9_4 (
            .in0(_gnd_net_),
            .in1(N__5183),
            .in2(_gnd_net_),
            .in3(N__4774),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_4_9_5.C_ON=1'b1;
    defparam beamX_6_LC_4_9_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_4_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_4_9_5 (
            .in0(_gnd_net_),
            .in1(N__5142),
            .in2(_gnd_net_),
            .in3(N__4771),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_4_9_6.C_ON=1'b1;
    defparam beamX_7_LC_4_9_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_4_9_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_4_9_6 (
            .in0(_gnd_net_),
            .in1(N__6911),
            .in2(_gnd_net_),
            .in3(N__4768),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_4_9_7.C_ON=1'b1;
    defparam beamX_8_LC_4_9_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_4_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_4_9_7 (
            .in0(_gnd_net_),
            .in1(N__5103),
            .in2(_gnd_net_),
            .in3(N__4765),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__9812),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_4_10_0.C_ON=1'b1;
    defparam beamX_9_LC_4_10_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_4_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_4_10_0 (
            .in0(_gnd_net_),
            .in1(N__5069),
            .in2(_gnd_net_),
            .in3(N__4762),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__9813),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_4_10_1.C_ON=1'b0;
    defparam beamX_10_LC_4_10_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_4_10_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_4_10_1 (
            .in0(N__8623),
            .in1(N__8203),
            .in2(_gnd_net_),
            .in3(N__4759),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9813),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_66_LC_4_10_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_66_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_66_LC_4_10_2.LUT_INIT=16'b0001000111001110;
    LogicCell40 Pixel_1_esr_RNO_66_LC_4_10_2 (
            .in0(N__10810),
            .in1(N__9725),
            .in2(N__4795),
            .in3(N__9638),
            .lcout(),
            .ltout(N_7_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_51_LC_4_10_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_51_LC_4_10_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_51_LC_4_10_3.LUT_INIT=16'b0000111111111111;
    LogicCell40 Pixel_1_esr_RNO_51_LC_4_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4798),
            .in3(N__5302),
            .lcout(g0_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_70_LC_4_10_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_70_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_70_LC_4_10_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 Pixel_1_esr_RNO_70_LC_4_10_5 (
            .in0(_gnd_net_),
            .in1(N__10492),
            .in2(_gnd_net_),
            .in3(N__11074),
            .lcout(g2_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_53_LC_4_11_0.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_53_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_53_LC_4_11_0.LUT_INIT=16'b0101010101110111;
    LogicCell40 Pixel_1_esr_RNO_53_LC_4_11_0 (
            .in0(N__10820),
            .in1(N__10572),
            .in2(_gnd_net_),
            .in3(N__11096),
            .lcout(),
            .ltout(N_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_30_LC_4_11_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_30_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_30_LC_4_11_1.LUT_INIT=16'b0000000001010000;
    LogicCell40 Pixel_1_esr_RNO_30_LC_4_11_1 (
            .in0(N__9648),
            .in1(_gnd_net_),
            .in2(N__4786),
            .in3(N__9759),
            .lcout(G_25_i_a8_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_12_1.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_12_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_4_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_4_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9647),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_5_3_2.C_ON=1'b0;
    defparam beamY_2_LC_5_3_2.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_5_3_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 beamY_2_LC_5_3_2 (
            .in0(_gnd_net_),
            .in1(N__4812),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(N__8241),
            .sr(_gnd_net_));
    defparam beamY_5_LC_5_3_4.C_ON=1'b0;
    defparam beamY_5_LC_5_3_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_5_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_5_LC_5_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6780),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(N__8241),
            .sr(_gnd_net_));
    defparam beamY_6_LC_5_3_7.C_ON=1'b0;
    defparam beamY_6_LC_5_3_7.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_5_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_6_LC_5_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6831),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(N__8241),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIG57D_4_LC_5_4_0.C_ON=1'b0;
    defparam beamY_fast_RNIG57D_4_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIG57D_4_LC_5_4_0.LUT_INIT=16'b1111111011111010;
    LogicCell40 beamY_fast_RNIG57D_4_LC_5_4_0 (
            .in0(N__6768),
            .in1(N__4888),
            .in2(N__8828),
            .in3(N__5488),
            .lcout(),
            .ltout(beamY_fast_RNIG57DZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIQQEM_5_LC_5_4_1.C_ON=1'b0;
    defparam beamY_fast_RNIQQEM_5_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIQQEM_5_LC_5_4_1.LUT_INIT=16'b1111000011101110;
    LogicCell40 beamY_fast_RNIQQEM_5_LC_5_4_1 (
            .in0(N__8812),
            .in1(N__6769),
            .in2(N__4846),
            .in3(N__5451),
            .lcout(un5_visibley_c5),
            .ltout(un5_visibley_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIK3TH2_7_LC_5_4_2.C_ON=1'b0;
    defparam beamY_RNIK3TH2_7_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIK3TH2_7_LC_5_4_2.LUT_INIT=16'b0110100100010010;
    LogicCell40 beamY_RNIK3TH2_7_LC_5_4_2 (
            .in0(N__8741),
            .in1(N__6733),
            .in2(N__4843),
            .in3(N__6684),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_4_LC_5_4_3.C_ON=1'b0;
    defparam beamY_fast_4_LC_5_4_3.SEQ_MODE=4'b1000;
    defparam beamY_fast_4_LC_5_4_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_fast_4_LC_5_4_3 (
            .in0(N__4825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8156),
            .lcout(beamY_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9822),
            .ce(N__8224),
            .sr(_gnd_net_));
    defparam beamY_fast_3_LC_5_4_6.C_ON=1'b0;
    defparam beamY_fast_3_LC_5_4_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_3_LC_5_4_6.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_fast_3_LC_5_4_6 (
            .in0(N__8155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4839),
            .lcout(beamY_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9822),
            .ce(N__8224),
            .sr(_gnd_net_));
    defparam beamY_4_LC_5_4_7.C_ON=1'b0;
    defparam beamY_4_LC_5_4_7.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_5_4_7.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_4_LC_5_4_7 (
            .in0(N__4824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8154),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9822),
            .ce(N__8224),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIBVU7_2_LC_5_5_1.C_ON=1'b0;
    defparam beamY_fast_RNIBVU7_2_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIBVU7_2_LC_5_5_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_fast_RNIBVU7_2_LC_5_5_1 (
            .in0(_gnd_net_),
            .in1(N__5445),
            .in2(_gnd_net_),
            .in3(N__5484),
            .lcout(un5_visibley_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_2_LC_5_5_2.C_ON=1'b0;
    defparam beamY_fast_2_LC_5_5_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_2_LC_5_5_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_fast_2_LC_5_5_2 (
            .in0(N__4816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9819),
            .ce(N__8228),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIT5UF_8_LC_5_5_3.C_ON=1'b0;
    defparam beamY_fast_RNIT5UF_8_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIT5UF_8_LC_5_5_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_fast_RNIT5UF_8_LC_5_5_3 (
            .in0(N__4886),
            .in1(N__5443),
            .in2(N__4897),
            .in3(N__5482),
            .lcout(un5_visibley_ac0_11_d),
            .ltout(un5_visibley_ac0_11_d_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI45FM_7_LC_5_5_4.C_ON=1'b0;
    defparam beamY_fast_RNI45FM_7_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI45FM_7_LC_5_5_4.LUT_INIT=16'b1100110011001001;
    LogicCell40 beamY_fast_RNI45FM_7_LC_5_5_4 (
            .in0(N__6488),
            .in1(N__7785),
            .in2(N__4801),
            .in3(N__7849),
            .lcout(beamY_fast_RNI45FMZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_8_LC_5_5_6.C_ON=1'b0;
    defparam beamY_fast_8_LC_5_5_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_8_LC_5_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_8_LC_5_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5544),
            .lcout(beamY_fastZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9819),
            .ce(N__8228),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIG57D_0_4_LC_5_5_7.C_ON=1'b0;
    defparam beamY_fast_RNIG57D_0_4_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIG57D_0_4_LC_5_5_7.LUT_INIT=16'b1000011100001111;
    LogicCell40 beamY_fast_RNIG57D_0_4_LC_5_5_7 (
            .in0(N__4887),
            .in1(N__5444),
            .in2(N__7869),
            .in3(N__5483),
            .lcout(beamY_fast_RNIG57D_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI24GA_2_LC_5_6_0.C_ON=1'b0;
    defparam beamY_fast_RNI24GA_2_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI24GA_2_LC_5_6_0.LUT_INIT=16'b1000011100001111;
    LogicCell40 beamY_fast_RNI24GA_2_LC_5_6_0 (
            .in0(N__7939),
            .in1(N__5452),
            .in2(N__8751),
            .in3(N__5485),
            .lcout(),
            .ltout(beamY_fast_RNI24GAZ0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGTNJ_7_LC_5_6_1.C_ON=1'b0;
    defparam beamY_RNIGTNJ_7_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIGTNJ_7_LC_5_6_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 beamY_RNIGTNJ_7_LC_5_6_1 (
            .in0(_gnd_net_),
            .in1(N__8737),
            .in2(N__4873),
            .in3(N__6802),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum),
            .ltout(un1_beamY_if_generate_plus_mult1_un40_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2GUN3_9_LC_5_6_2.C_ON=1'b0;
    defparam beamY_RNI2GUN3_9_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2GUN3_9_LC_5_6_2.LUT_INIT=16'b1001001000010110;
    LogicCell40 beamY_RNI2GUN3_9_LC_5_6_2 (
            .in0(N__8461),
            .in1(N__5757),
            .in2(N__4870),
            .in3(N__8406),
            .lcout(beamY_RNI2GUN3Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIO3Q1A_7_LC_5_6_3.C_ON=1'b0;
    defparam beamY_RNIO3Q1A_7_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIO3Q1A_7_LC_5_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 beamY_RNIO3Q1A_7_LC_5_6_3 (
            .in0(N__4977),
            .in1(N__4858),
            .in2(_gnd_net_),
            .in3(N__4867),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un54_sum_axbxc5_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNITVFT2_3_LC_5_6_4.C_ON=1'b0;
    defparam beamY_fast_RNITVFT2_3_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNITVFT2_3_LC_5_6_4.LUT_INIT=16'b0000011000000100;
    LogicCell40 beamY_fast_RNITVFT2_3_LC_5_6_4 (
            .in0(N__8333),
            .in1(N__8454),
            .in2(N__5503),
            .in3(N__6685),
            .lcout(),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_7_0_i4_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI47PR6_8_LC_5_6_5.C_ON=1'b0;
    defparam beamY_RNI47PR6_8_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI47PR6_8_LC_5_6_5.LUT_INIT=16'b0011101011001010;
    LogicCell40 beamY_RNI47PR6_8_LC_5_6_5 (
            .in0(N__4852),
            .in1(N__6691),
            .in2(N__4861),
            .in3(N__6734),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un54_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2GUN3_0_9_LC_5_6_6.C_ON=1'b0;
    defparam beamY_RNI2GUN3_0_9_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI2GUN3_0_9_LC_5_6_6.LUT_INIT=16'b0110110111101001;
    LogicCell40 beamY_RNI2GUN3_0_9_LC_5_6_6 (
            .in0(N__8332),
            .in1(N__5758),
            .in2(N__8474),
            .in3(N__8407),
            .lcout(beamY_RNI2GUN3_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIAI342_9_LC_5_6_7.C_ON=1'b0;
    defparam beamY_fast_RNIAI342_9_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIAI342_9_LC_5_6_7.LUT_INIT=16'b0101100010000101;
    LogicCell40 beamY_fast_RNIAI342_9_LC_5_6_7 (
            .in0(N__8408),
            .in1(N__7498),
            .in2(N__8469),
            .in3(N__8331),
            .lcout(d_i4_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDRE6H_0_3_LC_5_7_0.C_ON=1'b0;
    defparam beamY_RNIDRE6H_0_3_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIDRE6H_0_3_LC_5_7_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIDRE6H_0_3_LC_5_7_0 (
            .in0(N__7507),
            .in1(N__7653),
            .in2(N__4918),
            .in3(N__4938),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICDD7F_5_LC_5_7_1.C_ON=1'b0;
    defparam beamY_RNICDD7F_5_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNICDD7F_5_LC_5_7_1.LUT_INIT=16'b1110111010101010;
    LogicCell40 beamY_RNICDD7F_5_LC_5_7_1 (
            .in0(N__5733),
            .in1(N__6645),
            .in2(_gnd_net_),
            .in3(N__7508),
            .lcout(),
            .ltout(beamY_RNICDD7FZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRJ4CH2_3_LC_5_7_2.C_ON=1'b0;
    defparam beamY_RNIRJ4CH2_3_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIRJ4CH2_3_LC_5_7_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 beamY_RNIRJ4CH2_3_LC_5_7_2 (
            .in0(N__7981),
            .in1(N__4960),
            .in2(N__4981),
            .in3(N__5920),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUBM4F_7_LC_5_7_3.C_ON=1'b0;
    defparam beamY_RNIUBM4F_7_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIUBM4F_7_LC_5_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIUBM4F_7_LC_5_7_3 (
            .in0(N__4978),
            .in1(N__8281),
            .in2(N__4939),
            .in3(N__6999),
            .lcout(beamY_RNIUBM4FZ0Z_7),
            .ltout(beamY_RNIUBM4FZ0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKUC181_5_LC_5_7_4.C_ON=1'b0;
    defparam beamY_RNIKUC181_5_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIKUC181_5_LC_5_7_4.LUT_INIT=16'b0110111100000110;
    LogicCell40 beamY_RNIKUC181_5_LC_5_7_4 (
            .in0(N__7002),
            .in1(N__5707),
            .in2(N__4963),
            .in3(N__5659),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un61_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIA9P0Q_4_LC_5_7_5.C_ON=1'b0;
    defparam beamY_RNIA9P0Q_4_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIA9P0Q_4_LC_5_7_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIA9P0Q_4_LC_5_7_5 (
            .in0(N__4937),
            .in1(N__4913),
            .in2(N__6622),
            .in3(N__7001),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI52RJO_5_LC_5_7_6.C_ON=1'b0;
    defparam beamY_RNI52RJO_5_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI52RJO_5_LC_5_7_6.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNI52RJO_5_LC_5_7_6 (
            .in0(N__7000),
            .in1(N__5706),
            .in2(N__4917),
            .in3(N__4936),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5_m3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDRE6H_3_LC_5_7_7.C_ON=1'b0;
    defparam beamY_RNIDRE6H_3_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIDRE6H_3_LC_5_7_7.LUT_INIT=16'b1001000011111001;
    LogicCell40 beamY_RNIDRE6H_3_LC_5_7_7 (
            .in0(N__4932),
            .in1(N__4909),
            .in2(N__7667),
            .in3(N__7506),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un61_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICIBSR6_2_LC_5_8_0.C_ON=1'b0;
    defparam beamY_RNICIBSR6_2_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam beamY_RNICIBSR6_2_LC_5_8_0.LUT_INIT=16'b0001000111101110;
    LogicCell40 beamY_RNICIBSR6_2_LC_5_8_0 (
            .in0(N__5835),
            .in1(N__5814),
            .in2(_gnd_net_),
            .in3(N__8991),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un1_sum_axb2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIID28F1_0_3_LC_5_8_1.C_ON=1'b0;
    defparam beamY_RNIID28F1_0_3_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIID28F1_0_3_LC_5_8_1.LUT_INIT=16'b0101101001101001;
    LogicCell40 beamY_RNIID28F1_0_3_LC_5_8_1 (
            .in0(N__5893),
            .in1(N__5632),
            .in2(N__7677),
            .in3(N__5688),
            .lcout(),
            .ltout(beamY_RNIID28F1_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHMJMF3_3_LC_5_8_2.C_ON=1'b0;
    defparam beamY_RNIHMJMF3_3_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIHMJMF3_3_LC_5_8_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNIHMJMF3_3_LC_5_8_2 (
            .in0(_gnd_net_),
            .in1(N__5661),
            .in2(N__5041),
            .in3(N__5026),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un68_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI4AB1_5_LC_5_8_3.C_ON=1'b0;
    defparam beamX_RNI4AB1_5_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam beamX_RNI4AB1_5_LC_5_8_3.LUT_INIT=16'b1110000010100000;
    LogicCell40 beamX_RNI4AB1_5_LC_5_8_3 (
            .in0(N__5139),
            .in1(N__5178),
            .in2(N__6912),
            .in3(N__5038),
            .lcout(un13_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNII5M_9_LC_5_8_4.C_ON=1'b0;
    defparam beamX_RNII5M_9_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam beamX_RNII5M_9_LC_5_8_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNII5M_9_LC_5_8_4 (
            .in0(N__5101),
            .in1(N__6903),
            .in2(N__5074),
            .in3(N__5138),
            .lcout(),
            .ltout(un18_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_5_LC_5_8_5.C_ON=1'b0;
    defparam beamX_RNIVEM1_5_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_5_LC_5_8_5.LUT_INIT=16'b1111000011000000;
    LogicCell40 beamX_RNIVEM1_5_LC_5_8_5 (
            .in0(_gnd_net_),
            .in1(N__5037),
            .in2(N__5029),
            .in3(N__5177),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIID28F1_3_LC_5_8_6.C_ON=1'b0;
    defparam beamY_RNIID28F1_3_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIID28F1_3_LC_5_8_6.LUT_INIT=16'b1001001101101100;
    LogicCell40 beamY_RNIID28F1_3_LC_5_8_6 (
            .in0(N__5689),
            .in1(N__7668),
            .in2(N__5637),
            .in3(N__5892),
            .lcout(beamY_RNIID28F1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_5_8_7.C_ON=1'b0;
    defparam beamX_1_LC_5_8_7.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_5_8_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_5_8_7 (
            .in0(_gnd_net_),
            .in1(N__5020),
            .in2(_gnd_net_),
            .in3(N__10649),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9815),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_5_9_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_5_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10650),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_5_9_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_5_9_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5018),
            .in3(N__4984),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_5_9_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_5_9_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5275),
            .in3(N__5251),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_5_9_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_5_9_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_5_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_5_9_3 (
            .in0(_gnd_net_),
            .in1(N__9075),
            .in2(N__5248),
            .in3(N__5221),
            .lcout(un1_visiblex_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_5_9_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_5_9_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_5_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5218),
            .in3(N__5188),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_5_9_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_5_9_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_5_9_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_5_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5184),
            .in3(N__5146),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_5_9_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_5_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(N__9076),
            .in2(N__5143),
            .in3(N__5110),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_5_9_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_5_9_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_5_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_5_9_7 (
            .in0(_gnd_net_),
            .in1(N__6902),
            .in2(_gnd_net_),
            .in3(N__5107),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_5_10_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_5_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__9053),
            .in2(N__5104),
            .in3(N__5077),
            .lcout(un5_visiblex_cry_7_c_RNIVZ0Z952),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_5_10_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_5_10_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(N__5062),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHS3_LC_5_10_2.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHS3_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHS3_LC_5_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHS3_LC_5_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5970),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_c_RNIFHSZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBT9_LC_5_10_3.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBT9_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBT9_LC_5_10_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBT9_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5305),
            .in3(N__5944),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNITBTZ0Z9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_5_10_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_5_10_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_3_LC_5_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_3_LC_5_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9539),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_s_2_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_67_LC_5_10_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_67_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_67_LC_5_10_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 Pixel_1_esr_RNO_67_LC_5_10_6 (
            .in0(N__9540),
            .in1(N__6263),
            .in2(N__10934),
            .in3(N__6191),
            .lcout(g0_0_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_5_10_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_5_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6254),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_5_11_0.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_5_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(N__6186),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOV5_LC_5_11_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOV5_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOV5_LC_5_11_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOV5_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5296),
            .in3(N__5287),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1_c_RNIDOVZ0Z5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQ06_LC_5_11_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQ06_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQ06_LC_5_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQ06_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(N__9035),
            .in2(N__5341),
            .in3(N__5284),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_RNIEQZ0Z06),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_5_11_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_5_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_5_11_3 (
            .in0(_gnd_net_),
            .in1(N__9544),
            .in2(_gnd_net_),
            .in3(N__5281),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_5_11_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_5_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_5_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5278),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_5_11_5.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_5_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_5_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9546),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_5_11_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_5_11_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9563),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_5_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_2_LC_5_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_2_LC_5_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9545),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_5_12_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_5_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__6196),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_5_12_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_5_12_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(N__5332),
            .in2(_gnd_net_),
            .in3(N__5326),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_5_12_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_5_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__5323),
            .in2(N__9052),
            .in3(N__5317),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_5_12_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_5_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_5_12_3 (
            .in0(_gnd_net_),
            .in1(N__9565),
            .in2(_gnd_net_),
            .in3(N__5314),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_5_12_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_5_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5311),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO),
            .ltout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_5_12_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_5_12_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_5_12_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_5_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5308),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_12_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_12_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_5_13_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_5_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_5_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_5_13_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_5_13_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_5_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_5_13_1 (
            .in0(_gnd_net_),
            .in1(N__5404),
            .in2(N__6151),
            .in3(N__5398),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_5_13_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_5_13_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_5_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_5_13_2 (
            .in0(_gnd_net_),
            .in1(N__5358),
            .in2(N__5395),
            .in3(N__5386),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_5_13_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_5_13_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_5_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_5_13_3 (
            .in0(N__6324),
            .in1(N__5347),
            .in2(N__5383),
            .in3(N__5374),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_5_13_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_5_13_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_5_13_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_5_13_4 (
            .in0(N__5371),
            .in1(N__5359),
            .in2(N__9579),
            .in3(N__5365),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31),
            .ltout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_5_13_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_5_13_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_5_13_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_5_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5362),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_5_13_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_5_13_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_5_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_5_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5357),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIM4P7_0_2_LC_6_4_0.C_ON=1'b0;
    defparam beamY_fast_RNIM4P7_0_2_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIM4P7_0_2_LC_6_4_0.LUT_INIT=16'b1000011100001111;
    LogicCell40 beamY_fast_RNIM4P7_0_2_LC_6_4_0 (
            .in0(N__8888),
            .in1(N__7931),
            .in2(N__8827),
            .in3(N__5487),
            .lcout(),
            .ltout(beamY_fast_RNIM4P7_0Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIO71D_3_LC_6_4_1.C_ON=1'b0;
    defparam beamY_fast_RNIO71D_3_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIO71D_3_LC_6_4_1.LUT_INIT=16'b1111000000110011;
    LogicCell40 beamY_fast_RNIO71D_3_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(N__8807),
            .in2(N__5506),
            .in3(N__5450),
            .lcout(beamY_fast_RNIO71DZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIM4P7_2_LC_6_4_4.C_ON=1'b0;
    defparam beamY_fast_RNIM4P7_2_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIM4P7_2_LC_6_4_4.LUT_INIT=16'b1110000110100101;
    LogicCell40 beamY_fast_RNIM4P7_2_LC_6_4_4 (
            .in0(N__8886),
            .in1(N__7930),
            .in2(N__8826),
            .in3(N__5486),
            .lcout(),
            .ltout(beamY_fast_RNIM4P7Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIJP9E_3_LC_6_4_5.C_ON=1'b0;
    defparam beamY_fast_RNIJP9E_3_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIJP9E_3_LC_6_4_5.LUT_INIT=16'b1111000010011001;
    LogicCell40 beamY_fast_RNIJP9E_3_LC_6_4_5 (
            .in0(N__8808),
            .in1(N__8887),
            .in2(N__5455),
            .in3(N__5449),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_6_4_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_6_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_6_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8340),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_6_5_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_6_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(N__6727),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9A1_LC_6_5_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9A1_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9A1_LC_6_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9A1_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(N__5599),
            .in2(N__9109),
            .in3(N__5416),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNIDT9AZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAA1_LC_6_5_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAA1_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAA1_LC_6_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAA1_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(N__6680),
            .in2(N__9110),
            .in3(N__5413),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNIEVAAZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_6_5_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_6_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5410),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_6_5_4.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_6_5_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_6_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5407),
            .in3(N__6558),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9KEQ_8_LC_6_5_5.C_ON=1'b0;
    defparam beamY_RNI9KEQ_8_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI9KEQ_8_LC_6_5_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 beamY_RNI9KEQ_8_LC_6_5_5 (
            .in0(N__6472),
            .in1(N__5614),
            .in2(_gnd_net_),
            .in3(N__7853),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIK0NV_9_LC_6_5_6.C_ON=1'b0;
    defparam beamY_RNIK0NV_9_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIK0NV_9_LC_6_5_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 beamY_RNIK0NV_9_LC_6_5_6 (
            .in0(N__7786),
            .in1(N__6798),
            .in2(_gnd_net_),
            .in3(N__5608),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIK0NV_0_9_LC_6_5_7.C_ON=1'b0;
    defparam beamY_RNIK0NV_0_9_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIK0NV_0_9_LC_6_5_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 beamY_RNIK0NV_0_9_LC_6_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5602),
            .in3(_gnd_net_),
            .lcout(beamY_RNIK0NV_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIPE7D_6_LC_6_6_2.C_ON=1'b0;
    defparam beamY_fast_RNIPE7D_6_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIPE7D_6_LC_6_6_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_fast_RNIPE7D_6_LC_6_6_2 (
            .in0(N__6820),
            .in1(N__7854),
            .in2(N__6493),
            .in3(N__6762),
            .lcout(),
            .ltout(un5_visibley_c7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUUSO1_9_LC_6_6_3.C_ON=1'b0;
    defparam beamY_RNIUUSO1_9_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIUUSO1_9_LC_6_6_3.LUT_INIT=16'b0000001010101000;
    LogicCell40 beamY_RNIUUSO1_9_LC_6_6_3 (
            .in0(N__6729),
            .in1(N__5593),
            .in2(N__5587),
            .in3(N__7787),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5tt_N_3_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_9_LC_6_6_4.C_ON=1'b0;
    defparam beamY_9_LC_6_6_4.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_6_6_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_9_LC_6_6_4 (
            .in0(N__8152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5584),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9820),
            .ce(N__8250),
            .sr(_gnd_net_));
    defparam beamY_fast_7_LC_6_6_5.C_ON=1'b0;
    defparam beamY_fast_7_LC_6_6_5.SEQ_MODE=4'b1000;
    defparam beamY_fast_7_LC_6_6_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 beamY_fast_7_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(N__8153),
            .in2(_gnd_net_),
            .in3(N__5566),
            .lcout(beamY_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9820),
            .ce(N__8250),
            .sr(_gnd_net_));
    defparam beamY_8_LC_6_6_6.C_ON=1'b0;
    defparam beamY_8_LC_6_6_6.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_6_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_8_LC_6_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5548),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9820),
            .ce(N__8250),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI1QVS_9_LC_6_6_7.C_ON=1'b0;
    defparam beamY_fast_RNI1QVS_9_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI1QVS_9_LC_6_6_7.LUT_INIT=16'b1010011110001111;
    LogicCell40 beamY_fast_RNI1QVS_9_LC_6_6_7 (
            .in0(N__7855),
            .in1(N__5530),
            .in2(N__5521),
            .in3(N__8764),
            .lcout(beamY_fast_RNI1QVSZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9N7M7_5_LC_6_7_0.C_ON=1'b0;
    defparam beamY_RNI9N7M7_5_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI9N7M7_5_LC_6_7_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNI9N7M7_5_LC_6_7_0 (
            .in0(N__8412),
            .in1(N__7027),
            .in2(N__7003),
            .in3(N__7520),
            .lcout(beamY_RNI9N7M7Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2GUN3_1_9_LC_6_7_1.C_ON=1'b0;
    defparam beamY_RNI2GUN3_1_9_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI2GUN3_1_9_LC_6_7_1.LUT_INIT=16'b0100010110101110;
    LogicCell40 beamY_RNI2GUN3_1_9_LC_6_7_1 (
            .in0(N__5756),
            .in1(N__8409),
            .in2(N__8476),
            .in3(N__8324),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un47_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI3M5H7_0_3_LC_6_7_2.C_ON=1'b0;
    defparam beamY_fast_RNI3M5H7_0_3_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI3M5H7_0_3_LC_6_7_2.LUT_INIT=16'b0101000000000101;
    LogicCell40 beamY_fast_RNI3M5H7_0_3_LC_6_7_2 (
            .in0(N__8410),
            .in1(_gnd_net_),
            .in2(N__5743),
            .in3(N__7026),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un54_sum_ac0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0RA9O_5_LC_6_7_3.C_ON=1'b0;
    defparam beamY_RNI0RA9O_5_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI0RA9O_5_LC_6_7_3.LUT_INIT=16'b0011011000111100;
    LogicCell40 beamY_RNI0RA9O_5_LC_6_7_3 (
            .in0(N__7519),
            .in1(N__6967),
            .in2(N__5722),
            .in3(N__6637),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIRRO4H1_3_LC_6_7_4.C_ON=1'b0;
    defparam beamY_RNIRRO4H1_3_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIRRO4H1_3_LC_6_7_4.LUT_INIT=16'b0111101100000000;
    LogicCell40 beamY_RNIRRO4H1_3_LC_6_7_4 (
            .in0(N__6638),
            .in1(N__7666),
            .in2(N__5719),
            .in3(N__5716),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un68_sum_c5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKUC181_0_5_LC_6_7_5.C_ON=1'b0;
    defparam beamY_RNIKUC181_0_5_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIKUC181_0_5_LC_6_7_5.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNIKUC181_0_5_LC_6_7_5 (
            .in0(N__5633),
            .in1(N__5697),
            .in2(_gnd_net_),
            .in3(N__5667),
            .lcout(beamY_RNIKUC181_0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI779U3_5_LC_6_7_6.C_ON=1'b0;
    defparam beamY_RNI779U3_5_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI779U3_5_LC_6_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNI779U3_5_LC_6_7_6 (
            .in0(N__8411),
            .in1(N__7025),
            .in2(_gnd_net_),
            .in3(N__7518),
            .lcout(beamY_RNI779U3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKPNA02_5_LC_6_7_7.C_ON=1'b0;
    defparam beamY_RNIKPNA02_5_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIKPNA02_5_LC_6_7_7.LUT_INIT=16'b1000000101111110;
    LogicCell40 beamY_RNIKPNA02_5_LC_6_7_7 (
            .in0(N__5698),
            .in1(N__5668),
            .in2(N__5638),
            .in3(N__5894),
            .lcout(beamY_RNIKPNA02Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5AJJ02_3_LC_6_8_0.C_ON=1'b0;
    defparam beamY_RNI5AJJ02_3_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI5AJJ02_3_LC_6_8_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNI5AJJ02_3_LC_6_8_0 (
            .in0(N__5918),
            .in1(N__5896),
            .in2(N__7678),
            .in3(N__7522),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un68_sum_axb4_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5F8A81_3_LC_6_8_1.C_ON=1'b0;
    defparam beamY_RNI5F8A81_3_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI5F8A81_3_LC_6_8_1.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI5F8A81_3_LC_6_8_1 (
            .in0(N__7521),
            .in1(N__7672),
            .in2(_gnd_net_),
            .in3(N__5917),
            .lcout(),
            .ltout(beamY_RNI5F8A81Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7VNCG5_3_LC_6_8_2.C_ON=1'b0;
    defparam beamY_RNI7VNCG5_3_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI7VNCG5_3_LC_6_8_2.LUT_INIT=16'b1000000000001000;
    LogicCell40 beamY_RNI7VNCG5_3_LC_6_8_2 (
            .in0(N__8103),
            .in1(N__5844),
            .in2(N__5899),
            .in3(N__5895),
            .lcout(),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un68_sum_ac0_7_d_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIAJLT9A_3_LC_6_8_3.C_ON=1'b0;
    defparam beamY_RNIAJLT9A_3_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIAJLT9A_3_LC_6_8_3.LUT_INIT=16'b0011011011001001;
    LogicCell40 beamY_RNIAJLT9A_3_LC_6_8_3 (
            .in0(N__5872),
            .in1(N__5853),
            .in2(N__5866),
            .in3(N__5863),
            .lcout(beamY_RNIAJLT9AZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1UL7G5_3_LC_6_8_4.C_ON=1'b0;
    defparam beamY_RNI1UL7G5_3_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI1UL7G5_3_LC_6_8_4.LUT_INIT=16'b1101110001010000;
    LogicCell40 beamY_RNI1UL7G5_3_LC_6_8_4 (
            .in0(N__7673),
            .in1(N__8104),
            .in2(N__5857),
            .in3(N__5845),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un68_sum_c4),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un68_sum_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQBCMCE_3_LC_6_8_5.C_ON=1'b0;
    defparam beamY_RNIQBCMCE_3_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIQBCMCE_3_LC_6_8_5.LUT_INIT=16'b0101101001101001;
    LogicCell40 beamY_RNIQBCMCE_3_LC_6_8_5 (
            .in0(N__5790),
            .in1(N__5836),
            .in2(N__5824),
            .in3(N__5821),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_axbxc5_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISDALMO_2_LC_6_8_7.C_ON=1'b0;
    defparam beamY_RNISDALMO_2_LC_6_8_7.SEQ_MODE=4'b0000;
    defparam beamY_RNISDALMO_2_LC_6_8_7.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNISDALMO_2_LC_6_8_7 (
            .in0(N__5803),
            .in1(N__5797),
            .in2(N__5791),
            .in3(N__6853),
            .lcout(font_un42_pixel_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_9_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__9718),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_6_9_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_6_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_6_9_1 (
            .in0(_gnd_net_),
            .in1(N__5982),
            .in2(N__5779),
            .in3(N__5764),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_60_LC_6_9_2.C_ON=1'b1;
    defparam Pixel_1_esr_RNO_60_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_60_LC_6_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_esr_RNO_60_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__7213),
            .in2(N__7111),
            .in3(N__5761),
            .lcout(Pixel_1_esr_RNOZ0Z_60),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_6_9_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_6_9_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_6_9_3 (
            .in0(N__7212),
            .in1(N__5983),
            .in2(N__7252),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOC_LC_6_9_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOC_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOC_LC_6_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOC_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__7237),
            .in2(_gnd_net_),
            .in3(N__5974),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNILFQOCZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIO1J8_LC_6_9_5.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIO1J8_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIO1J8_LC_6_9_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 un5_visiblex_cry_7_c_RNIO1J8_LC_6_9_5 (
            .in0(N__6262),
            .in1(N__6193),
            .in2(N__10933),
            .in3(N__9562),
            .lcout(G_25_i_o8_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_21_LC_6_9_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_21_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_21_LC_6_9_6.LUT_INIT=16'b1110111000000000;
    LogicCell40 Pixel_1_esr_RNO_21_LC_6_9_6 (
            .in0(N__10829),
            .in1(N__9719),
            .in2(_gnd_net_),
            .in3(N__9639),
            .lcout(G_25_i_a8_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_65_LC_6_9_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_65_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_65_LC_6_9_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 Pixel_1_esr_RNO_65_LC_6_9_7 (
            .in0(N__6261),
            .in1(N__6192),
            .in2(N__10932),
            .in3(N__9561),
            .lcout(g0_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNISG94_LC_6_10_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNISG94_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNISG94_LC_6_10_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un5_visiblex_cry_7_c_RNISG94_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(N__6252),
            .in2(_gnd_net_),
            .in3(N__6194),
            .lcout(un22_visibley_2),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2G_LC_6_10_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2G_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2G_LC_6_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2G_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(N__5971),
            .in2(N__6147),
            .in3(N__5959),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1_c_RNIOF2GZ0),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJ_LC_6_10_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJ_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJ_LC_6_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJ_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(N__6060),
            .in2(N__5956),
            .in3(N__5947),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI70UJZ0),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI273E1_LC_6_10_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI273E1_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI273E1_LC_6_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI273E1_LC_6_10_3 (
            .in0(N__6030),
            .in1(N__5943),
            .in2(N__5932),
            .in3(N__5923),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_LC_6_10_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_LC_6_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_LC_6_10_4 (
            .in0(N__6067),
            .in1(N__6061),
            .in2(N__9564),
            .in3(N__6052),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82KZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_0_LC_6_10_5.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_0_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_0_LC_6_10_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIB82K_0_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6049),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_8_LC_6_10_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_8_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_8_LC_6_10_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 Pixel_1_esr_RNO_8_LC_6_10_6 (
            .in0(N__6046),
            .in1(N__6253),
            .in2(_gnd_net_),
            .in3(N__6195),
            .lcout(g0_i_o4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_20_LC_6_10_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_20_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_20_LC_6_10_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 Pixel_1_esr_RNO_20_LC_6_10_7 (
            .in0(N__9726),
            .in1(N__11105),
            .in2(N__10548),
            .in3(N__10847),
            .lcout(un22_visibleylt9_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_6_11_0.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_6_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10941),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEM_LC_6_11_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEM_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEM_LC_6_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEM_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__6040),
            .in2(N__6000),
            .in3(N__6034),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1_c_RNIGCEMZ0),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICND41_LC_6_11_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICND41_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICND41_LC_6_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICND41_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(N__6031),
            .in2(N__6019),
            .in3(N__6010),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNICNDZ0Z41),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNI9KOM2_LC_6_11_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNI9KOM2_LC_6_11_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNI9KOM2_LC_6_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNI9KOM2_LC_6_11_3 (
            .in0(N__6126),
            .in1(N__6007),
            .in2(N__6001),
            .in3(N__5986),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_LC_6_11_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_LC_6_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(N__6208),
            .in2(_gnd_net_),
            .in3(N__6202),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEEZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_0_LC_6_11_5.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_0_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_0_LC_6_11_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIDAEE1_0_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6199),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_6_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_6_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_6_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6187),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIK454_LC_6_12_0.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIK454_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIK454_LC_6_12_0.LUT_INIT=16'b0001000100010001;
    LogicCell40 un5_visiblex_cry_5_c_RNIK454_LC_6_12_0 (
            .in0(N__10925),
            .in1(N__9640),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un22_visibley_3),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9J1_LC_6_12_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9J1_LC_6_12_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9J1_LC_6_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9J1_LC_6_12_1 (
            .in0(_gnd_net_),
            .in1(N__6334),
            .in2(N__6096),
            .in3(N__6130),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1_c_RNINV9JZ0Z1),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAM72_LC_6_12_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAM72_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAM72_LC_6_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAM72_LC_6_12_2 (
            .in0(_gnd_net_),
            .in1(N__6127),
            .in2(N__6115),
            .in3(N__6106),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_RNIDAMZ0Z72),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI53BF5_LC_6_12_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI53BF5_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI53BF5_LC_6_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI53BF5_LC_6_12_3 (
            .in0(N__7182),
            .in1(N__6103),
            .in2(N__6097),
            .in3(N__6082),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_LC_6_12_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_LC_6_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(N__6079),
            .in2(_gnd_net_),
            .in3(N__6073),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKPZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_0_LC_6_12_5.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_0_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_0_LC_6_12_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRBKP2_0_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6070),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_6_12_6.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_6_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_6_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9641),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_7.LUT_INIT=16'b0011001100110011;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(N__10924),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_13_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_13_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(N__10942),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_6_13_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_6_13_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_6_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_6_13_1 (
            .in0(_gnd_net_),
            .in1(N__6300),
            .in2(N__6217),
            .in3(N__6328),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_6_13_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_6_13_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_6_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(N__6325),
            .in2(N__6313),
            .in3(N__6304),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI31V25_LC_6_13_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI31V25_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI31V25_LC_6_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI31V25_LC_6_13_3 (
            .in0(N__7322),
            .in1(N__6301),
            .in2(N__6292),
            .in3(N__6283),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_6_13_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_6_13_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_6_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_6_13_4 (
            .in0(_gnd_net_),
            .in1(N__6280),
            .in2(_gnd_net_),
            .in3(N__6274),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_13_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_13_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_6_13_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_6_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6271),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_3_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__7516),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__6419),
            .in2(N__6361),
            .in3(N__6376),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__6343),
            .in2(N__6424),
            .in3(N__6373),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58S32_LC_7_3_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58S32_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58S32_LC_7_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58S32_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(N__6423),
            .in2(N__6460),
            .in3(N__6370),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI58SZ0Z32),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNISMP75_LC_7_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNISMP75_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNISMP75_LC_7_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNISMP75_LC_7_3_4 (
            .in0(N__7420),
            .in1(N__6400),
            .in2(N__6448),
            .in3(N__6367),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_LC_7_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_LC_7_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_LC_7_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_LC_7_3_5 (
            .in0(_gnd_net_),
            .in1(N__6436),
            .in2(_gnd_net_),
            .in3(N__6364),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_3_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_7_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8377),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_3_LC_7_3_7.C_ON=1'b0;
    defparam beamY_RNIBFP3_3_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_3_LC_7_3_7.LUT_INIT=16'b0111011110001000;
    LogicCell40 beamY_RNIBFP3_3_LC_7_3_7 (
            .in0(N__8034),
            .in1(N__8969),
            .in2(_gnd_net_),
            .in3(N__7958),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_4_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__8402),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_7_4_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_7_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__6514),
            .in2(N__6352),
            .in3(N__6337),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48A1_LC_7_4_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48A1_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48A1_LC_7_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48A1_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__6385),
            .in2(N__6520),
            .in3(N__6451),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNIL48AZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5Q1_LC_7_4_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5Q1_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5Q1_LC_7_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5Q1_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__6518),
            .in2(N__6589),
            .in3(N__6439),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIRH5QZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIGK8A2_LC_7_4_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIGK8A2_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIGK8A2_LC_7_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIGK8A2_LC_7_4_4 (
            .in0(N__6418),
            .in1(N__6499),
            .in2(N__6571),
            .in3(N__6430),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_7_4_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_7_4_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_7_4_5 (
            .in0(N__6538),
            .in1(N__6519),
            .in2(N__6559),
            .in3(N__6427),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_4_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_4_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_7_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6403),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9KEQ_0_8_LC_7_4_7.C_ON=1'b0;
    defparam beamY_RNI9KEQ_0_8_LC_7_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI9KEQ_0_8_LC_7_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 beamY_RNI9KEQ_0_8_LC_7_4_7 (
            .in0(N__6728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_RNI9KEQ_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_5_0 (
            .in0(_gnd_net_),
            .in1(N__8341),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8R_LC_7_5_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8R_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8R_LC_7_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8R_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(N__9102),
            .in2(N__6394),
            .in3(N__6379),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI0Q8RZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555B1_LC_7_5_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555B1_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555B1_LC_7_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555B1_LC_7_5_2 (
            .in0(_gnd_net_),
            .in1(N__6595),
            .in2(N__9111),
            .in3(N__6580),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNI555BZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797B1_LC_7_5_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797B1_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797B1_LC_7_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797B1_LC_7_5_3 (
            .in0(_gnd_net_),
            .in1(N__6577),
            .in2(N__9112),
            .in3(N__6562),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNI797BZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_5_4 (
            .in0(_gnd_net_),
            .in1(N__6554),
            .in2(_gnd_net_),
            .in3(N__6532),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_5_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_5_5 (
            .in0(_gnd_net_),
            .in1(N__6529),
            .in2(_gnd_net_),
            .in3(N__6523),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_5_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_5_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6502),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIRPUB_6_LC_7_5_7.C_ON=1'b0;
    defparam beamY_fast_RNIRPUB_6_LC_7_5_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIRPUB_6_LC_7_5_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamY_fast_RNIRPUB_6_LC_7_5_7 (
            .in0(N__6489),
            .in1(N__6819),
            .in2(_gnd_net_),
            .in3(N__6758),
            .lcout(un5_visibley_c6_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_0_5_LC_7_6_0.C_ON=1'b0;
    defparam beamY_RNI6125_0_5_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_0_5_LC_7_6_0.LUT_INIT=16'b0010010000000100;
    LogicCell40 beamY_RNI6125_0_5_LC_7_6_0 (
            .in0(N__8048),
            .in1(N__8914),
            .in2(N__7966),
            .in3(N__8996),
            .lcout(),
            .ltout(un11_visibleylto9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIICI12_5_LC_7_6_1.C_ON=1'b0;
    defparam beamY_RNIICI12_5_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIICI12_5_LC_7_6_1.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNIICI12_5_LC_7_6_1 (
            .in0(N__8415),
            .in1(N__8339),
            .in2(N__6466),
            .in3(N__6735),
            .lcout(),
            .ltout(un11_visibleylto9_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6D913_9_LC_7_6_2.C_ON=1'b0;
    defparam beamY_RNI6D913_9_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI6D913_9_LC_7_6_2.LUT_INIT=16'b0000000011110000;
    LogicCell40 beamY_RNI6D913_9_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6463),
            .in3(N__6689),
            .lcout(un11_visibley),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_6_LC_7_6_5.C_ON=1'b0;
    defparam beamY_fast_6_LC_7_6_5.SEQ_MODE=4'b1000;
    defparam beamY_fast_6_LC_7_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_6_LC_7_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6838),
            .lcout(beamY_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9823),
            .ce(N__8229),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIH5V7_6_LC_7_6_6.C_ON=1'b0;
    defparam beamY_fast_RNIH5V7_6_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIH5V7_6_LC_7_6_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 beamY_fast_RNIH5V7_6_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(N__6818),
            .in2(_gnd_net_),
            .in3(N__6757),
            .lcout(un5_visibley_c6_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_5_LC_7_6_7.C_ON=1'b0;
    defparam beamY_fast_5_LC_7_6_7.SEQ_MODE=4'b1000;
    defparam beamY_fast_5_LC_7_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_5_LC_7_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6787),
            .lcout(beamY_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9823),
            .ce(N__8229),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0DB_9_LC_7_7_0.C_ON=1'b0;
    defparam beamY_RNIJ0DB_9_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0DB_9_LC_7_7_0.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamY_RNIJ0DB_9_LC_7_7_0 (
            .in0(N__6961),
            .in1(N__7800),
            .in2(N__6610),
            .in3(N__7868),
            .lcout(beamY_RNIJ0DBZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIECTA3_8_LC_7_7_1.C_ON=1'b0;
    defparam beamY_RNIECTA3_8_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIECTA3_8_LC_7_7_1.LUT_INIT=16'b0011110010000111;
    LogicCell40 beamY_RNIECTA3_8_LC_7_7_1 (
            .in0(N__8343),
            .in1(N__6736),
            .in2(N__8470),
            .in3(N__6690),
            .lcout(beamY_RNIECTA3Z0Z_8),
            .ltout(beamY_RNIECTA3Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI3M5H7_3_LC_7_7_2.C_ON=1'b0;
    defparam beamY_fast_RNI3M5H7_3_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI3M5H7_3_LC_7_7_2.LUT_INIT=16'b1001011010010110;
    LogicCell40 beamY_fast_RNI3M5H7_3_LC_7_7_2 (
            .in0(N__8414),
            .in1(N__6995),
            .in2(N__6649),
            .in3(_gnd_net_),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un54_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICE7B5_4_LC_7_7_3.C_ON=1'b0;
    defparam beamY_RNICE7B5_4_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNICE7B5_4_LC_7_7_3.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNICE7B5_4_LC_7_7_3 (
            .in0(N__6601),
            .in1(N__7024),
            .in2(_gnd_net_),
            .in3(N__7959),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un75_sum_c5tt_m1_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_1_5_LC_7_7_4.C_ON=1'b0;
    defparam beamY_RNI6125_1_5_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_1_5_LC_7_7_4.LUT_INIT=16'b0000000000010101;
    LogicCell40 beamY_RNI6125_1_5_LC_7_7_4 (
            .in0(N__8846),
            .in1(N__9004),
            .in2(N__10345),
            .in3(N__8921),
            .lcout(un1_beamylto9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI4H1V1_0_9_LC_7_7_5.C_ON=1'b0;
    defparam beamY_fast_RNI4H1V1_0_9_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI4H1V1_0_9_LC_7_7_5.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_fast_RNI4H1V1_0_9_LC_7_7_5 (
            .in0(N__8344),
            .in1(N__8465),
            .in2(_gnd_net_),
            .in3(N__8413),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0),
            .ltout(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIKDT19_9_LC_7_7_6.C_ON=1'b0;
    defparam beamY_fast_RNIKDT19_9_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIKDT19_9_LC_7_7_6.LUT_INIT=16'b0110100101101001;
    LogicCell40 beamY_fast_RNIKDT19_9_LC_7_7_6 (
            .in0(N__7023),
            .in1(N__6994),
            .in2(N__6970),
            .in3(_gnd_net_),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un61_sum_axbxc5_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGKP3_7_LC_7_7_7.C_ON=1'b0;
    defparam beamY_RNIGKP3_7_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIGKP3_7_LC_7_7_7.LUT_INIT=16'b0000000000010001;
    LogicCell40 beamY_RNIGKP3_7_LC_7_7_7 (
            .in0(N__8065),
            .in1(N__8767),
            .in2(_gnd_net_),
            .in3(N__7960),
            .lcout(un1_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_46_LC_7_8_0.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_46_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_46_LC_7_8_0.LUT_INIT=16'b1001100010100010;
    LogicCell40 Pixel_1_esr_RNO_46_LC_7_8_0 (
            .in0(N__6946),
            .in1(N__9754),
            .in2(N__10849),
            .in3(N__6955),
            .lcout(un27lt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_45_LC_7_8_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_45_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_45_LC_7_8_1.LUT_INIT=16'b0101110110100010;
    LogicCell40 Pixel_1_esr_RNO_45_LC_7_8_1 (
            .in0(N__6954),
            .in1(N__6945),
            .in2(N__9763),
            .in3(N__6937),
            .lcout(un1_visiblex_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_52_LC_7_8_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_52_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_52_LC_7_8_2.LUT_INIT=16'b1100110001010101;
    LogicCell40 Pixel_1_esr_RNO_52_LC_7_8_2 (
            .in0(N__6872),
            .in1(N__6855),
            .in2(_gnd_net_),
            .in3(N__9007),
            .lcout(),
            .ltout(g1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_29_LC_7_8_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_29_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_29_LC_7_8_3.LUT_INIT=16'b1110000100011110;
    LogicCell40 Pixel_1_esr_RNO_29_LC_7_8_3 (
            .in0(N__10356),
            .in1(N__10034),
            .in2(N__6931),
            .in3(N__8060),
            .lcout(g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI34L6_10_LC_7_8_5.C_ON=1'b0;
    defparam beamX_RNI34L6_10_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam beamX_RNI34L6_10_LC_7_8_5.LUT_INIT=16'b0000000000000100;
    LogicCell40 beamX_RNI34L6_10_LC_7_8_5 (
            .in0(N__8636),
            .in1(N__8584),
            .in2(N__6928),
            .in3(N__6916),
            .lcout(un1_beamx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILTIMMO_3_LC_7_8_6.C_ON=1'b0;
    defparam beamY_RNILTIMMO_3_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNILTIMMO_3_LC_7_8_6.LUT_INIT=16'b0110011010100101;
    LogicCell40 beamY_RNILTIMMO_3_LC_7_8_6 (
            .in0(N__8059),
            .in1(N__6854),
            .in2(N__6874),
            .in3(N__9005),
            .lcout(font_un78_pixellto3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_50_LC_7_8_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_50_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_50_LC_7_8_7.LUT_INIT=16'b0100111010110001;
    LogicCell40 Pixel_1_esr_RNO_50_LC_7_8_7 (
            .in0(N__9006),
            .in1(N__6873),
            .in2(N__6859),
            .in3(N__8061),
            .lcout(g1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_0_LC_7_9_0.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_0_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_0_LC_7_9_0.LUT_INIT=16'b0100010000100010;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_0_LC_7_9_0 (
            .in0(N__10543),
            .in1(N__10722),
            .in2(_gnd_net_),
            .in3(N__10429),
            .lcout(),
            .ltout(r_i1_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI6J1NH2_0_LC_7_9_1.C_ON=1'b0;
    defparam beamX_RNI6J1NH2_0_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam beamX_RNI6J1NH2_0_LC_7_9_1.LUT_INIT=16'b1000110001001100;
    LogicCell40 beamX_RNI6J1NH2_0_LC_7_9_1 (
            .in0(N__10681),
            .in1(N__8544),
            .in2(N__7096),
            .in3(N__9121),
            .lcout(Pixel_3_sqmuxa_1_1),
            .ltout(Pixel_3_sqmuxa_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEC74VJ1_1_LC_7_9_2.C_ON=1'b0;
    defparam beamY_RNIEC74VJ1_1_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIEC74VJ1_1_LC_7_9_2.LUT_INIT=16'b0011000001100000;
    LogicCell40 beamY_RNIEC74VJ1_1_LC_7_9_2 (
            .in0(N__10358),
            .in1(N__7093),
            .in2(N__7087),
            .in3(N__10033),
            .lcout(Pixel_7_sqmuxa_1),
            .ltout(Pixel_7_sqmuxa_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_9_LC_7_9_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_9_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_9_LC_7_9_3.LUT_INIT=16'b0000000011101111;
    LogicCell40 Pixel_1_esr_RNO_9_LC_7_9_3 (
            .in0(N__7084),
            .in1(N__7131),
            .in2(N__7075),
            .in3(N__8512),
            .lcout(G_25_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_28_LC_7_9_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_28_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_28_LC_7_9_4.LUT_INIT=16'b0000000100001000;
    LogicCell40 Pixel_1_esr_RNO_28_LC_7_9_4 (
            .in0(N__10544),
            .in1(N__10723),
            .in2(N__7072),
            .in3(N__10430),
            .lcout(),
            .ltout(g0_0_4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_11_LC_7_9_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_11_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_11_LC_7_9_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 Pixel_1_esr_RNO_11_LC_7_9_5 (
            .in0(N__7057),
            .in1(N__7048),
            .in2(N__7051),
            .in3(N__7036),
            .lcout(G_25_i_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_27_LC_7_9_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_27_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_27_LC_7_9_6.LUT_INIT=16'b1101110110011001;
    LogicCell40 Pixel_1_esr_RNO_27_LC_7_9_6 (
            .in0(N__10217),
            .in1(N__10357),
            .in2(_gnd_net_),
            .in3(N__10032),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_49_LC_7_9_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_49_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_49_LC_7_9_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 Pixel_1_esr_RNO_49_LC_7_9_7 (
            .in0(N__7042),
            .in1(N__7159),
            .in2(_gnd_net_),
            .in3(N__7035),
            .lcout(g0_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_4_LC_7_10_0.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_4_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_4_LC_7_10_0.LUT_INIT=16'b0000000000101010;
    LogicCell40 Pixel_1_esr_RNO_4_LC_7_10_0 (
            .in0(N__7120),
            .in1(N__7279),
            .in2(N__7582),
            .in3(N__7294),
            .lcout(Pixel_9_u_ns_sn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_7_10_1.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_7_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_7_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11103),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_35_LC_7_10_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_35_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_35_LC_7_10_2.LUT_INIT=16'b1110111111011111;
    LogicCell40 Pixel_1_esr_RNO_35_LC_7_10_2 (
            .in0(N__10563),
            .in1(N__10359),
            .in2(N__10219),
            .in3(N__10442),
            .lcout(g1_0_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_15_LC_7_10_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_15_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_15_LC_7_10_3.LUT_INIT=16'b0010001000010001;
    LogicCell40 Pixel_1_esr_RNO_15_LC_7_10_3 (
            .in0(N__10443),
            .in1(N__10363),
            .in2(_gnd_net_),
            .in3(N__10564),
            .lcout(g1_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_24_LC_7_10_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_24_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_24_LC_7_10_4.LUT_INIT=16'b1001000000001001;
    LogicCell40 Pixel_1_esr_RNO_24_LC_7_10_4 (
            .in0(N__10677),
            .in1(N__10726),
            .in2(N__10578),
            .in3(N__10444),
            .lcout(G_25_i_a8_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_17_LC_7_10_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_17_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_17_LC_7_10_5.LUT_INIT=16'b1010101011101110;
    LogicCell40 Pixel_1_esr_RNO_17_LC_7_10_5 (
            .in0(N__10218),
            .in1(N__10076),
            .in2(_gnd_net_),
            .in3(N__10676),
            .lcout(g2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_64_LC_7_10_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_64_LC_7_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_64_LC_7_10_6.LUT_INIT=16'b0001000111001110;
    LogicCell40 Pixel_1_esr_RNO_64_LC_7_10_6 (
            .in0(N__10846),
            .in1(N__9762),
            .in2(N__9139),
            .in3(N__9657),
            .lcout(N_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_12_LC_7_10_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_12_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_12_LC_7_10_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_esr_RNO_12_LC_7_10_7 (
            .in0(N__7150),
            .in1(N__9268),
            .in2(N__7138),
            .in3(N__7119),
            .lcout(N_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_11_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_7_11_0 (
            .in0(_gnd_net_),
            .in1(N__9655),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_7_11_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_7_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_7_11_1 (
            .in0(_gnd_net_),
            .in1(N__7300),
            .in2(N__10861),
            .in3(N__7099),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_7_11_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_7_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(N__7327),
            .in2(N__7264),
            .in3(N__7240),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIP79LC_LC_7_11_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIP79LC_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIP79LC_LC_7_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIP79LC_LC_7_11_3 (
            .in0(N__7211),
            .in1(N__7333),
            .in2(N__7351),
            .in3(N__7228),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109G5_LC_7_11_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109G5_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109G5_LC_7_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109G5_LC_7_11_4 (
            .in0(_gnd_net_),
            .in1(N__7225),
            .in2(_gnd_net_),
            .in3(N__7216),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI109GZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_56_LC_7_11_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_56_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_56_LC_7_11_5.LUT_INIT=16'b1010101010001000;
    LogicCell40 Pixel_1_esr_RNO_56_LC_7_11_5 (
            .in0(N__9656),
            .in1(N__10843),
            .in2(_gnd_net_),
            .in3(N__9758),
            .lcout(un28_visibleylt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_37_LC_7_11_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_37_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_37_LC_7_11_6.LUT_INIT=16'b1011101111101110;
    LogicCell40 Pixel_1_esr_RNO_37_LC_7_11_6 (
            .in0(N__10675),
            .in1(N__10571),
            .in2(_gnd_net_),
            .in3(N__10445),
            .lcout(),
            .ltout(g0_10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_16_LC_7_11_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_16_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_16_LC_7_11_7.LUT_INIT=16'b1111000011110100;
    LogicCell40 Pixel_1_esr_RNO_16_LC_7_11_7 (
            .in0(N__10074),
            .in1(N__10192),
            .in2(N__7195),
            .in3(N__10368),
            .lcout(g1_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(N__9752),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17M43_LC_7_12_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17M43_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17M43_LC_7_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17M43_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(N__7192),
            .in2(N__7380),
            .in3(N__7186),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1_c_RNI17MZ0Z43),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VL4_LC_7_12_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VL4_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VL4_LC_7_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VL4_LC_7_12_2 (
            .in0(_gnd_net_),
            .in1(N__7183),
            .in2(N__7171),
            .in3(N__7162),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI08VLZ0Z4),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNICOQ2B_LC_7_12_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNICOQ2B_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNICOQ2B_LC_7_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNICOQ2B_LC_7_12_3 (
            .in0(N__9390),
            .in1(N__7387),
            .in2(N__7381),
            .in3(N__7366),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_LC_7_12_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_LC_7_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_LC_7_12_4 (
            .in0(_gnd_net_),
            .in1(N__7363),
            .in2(_gnd_net_),
            .in3(N__7357),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EOZ0Z5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_0_LC_7_12_5.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_0_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_0_LC_7_12_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIL3EO5_0_LC_7_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7354),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KK4_LC_7_12_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KK4_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KK4_LC_7_12_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KK4_LC_7_12_6 (
            .in0(N__7347),
            .in1(_gnd_net_),
            .in2(N__7326),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI77KKZ0Z4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_7_12_7.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_7_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_7_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7318),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_13_LC_7_13_0.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_13_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_13_LC_7_13_0.LUT_INIT=16'b0000000111000101;
    LogicCell40 Pixel_1_esr_RNO_13_LC_7_13_0 (
            .in0(N__7588),
            .in1(N__7275),
            .in2(N__7531),
            .in3(N__7572),
            .lcout(Pixel_9_sn_N_7_mux_1_tz),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIVFV5_LC_7_13_1.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIVFV5_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIVFV5_LC_7_13_1.LUT_INIT=16'b1100110010001000;
    LogicCell40 un5_visiblex_cry_1_c_RNIVFV5_LC_7_13_1 (
            .in0(N__10844),
            .in1(N__9760),
            .in2(_gnd_net_),
            .in3(N__11106),
            .lcout(),
            .ltout(un16_visibleylt9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNISDFC_LC_7_13_2.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNISDFC_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNISDFC_LC_7_13_2.LUT_INIT=16'b0000000000001100;
    LogicCell40 un5_visiblex_cry_8_c_RNISDFC_LC_7_13_2 (
            .in0(_gnd_net_),
            .in1(N__7550),
            .in2(N__7282),
            .in3(N__9580),
            .lcout(un16_visibley_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_33_LC_7_13_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_33_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_33_LC_7_13_5.LUT_INIT=16'b0000000100000000;
    LogicCell40 Pixel_1_esr_RNO_33_LC_7_13_5 (
            .in0(N__7597),
            .in1(N__10944),
            .in2(N__9586),
            .in3(N__7551),
            .lcout(Pixel_7_sqmuxa_3_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_55_LC_7_13_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_55_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_55_LC_7_13_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 Pixel_1_esr_RNO_55_LC_7_13_6 (
            .in0(N__9761),
            .in1(N__11107),
            .in2(N__10579),
            .in3(N__10845),
            .lcout(),
            .ltout(un22_visibleylt9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_32_LC_7_13_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_32_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_32_LC_7_13_7.LUT_INIT=16'b0000010000000000;
    LogicCell40 Pixel_1_esr_RNO_32_LC_7_13_7 (
            .in0(N__9584),
            .in1(N__7571),
            .in2(N__7555),
            .in3(N__7552),
            .lcout(un22_visibley),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_3_2.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_3_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7517),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_0_LC_8_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_0_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_0_LC_8_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIGVUJ2_0_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_4_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_4_0 (
            .in0(_gnd_net_),
            .in1(N__7622),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51F3_LC_8_4_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51F3_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51F3_LC_8_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51F3_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__7421),
            .in2(N__7447),
            .in3(N__7438),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIR51FZ0Z3),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNU3_LC_8_4_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNU3_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNU3_LC_8_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNU3_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__7435),
            .in2(N__7426),
            .in3(N__7429),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNICSNUZ0Z3),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKE4_LC_8_4_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKE4_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKE4_LC_8_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKE4_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(N__7425),
            .in2(N__7399),
            .in3(N__7390),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIRRKEZ0Z4),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIC4FVA_LC_8_4_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIC4FVA_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIC4FVA_LC_8_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIC4FVA_LC_8_4_4 (
            .in0(N__8505),
            .in1(N__7750),
            .in2(N__7744),
            .in3(N__7735),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_LC_8_4_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_LC_8_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_LC_8_4_5 (
            .in0(_gnd_net_),
            .in1(N__7732),
            .in2(_gnd_net_),
            .in3(N__7726),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANNZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_5_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(N__8092),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6V5_LC_8_5_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6V5_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6V5_LC_8_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6V5_LC_8_5_1 (
            .in0(_gnd_net_),
            .in1(N__8500),
            .in2(N__7606),
            .in3(N__7723),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIAG6VZ0Z5),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINI399_LC_8_5_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINI399_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINI399_LC_8_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINI399_LC_8_5_2 (
            .in0(_gnd_net_),
            .in1(N__7720),
            .in2(N__8506),
            .in3(N__7714),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNINIZ0Z399),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BRO9_LC_8_5_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BRO9_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BRO9_LC_8_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BRO9_LC_8_5_3 (
            .in0(_gnd_net_),
            .in1(N__8504),
            .in2(N__7711),
            .in3(N__7702),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI9BROZ0Z9),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAPMAL_LC_8_5_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAPMAL_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAPMAL_LC_8_5_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIAPMAL_LC_8_5_4 (
            .in0(N__9443),
            .in1(N__8482),
            .in2(N__7699),
            .in3(N__7690),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1B_LC_8_5_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1B_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1B_LC_8_5_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1B_LC_8_5_5 (
            .in0(_gnd_net_),
            .in1(N__7687),
            .in2(_gnd_net_),
            .in3(N__7681),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIHCT1BZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_5_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7635),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_0_LC_8_5_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_0_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_0_LC_8_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIQANN5_0_LC_8_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8499),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI4H1V1_9_LC_8_6_0.C_ON=1'b0;
    defparam beamY_fast_RNI4H1V1_9_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI4H1V1_9_LC_8_6_0.LUT_INIT=16'b1000100011101110;
    LogicCell40 beamY_fast_RNI4H1V1_9_LC_8_6_0 (
            .in0(N__8475),
            .in1(N__8416),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(font_un42_pixel_if_generate_plus_mult1_un47_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2ROB_9_LC_8_6_1.C_ON=1'b0;
    defparam beamY_RNI2ROB_9_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI2ROB_9_LC_8_6_1.LUT_INIT=16'b0000000000010011;
    LogicCell40 beamY_RNI2ROB_9_LC_8_6_1 (
            .in0(N__7965),
            .in1(N__7801),
            .in2(N__8269),
            .in3(N__7870),
            .lcout(un8_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_8_6_2.C_ON=1'b0;
    defparam beamY_1_LC_8_6_2.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_8_6_2.LUT_INIT=16'b0101000001111000;
    LogicCell40 beamY_1_LC_8_6_2 (
            .in0(N__8254),
            .in1(N__10213),
            .in2(N__10346),
            .in3(N__8158),
            .lcout(un28lto1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9826),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_8_6_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_8_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8102),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_8_7_0.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_8_7_0.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIHUG2_0_3_LC_8_7_0 (
            .in0(N__8995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8047),
            .lcout(un4_beamylt6),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_5_LC_8_7_1.C_ON=1'b0;
    defparam beamY_RNI2KA6_5_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_5_LC_8_7_1.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI2KA6_5_LC_8_7_1 (
            .in0(N__8842),
            .in1(N__8922),
            .in2(N__7969),
            .in3(N__7961),
            .lcout(),
            .ltout(un4_beamylt8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_9_LC_8_7_2.C_ON=1'b0;
    defparam beamY_RNISI4A_9_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_9_LC_8_7_2.LUT_INIT=16'b1111111000000000;
    LogicCell40 beamY_RNISI4A_9_LC_8_7_2 (
            .in0(N__7880),
            .in1(N__8765),
            .in2(N__7813),
            .in3(N__7809),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_7_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_7_5 (
            .in0(N__9923),
            .in1(N__9095),
            .in2(_gnd_net_),
            .in3(N__8994),
            .lcout(beamY_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIMJIF_7_LC_8_7_6.C_ON=1'b0;
    defparam beamY_RNIMJIF_7_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIMJIF_7_LC_8_7_6.LUT_INIT=16'b0000000000000100;
    LogicCell40 beamY_RNIMJIF_7_LC_8_7_6 (
            .in0(N__8923),
            .in1(N__8854),
            .in2(N__8848),
            .in3(N__8766),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_3_LC_8_8_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_3_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_3_LC_8_8_1.LUT_INIT=16'b1111101111110000;
    LogicCell40 Pixel_1_esr_RNO_3_LC_8_8_1 (
            .in0(N__8560),
            .in1(N__8583),
            .in2(N__8698),
            .in3(N__8590),
            .lcout(),
            .ltout(Pixel_1_sqmuxa_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_0_LC_8_8_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_0_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_0_LC_8_8_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 Pixel_1_esr_RNO_0_LC_8_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8701),
            .in3(N__9875),
            .lcout(Pixel_1_sqmuxa_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_8_8_3.C_ON=1'b0;
    defparam HSync_1_LC_8_8_3.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_8_8_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 HSync_1_LC_8_8_3 (
            .in0(N__8697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9821),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNINAS01_10_LC_8_8_5.C_ON=1'b0;
    defparam beamX_RNINAS01_10_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam beamX_RNINAS01_10_LC_8_8_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNINAS01_10_LC_8_8_5 (
            .in0(N__8653),
            .in1(N__8647),
            .in2(N__8638),
            .in3(N__8596),
            .lcout(un15_beamy_2),
            .ltout(un15_beamy_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_44_LC_8_8_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_44_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_44_LC_8_8_6.LUT_INIT=16'b0000000011010000;
    LogicCell40 Pixel_1_esr_RNO_44_LC_8_8_6 (
            .in0(N__8582),
            .in1(N__8559),
            .in2(N__8548),
            .in3(N__8545),
            .lcout(),
            .ltout(Pixel_9_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_22_LC_8_8_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_22_LC_8_8_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_22_LC_8_8_7.LUT_INIT=16'b1110000000010000;
    LogicCell40 Pixel_1_esr_RNO_22_LC_8_8_7 (
            .in0(N__8527),
            .in1(N__8521),
            .in2(N__8515),
            .in3(N__9949),
            .lcout(Pixel_9_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_1_LC_8_9_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_1_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_1_LC_8_9_1.LUT_INIT=16'b1111111000010000;
    LogicCell40 Pixel_1_esr_RNO_1_LC_8_9_1 (
            .in0(N__9493),
            .in1(N__9244),
            .in2(N__9280),
            .in3(N__10585),
            .lcout(),
            .ltout(N_163_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_LC_8_9_2.C_ON=1'b0;
    defparam Pixel_1_esr_LC_8_9_2.SEQ_MODE=4'b1000;
    defparam Pixel_1_esr_LC_8_9_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 Pixel_1_esr_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__9232),
            .in2(N__9226),
            .in3(N__9145),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9816),
            .ce(N__9193),
            .sr(N__9889));
    defparam Pixel_1_esr_RNO_26_LC_8_9_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_26_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_26_LC_8_9_3.LUT_INIT=16'b0101011000000000;
    LogicCell40 Pixel_1_esr_RNO_26_LC_8_9_3 (
            .in0(N__9187),
            .in1(N__10070),
            .in2(N__10355),
            .in3(N__9181),
            .lcout(),
            .ltout(g0_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_10_LC_8_9_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_10_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_10_LC_8_9_4.LUT_INIT=16'b1111000001000000;
    LogicCell40 Pixel_1_esr_RNO_10_LC_8_9_4 (
            .in0(N__9253),
            .in1(N__9175),
            .in2(N__9169),
            .in3(N__10741),
            .lcout(),
            .ltout(G_25_i_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_2_LC_8_9_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_2_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_2_LC_8_9_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 Pixel_1_esr_RNO_2_LC_8_9_5 (
            .in0(N__9166),
            .in1(N__9160),
            .in2(N__9154),
            .in3(N__9151),
            .lcout(Pixel_9_u_ns_rn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_69_LC_8_10_0.C_ON=1'b1;
    defparam Pixel_1_esr_RNO_69_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_69_LC_8_10_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 Pixel_1_esr_RNO_69_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__10549),
            .in2(_gnd_net_),
            .in3(N__11104),
            .lcout(g2_1),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OT9_LC_8_10_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OT9_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OT9_LC_8_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OT9_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__9130),
            .in2(N__9330),
            .in3(N__9124),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI3OTZ0Z9),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JF21_LC_8_10_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JF21_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JF21_LC_8_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JF21_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__11041),
            .in2(N__10963),
            .in3(N__9115),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNI39JFZ0Z21),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3 (
            .in0(_gnd_net_),
            .in1(N__11011),
            .in2(N__9331),
            .in3(N__10958),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QB1_LC_8_10_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QB1_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QB1_LC_8_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QB1_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(N__10981),
            .in2(_gnd_net_),
            .in3(N__9316),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIK64QBZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_34_LC_8_10_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_34_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_34_LC_8_10_5.LUT_INIT=16'b1010111101010000;
    LogicCell40 Pixel_1_esr_RNO_34_LC_8_10_5 (
            .in0(N__10550),
            .in1(_gnd_net_),
            .in2(N__9313),
            .in3(N__10727),
            .lcout(),
            .ltout(font_un19_pixel_0_0_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_14_LC_8_10_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_14_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_14_LC_8_10_6.LUT_INIT=16'b1111111000001110;
    LogicCell40 Pixel_1_esr_RNO_14_LC_8_10_6 (
            .in0(N__10075),
            .in1(N__9310),
            .in2(N__9304),
            .in3(N__9400),
            .lcout(),
            .ltout(font_un237_pixel_6_ns_1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_5_LC_8_10_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_5_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_5_LC_8_10_7.LUT_INIT=16'b1000111110000000;
    LogicCell40 Pixel_1_esr_RNO_5_LC_8_10_7 (
            .in0(N__9301),
            .in1(N__9295),
            .in2(N__9289),
            .in3(N__9286),
            .lcout(font_un237_pixel_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_54_LC_8_11_0.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_54_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_54_LC_8_11_0.LUT_INIT=16'b1101111011101101;
    LogicCell40 Pixel_1_esr_RNO_54_LC_8_11_0 (
            .in0(N__10574),
            .in1(N__9262),
            .in2(N__10446),
            .in3(N__10682),
            .lcout(),
            .ltout(g2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_31_LC_8_11_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_31_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_31_LC_8_11_1.LUT_INIT=16'b1111000011010000;
    LogicCell40 Pixel_1_esr_RNO_31_LC_8_11_1 (
            .in0(N__10214),
            .in1(N__10350),
            .in2(N__9271),
            .in3(N__10073),
            .lcout(font_un83_pixel_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_LC_8_11_3.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_LC_8_11_3.LUT_INIT=16'b1100001111110000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un75_sum_cry_1_c_RNI8JV5C1_LC_8_11_3 (
            .in0(_gnd_net_),
            .in1(N__10573),
            .in2(N__10729),
            .in3(N__10422),
            .lcout(font_un19_pixel_23),
            .ltout(font_un19_pixel_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_25_LC_8_11_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_25_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_25_LC_8_11_4.LUT_INIT=16'b0001001101100100;
    LogicCell40 Pixel_1_esr_RNO_25_LC_8_11_4 (
            .in0(N__10072),
            .in1(N__10215),
            .in2(N__9256),
            .in3(N__10354),
            .lcout(font_un160_pixel_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_57_LC_8_11_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_57_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_57_LC_8_11_6.LUT_INIT=16'b0100100001001000;
    LogicCell40 Pixel_1_esr_RNO_57_LC_8_11_6 (
            .in0(N__10575),
            .in1(N__10683),
            .in2(N__10447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(g0_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_36_LC_8_11_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_36_LC_8_11_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_36_LC_8_11_7.LUT_INIT=16'b1110000001010000;
    LogicCell40 Pixel_1_esr_RNO_36_LC_8_11_7 (
            .in0(N__10216),
            .in1(N__10351),
            .in2(N__9403),
            .in3(N__10071),
            .lcout(g3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_8_12_0.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_8_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_LC_8_12_0 (
            .in0(_gnd_net_),
            .in1(N__10836),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4M96_LC_8_12_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4M96_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4M96_LC_8_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4M96_LC_8_12_1 (
            .in0(_gnd_net_),
            .in1(N__9667),
            .in2(N__9360),
            .in3(N__9394),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1_c_RNIN4MZ0Z96),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCC9_LC_8_12_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCC9_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCC9_LC_8_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCC9_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(N__9391),
            .in2(N__9379),
            .in3(N__9370),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI2GCCZ0Z9),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNISKRFM_LC_8_12_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNISKRFM_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNISKRFM_LC_8_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNISKRFM_LC_8_12_3 (
            .in0(N__11031),
            .in1(N__9367),
            .in2(N__9361),
            .in3(N__9346),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_LC_8_12_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_LC_8_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_LC_8_12_4 (
            .in0(_gnd_net_),
            .in1(N__9343),
            .in2(_gnd_net_),
            .in3(N__9337),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0),
            .ltout(font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_0_LC_8_12_5.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_0_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_0_LC_8_12_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQ15IB_0_LC_8_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9334),
            .in3(_gnd_net_),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_8_12_7.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_8_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_8_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9753),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_7_LC_8_13_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_7_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_7_LC_8_13_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 Pixel_1_esr_RNO_7_LC_8_13_5 (
            .in0(N__9661),
            .in1(N__10945),
            .in2(_gnd_net_),
            .in3(N__9585),
            .lcout(g0_i_o4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_6_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9924),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEB_LC_9_6_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEB_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEB_LC_9_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEB_LC_9_6_1 (
            .in0(_gnd_net_),
            .in1(N__9484),
            .in2(N__9444),
            .in3(N__9478),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI68NEBZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9H_LC_9_6_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9H_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9H_LC_9_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9H_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(N__9439),
            .in2(N__9475),
            .in3(N__9466),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIR7M9HZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_62_LC_9_6_3.C_ON=1'b1;
    defparam Pixel_1_esr_RNO_62_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_62_LC_9_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_esr_RNO_62_LC_9_6_3 (
            .in0(_gnd_net_),
            .in1(N__9463),
            .in2(N__9445),
            .in3(N__9457),
            .lcout(Pixel_1_esr_RNOZ0Z_62),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_6_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_6_4 (
            .in0(_gnd_net_),
            .in1(N__9418),
            .in2(N__9454),
            .in3(N__9435),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJL_LC_9_6_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJL_LC_9_6_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJL_LC_9_6_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJL_LC_9_6_5 (
            .in0(_gnd_net_),
            .in1(N__9412),
            .in2(_gnd_net_),
            .in3(N__9406),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIDACJLZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_68_LC_9_7_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_68_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_68_LC_9_7_1.LUT_INIT=16'b0001100010001000;
    LogicCell40 Pixel_1_esr_RNO_68_LC_9_7_1 (
            .in0(N__9933),
            .in1(N__9942),
            .in2(N__9925),
            .in3(N__9959),
            .lcout(),
            .ltout(un28lto4_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_63_LC_9_7_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_63_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_63_LC_9_7_2.LUT_INIT=16'b1000000001000000;
    LogicCell40 Pixel_1_esr_RNO_63_LC_9_7_2 (
            .in0(N__9960),
            .in1(N__10261),
            .in2(N__9973),
            .in3(N__9922),
            .lcout(),
            .ltout(un28lt10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_47_LC_9_7_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_47_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_47_LC_9_7_3.LUT_INIT=16'b0000011000000101;
    LogicCell40 Pixel_1_esr_RNO_47_LC_9_7_3 (
            .in0(N__9970),
            .in1(N__9895),
            .in2(N__9964),
            .in3(N__9961),
            .lcout(un28_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_61_LC_9_7_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_61_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_61_LC_9_7_6.LUT_INIT=16'b1110111011111111;
    LogicCell40 Pixel_1_esr_RNO_61_LC_9_7_6 (
            .in0(N__9943),
            .in1(N__9934),
            .in2(_gnd_net_),
            .in3(N__9921),
            .lcout(un1_beamY_if_generate_plus_mult1_un1_rem_adjust_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_9_8_4.C_ON=1'b0;
    defparam VSync_1_LC_9_8_4.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_9_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 VSync_1_LC_9_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9888),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9824),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_39_LC_9_8_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_39_LC_9_8_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_39_LC_9_8_6.LUT_INIT=16'b0010001001100110;
    LogicCell40 Pixel_1_esr_RNO_39_LC_9_8_6 (
            .in0(N__10305),
            .in1(N__10191),
            .in2(_gnd_net_),
            .in3(N__10046),
            .lcout(Pixel_1_esr_RNOZ0Z_39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_58_LC_9_9_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_58_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_58_LC_9_9_1.LUT_INIT=16'b0101101001011010;
    LogicCell40 Pixel_1_esr_RNO_58_LC_9_9_1 (
            .in0(N__10546),
            .in1(_gnd_net_),
            .in2(N__10448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(g1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_38_LC_9_9_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_38_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_38_LC_9_9_2.LUT_INIT=16'b0011110010101111;
    LogicCell40 Pixel_1_esr_RNO_38_LC_9_9_2 (
            .in0(N__10209),
            .in1(N__10319),
            .in2(N__9775),
            .in3(N__10063),
            .lcout(),
            .ltout(N_1304_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_18_LC_9_9_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_18_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_18_LC_9_9_3.LUT_INIT=16'b1110001010111000;
    LogicCell40 Pixel_1_esr_RNO_18_LC_9_9_3 (
            .in0(N__9772),
            .in1(N__10750),
            .in2(N__9766),
            .in3(N__10725),
            .lcout(N_156_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_40_LC_9_9_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_40_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_40_LC_9_9_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 Pixel_1_esr_RNO_40_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(N__10545),
            .in2(_gnd_net_),
            .in3(N__10431),
            .lcout(g1_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_48_LC_9_9_5.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_48_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_48_LC_9_9_5.LUT_INIT=16'b0101000000001010;
    LogicCell40 Pixel_1_esr_RNO_48_LC_9_9_5 (
            .in0(N__10547),
            .in1(_gnd_net_),
            .in2(N__10449),
            .in3(N__10724),
            .lcout(),
            .ltout(N_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_23_LC_9_9_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_23_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_23_LC_9_9_6.LUT_INIT=16'b0000000001100000;
    LogicCell40 Pixel_1_esr_RNO_23_LC_9_9_6 (
            .in0(N__10210),
            .in1(N__10320),
            .in2(N__10744),
            .in3(N__10064),
            .lcout(G_25_i_a8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_59_LC_9_10_1.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_59_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_59_LC_9_10_1.LUT_INIT=16'b0101101001011010;
    LogicCell40 Pixel_1_esr_RNO_59_LC_9_10_1 (
            .in0(N__10577),
            .in1(_gnd_net_),
            .in2(N__10450),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(g1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_41_LC_9_10_2.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_41_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_41_LC_9_10_2.LUT_INIT=16'b1100011101111110;
    LogicCell40 Pixel_1_esr_RNO_41_LC_9_10_2 (
            .in0(N__10078),
            .in1(N__10212),
            .in2(N__10735),
            .in3(N__10353),
            .lcout(),
            .ltout(N_1302_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_19_LC_9_10_3.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_19_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_19_LC_9_10_3.LUT_INIT=16'b1110001010111000;
    LogicCell40 Pixel_1_esr_RNO_19_LC_9_10_3 (
            .in0(N__9979),
            .in1(N__10375),
            .in2(N__10732),
            .in3(N__10728),
            .lcout(),
            .ltout(N_159_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_6_LC_9_10_4.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_6_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_6_LC_9_10_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 Pixel_1_esr_RNO_6_LC_9_10_4 (
            .in0(_gnd_net_),
            .in1(N__10684),
            .in2(N__10594),
            .in3(N__10591),
            .lcout(font_un314_pixel_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_43_LC_9_10_6.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_43_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_43_LC_9_10_6.LUT_INIT=16'b1111111100110011;
    LogicCell40 Pixel_1_esr_RNO_43_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(N__10576),
            .in2(_gnd_net_),
            .in3(N__10438),
            .lcout(g1_3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_esr_RNO_42_LC_9_10_7.C_ON=1'b0;
    defparam Pixel_1_esr_RNO_42_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam Pixel_1_esr_RNO_42_LC_9_10_7.LUT_INIT=16'b0010001001100110;
    LogicCell40 Pixel_1_esr_RNO_42_LC_9_10_7 (
            .in0(N__10352),
            .in1(N__10211),
            .in2(_gnd_net_),
            .in3(N__10077),
            .lcout(N_1303_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_11_0.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(N__11095),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLB_LC_9_11_1.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLB_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLB_LC_9_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLB_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(N__10756),
            .in2(N__10995),
            .in3(N__11035),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1_c_RNI1KSLBZ0),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTH_LC_9_11_2.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTH_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTH_LC_9_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTH_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(N__11032),
            .in2(N__11020),
            .in3(N__11005),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_RNI40KTHZ0),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI102IB1_LC_9_11_3.C_ON=1'b1;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI102IB1_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI102IB1_LC_9_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI102IB1_LC_9_11_3 (
            .in0(N__10962),
            .in1(N__11002),
            .in2(N__10996),
            .in3(N__10975),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHM_LC_9_11_4.C_ON=1'b0;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHM_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHM_LC_9_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHM_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(N__10972),
            .in2(_gnd_net_),
            .in3(N__10966),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIHIMHMZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_11_6.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_9_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_9_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10943),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_9_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_9_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10848),
            .lcout(font_un19_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
