// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 18:20:45

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4848;
    wire N__4847;
    wire N__4846;
    wire N__4839;
    wire N__4838;
    wire N__4837;
    wire N__4830;
    wire N__4829;
    wire N__4828;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4715;
    wire N__4712;
    wire N__4711;
    wire N__4706;
    wire N__4703;
    wire N__4702;
    wire N__4699;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4681;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4669;
    wire N__4666;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4645;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4633;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4551;
    wire N__4546;
    wire N__4541;
    wire N__4538;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4530;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4471;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4418;
    wire N__4417;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4381;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4331;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4299;
    wire N__4298;
    wire N__4297;
    wire N__4296;
    wire N__4295;
    wire N__4294;
    wire N__4291;
    wire N__4290;
    wire N__4289;
    wire N__4286;
    wire N__4279;
    wire N__4276;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4261;
    wire N__4260;
    wire N__4257;
    wire N__4252;
    wire N__4243;
    wire N__4240;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4190;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4178;
    wire N__4177;
    wire N__4174;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4150;
    wire N__4147;
    wire N__4146;
    wire N__4145;
    wire N__4142;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4128;
    wire N__4125;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4107;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4058;
    wire N__4055;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__4049;
    wire N__4048;
    wire N__4047;
    wire N__4046;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3889;
    wire N__3888;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3880;
    wire N__3877;
    wire N__3868;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3796;
    wire N__3793;
    wire N__3792;
    wire N__3791;
    wire N__3784;
    wire N__3781;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3736;
    wire N__3733;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3697;
    wire N__3694;
    wire N__3693;
    wire N__3692;
    wire N__3685;
    wire N__3682;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3623;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3596;
    wire N__3595;
    wire N__3594;
    wire N__3593;
    wire N__3592;
    wire N__3589;
    wire N__3584;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3557;
    wire N__3556;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3533;
    wire N__3530;
    wire N__3521;
    wire N__3520;
    wire N__3519;
    wire N__3516;
    wire N__3511;
    wire N__3508;
    wire N__3507;
    wire N__3506;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3485;
    wire N__3482;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3458;
    wire N__3457;
    wire N__3454;
    wire N__3453;
    wire N__3450;
    wire N__3449;
    wire N__3448;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3433;
    wire N__3430;
    wire N__3419;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3411;
    wire N__3410;
    wire N__3405;
    wire N__3402;
    wire N__3401;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3389;
    wire N__3386;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3364;
    wire N__3363;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3351;
    wire N__3344;
    wire N__3343;
    wire N__3340;
    wire N__3339;
    wire N__3338;
    wire N__3335;
    wire N__3328;
    wire N__3323;
    wire N__3322;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3307;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3280;
    wire N__3277;
    wire N__3276;
    wire N__3275;
    wire N__3268;
    wire N__3265;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3232;
    wire N__3231;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3213;
    wire N__3210;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3152;
    wire N__3151;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3128;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3120;
    wire N__3119;
    wire N__3118;
    wire N__3117;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3083;
    wire N__3082;
    wire N__3081;
    wire N__3080;
    wire N__3079;
    wire N__3078;
    wire N__3073;
    wire N__3072;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3050;
    wire N__3047;
    wire N__3046;
    wire N__3043;
    wire N__3042;
    wire N__3041;
    wire N__3040;
    wire N__3039;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3019;
    wire N__3016;
    wire N__3005;
    wire N__3002;
    wire N__3001;
    wire N__3000;
    wire N__2999;
    wire N__2998;
    wire N__2997;
    wire N__2994;
    wire N__2989;
    wire N__2986;
    wire N__2981;
    wire N__2972;
    wire N__2969;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2945;
    wire N__2944;
    wire N__2943;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2918;
    wire N__2917;
    wire N__2916;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2904;
    wire N__2901;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2887;
    wire N__2886;
    wire N__2885;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2871;
    wire N__2868;
    wire N__2861;
    wire N__2858;
    wire N__2857;
    wire N__2856;
    wire N__2855;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2841;
    wire N__2838;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2804;
    wire N__2803;
    wire N__2802;
    wire N__2801;
    wire N__2796;
    wire N__2793;
    wire N__2792;
    wire N__2789;
    wire N__2784;
    wire N__2781;
    wire N__2774;
    wire N__2773;
    wire N__2772;
    wire N__2771;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2696;
    wire N__2693;
    wire N__2692;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2674;
    wire N__2669;
    wire N__2666;
    wire N__2665;
    wire N__2664;
    wire N__2661;
    wire N__2660;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2646;
    wire N__2643;
    wire N__2634;
    wire N__2631;
    wire N__2626;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2569;
    wire N__2568;
    wire N__2565;
    wire N__2562;
    wire N__2559;
    wire N__2556;
    wire N__2549;
    wire N__2548;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2540;
    wire N__2537;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2455;
    wire N__2454;
    wire N__2453;
    wire N__2444;
    wire N__2443;
    wire N__2442;
    wire N__2439;
    wire N__2434;
    wire N__2429;
    wire N__2428;
    wire N__2427;
    wire N__2426;
    wire N__2423;
    wire N__2422;
    wire N__2413;
    wire N__2410;
    wire N__2409;
    wire N__2406;
    wire N__2401;
    wire N__2396;
    wire N__2395;
    wire N__2392;
    wire N__2389;
    wire N__2388;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire VCCG0;
    wire \Clock50MHz.PixelClock ;
    wire Clock12MHz_c;
    wire GNDG0;
    wire bfn_7_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_;
    wire bfn_7_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire un5_visibley_cry_8_c_RNI3O5CZ0Z_0;
    wire un5_visibley_cry_7_c_RNI1L4CZ0Z_0;
    wire bfn_7_4_0_;
    wire un21_beamy_cry_1;
    wire beamY_RNO_0Z0Z_3;
    wire un21_beamy_cry_2;
    wire beamY_RNO_0Z0Z_4;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire beamY_RNO_0Z0Z_7;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire bfn_7_5_0_;
    wire beamY_RNO_0Z0Z_9;
    wire un3_beamx_5_cascade_;
    wire un3_beamx_7;
    wire beamY_RNO_0Z0Z_1;
    wire un5_beamx_3_0;
    wire un5_beamx_4;
    wire beamYZ0Z_0;
    wire bfn_7_7_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_7_8_0_;
    wire beamX_RNI5457Z0Z_5;
    wire un8_beamx_cry_9;
    wire bfn_8_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_axb_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_0;
    wire bfn_8_3_0_;
    wire un5_visibley_cry_2;
    wire un5_visibley_cry_3;
    wire un5_visibley_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un47_sum;
    wire un5_visibley_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un40_sum;
    wire un5_visibley_cry_6;
    wire un5_visibley_cry_7_c_RNI1L4CZ0;
    wire un5_visibley_cry_7;
    wire un5_visibley_cry_8;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_axb_3;
    wire beamYZ0Z_6;
    wire beamYZ0Z_5;
    wire un4_beamylt6_cascade_;
    wire un4_beamylt8_0_cascade_;
    wire beamYZ0Z_3;
    wire un1_beamylto9_2_cascade_;
    wire beamYZ0Z_4;
    wire VSync_c;
    wire beamYZ0Z_9;
    wire beamYZ0Z_8;
    wire un18_beamylt4;
    wire un18_beamylt4_cascade_;
    wire un13_beamylt7_cascade_;
    wire un8_beamy_2;
    wire un1_beamy_4;
    wire beamYZ0Z_7;
    wire un5_beamx_3;
    wire un8_beamylto9_1_cascade_;
    wire beamYZ0Z_2;
    wire bfn_8_6_0_;
    wire beamXZ0Z_0;
    wire beamXZ0Z_1;
    wire un5_visiblex_cry_0;
    wire beamXZ0Z_2;
    wire un5_visiblex_cry_1;
    wire un5_visiblex_cry_2;
    wire un5_visiblex_cry_3;
    wire un5_visiblex_cry_4;
    wire un5_visiblex_cry_5;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire bfn_8_7_0_;
    wire un5_visiblex_cry_8;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_;
    wire beamXZ0Z_5;
    wire beamXZ0Z_4;
    wire beamXZ0Z_3;
    wire beamXZ0Z_10;
    wire un1_beamxlt10_0_cascade_;
    wire HSync_c;
    wire beamXZ0Z_7;
    wire beamXZ0Z_6;
    wire un18_beamylto9_2;
    wire beamXZ0Z_8;
    wire beamXZ0Z_9;
    wire un1_beamx_2;
    wire bfn_9_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_;
    wire bfn_9_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_0;
    wire bfn_9_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un68_sum;
    wire un1_beamY_if_generate_plus_mult1_un61_sum;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_0;
    wire bfn_9_4_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6;
    wire G_6_i_a4_0_0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0;
    wire un5_visibley_i;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0;
    wire beamYZ0Z_1;
    wire Pixel_1_RNOZ0Z_12;
    wire N_8_cascade_;
    wire N_11;
    wire un15_0_1_cascade_;
    wire Pixel_c;
    wire PixelClock_g;
    wire un13_beamy;
    wire un4_beamy_0;
    wire un18_beamylt10_0;
    wire Pixel_0_sqmuxa_0;
    wire Pixel_0_sqmuxa_3;
    wire un1_visiblex_24;
    wire un14lt10;
    wire un1_visiblex_27;
    wire bfn_11_6_0_;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum;
    wire bfn_11_7_0_;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4;
    wire un5_visiblex_cry_8_c_RNI1D62Z0Z_0;
    wire CONSTANT_ONE_NET;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un40_sum_c5;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_i_8;
    wire un5_visiblex_cry_7_c_RNIVZ0Z952;
    wire un5_visiblex_i_24;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum;
    wire bfn_12_4_0_;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4;
    wire Pixel_1_RNOZ0Z_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum;
    wire bfn_12_5_0_;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6;
    wire bfn_12_6_0_;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__2237),
            .RESETB(N__4336),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__4866),
            .DIN(N__4865),
            .DOUT(N__4864),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__4866),
            .PADOUT(N__4865),
            .PADIN(N__4864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4082),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__4857),
            .DIN(N__4856),
            .DOUT(N__4855),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__4857),
            .PADOUT(N__4856),
            .PADIN(N__4855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__4848),
            .DIN(N__4847),
            .DOUT(N__4846),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__4848),
            .PADOUT(N__4847),
            .PADIN(N__4846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__4839),
            .DIN(N__4838),
            .DOUT(N__4837),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__4839),
            .PADOUT(N__4838),
            .PADIN(N__4837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4069),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__4830),
            .DIN(N__4829),
            .DOUT(N__4828),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__4830),
            .PADOUT(N__4829),
            .PADIN(N__4828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2831),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__4821),
            .DIN(N__4820),
            .DOUT(N__4819),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__4821),
            .PADOUT(N__4820),
            .PADIN(N__4819),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__4812),
            .DIN(N__4811),
            .DOUT(N__4810),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__4812),
            .PADOUT(N__4811),
            .PADIN(N__4810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1051 (
            .O(N__4793),
            .I(N__4790));
    LocalMux I__1050 (
            .O(N__4790),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__1049 (
            .O(N__4787),
            .I(N__4784));
    InMux I__1048 (
            .O(N__4784),
            .I(N__4781));
    LocalMux I__1047 (
            .O(N__4781),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i));
    CascadeMux I__1046 (
            .O(N__4778),
            .I(N__4775));
    InMux I__1045 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__1044 (
            .O(N__4772),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1));
    InMux I__1043 (
            .O(N__4769),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__1042 (
            .O(N__4766),
            .I(N__4763));
    InMux I__1041 (
            .O(N__4763),
            .I(N__4760));
    LocalMux I__1040 (
            .O(N__4760),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0));
    CascadeMux I__1039 (
            .O(N__4757),
            .I(N__4754));
    InMux I__1038 (
            .O(N__4754),
            .I(N__4751));
    LocalMux I__1037 (
            .O(N__4751),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332));
    InMux I__1036 (
            .O(N__4748),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1035 (
            .O(N__4745),
            .I(N__4742));
    LocalMux I__1034 (
            .O(N__4742),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__1033 (
            .O(N__4739),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1032 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__1031 (
            .O(N__4733),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__1030 (
            .O(N__4730),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7));
    InMux I__1029 (
            .O(N__4727),
            .I(N__4723));
    InMux I__1028 (
            .O(N__4726),
            .I(N__4720));
    LocalMux I__1027 (
            .O(N__4723),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2));
    LocalMux I__1026 (
            .O(N__4720),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2));
    CascadeMux I__1025 (
            .O(N__4715),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_));
    InMux I__1024 (
            .O(N__4712),
            .I(N__4706));
    InMux I__1023 (
            .O(N__4711),
            .I(N__4706));
    LocalMux I__1022 (
            .O(N__4706),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__1021 (
            .O(N__4703),
            .I(N__4699));
    InMux I__1020 (
            .O(N__4702),
            .I(N__4694));
    InMux I__1019 (
            .O(N__4699),
            .I(N__4694));
    LocalMux I__1018 (
            .O(N__4694),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831));
    InMux I__1017 (
            .O(N__4691),
            .I(N__4686));
    InMux I__1016 (
            .O(N__4690),
            .I(N__4681));
    InMux I__1015 (
            .O(N__4689),
            .I(N__4681));
    LocalMux I__1014 (
            .O(N__4686),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31));
    LocalMux I__1013 (
            .O(N__4681),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31));
    InMux I__1012 (
            .O(N__4676),
            .I(N__4673));
    LocalMux I__1011 (
            .O(N__4673),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62));
    CascadeMux I__1010 (
            .O(N__4670),
            .I(N__4666));
    InMux I__1009 (
            .O(N__4669),
            .I(N__4661));
    InMux I__1008 (
            .O(N__4666),
            .I(N__4661));
    LocalMux I__1007 (
            .O(N__4661),
            .I(N__4658));
    Odrv12 I__1006 (
            .O(N__4658),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1005 (
            .O(N__4655),
            .I(N__4652));
    InMux I__1004 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__1003 (
            .O(N__4649),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i));
    InMux I__1002 (
            .O(N__4646),
            .I(N__4640));
    InMux I__1001 (
            .O(N__4645),
            .I(N__4640));
    LocalMux I__1000 (
            .O(N__4640),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__999 (
            .O(N__4637),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__998 (
            .O(N__4634),
            .I(N__4628));
    InMux I__997 (
            .O(N__4633),
            .I(N__4628));
    LocalMux I__996 (
            .O(N__4628),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0));
    CascadeMux I__995 (
            .O(N__4625),
            .I(N__4622));
    InMux I__994 (
            .O(N__4622),
            .I(N__4619));
    LocalMux I__993 (
            .O(N__4619),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i));
    InMux I__992 (
            .O(N__4616),
            .I(N__4612));
    InMux I__991 (
            .O(N__4615),
            .I(N__4609));
    LocalMux I__990 (
            .O(N__4612),
            .I(N__4606));
    LocalMux I__989 (
            .O(N__4609),
            .I(N__4603));
    Span4Mux_s3_h I__988 (
            .O(N__4606),
            .I(N__4600));
    Span4Mux_s3_h I__987 (
            .O(N__4603),
            .I(N__4597));
    Odrv4 I__986 (
            .O(N__4600),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    Odrv4 I__985 (
            .O(N__4597),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum));
    InMux I__984 (
            .O(N__4592),
            .I(N__4589));
    LocalMux I__983 (
            .O(N__4589),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03));
    InMux I__982 (
            .O(N__4586),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__981 (
            .O(N__4583),
            .I(N__4580));
    InMux I__980 (
            .O(N__4580),
            .I(N__4577));
    LocalMux I__979 (
            .O(N__4577),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4));
    InMux I__978 (
            .O(N__4574),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__977 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__976 (
            .O(N__4568),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__975 (
            .O(N__4565),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__974 (
            .O(N__4562),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__973 (
            .O(N__4559),
            .I(N__4555));
    InMux I__972 (
            .O(N__4558),
            .I(N__4551));
    InMux I__971 (
            .O(N__4555),
            .I(N__4546));
    InMux I__970 (
            .O(N__4554),
            .I(N__4546));
    LocalMux I__969 (
            .O(N__4551),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6));
    LocalMux I__968 (
            .O(N__4546),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6));
    InMux I__967 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__966 (
            .O(N__4538),
            .I(N__4534));
    InMux I__965 (
            .O(N__4537),
            .I(N__4531));
    Span4Mux_v I__964 (
            .O(N__4534),
            .I(N__4525));
    LocalMux I__963 (
            .O(N__4531),
            .I(N__4525));
    InMux I__962 (
            .O(N__4530),
            .I(N__4522));
    Odrv4 I__961 (
            .O(N__4525),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_c5));
    LocalMux I__960 (
            .O(N__4522),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_c5));
    CascadeMux I__959 (
            .O(N__4517),
            .I(N__4514));
    InMux I__958 (
            .O(N__4514),
            .I(N__4511));
    LocalMux I__957 (
            .O(N__4511),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO));
    InMux I__956 (
            .O(N__4508),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__955 (
            .O(N__4505),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__954 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__953 (
            .O(N__4499),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    CascadeMux I__952 (
            .O(N__4496),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_));
    InMux I__951 (
            .O(N__4493),
            .I(N__4489));
    InMux I__950 (
            .O(N__4492),
            .I(N__4486));
    LocalMux I__949 (
            .O(N__4489),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0));
    LocalMux I__948 (
            .O(N__4486),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0));
    CascadeMux I__947 (
            .O(N__4481),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_));
    InMux I__946 (
            .O(N__4478),
            .I(N__4475));
    LocalMux I__945 (
            .O(N__4475),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__944 (
            .O(N__4472),
            .I(N__4466));
    InMux I__943 (
            .O(N__4471),
            .I(N__4466));
    LocalMux I__942 (
            .O(N__4466),
            .I(N__4463));
    Odrv4 I__941 (
            .O(N__4463),
            .I(un5_visiblex_cry_7_c_RNIVZ0Z952));
    CascadeMux I__940 (
            .O(N__4460),
            .I(N__4457));
    InMux I__939 (
            .O(N__4457),
            .I(N__4454));
    LocalMux I__938 (
            .O(N__4454),
            .I(un5_visiblex_i_24));
    CascadeMux I__937 (
            .O(N__4451),
            .I(N__4447));
    InMux I__936 (
            .O(N__4450),
            .I(N__4443));
    InMux I__935 (
            .O(N__4447),
            .I(N__4440));
    InMux I__934 (
            .O(N__4446),
            .I(N__4437));
    LocalMux I__933 (
            .O(N__4443),
            .I(N__4432));
    LocalMux I__932 (
            .O(N__4440),
            .I(N__4432));
    LocalMux I__931 (
            .O(N__4437),
            .I(N__4429));
    Span4Mux_s3_h I__930 (
            .O(N__4432),
            .I(N__4426));
    Span4Mux_s3_h I__929 (
            .O(N__4429),
            .I(N__4423));
    Odrv4 I__928 (
            .O(N__4426),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    Odrv4 I__927 (
            .O(N__4423),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum));
    InMux I__926 (
            .O(N__4418),
            .I(N__4412));
    InMux I__925 (
            .O(N__4417),
            .I(N__4412));
    LocalMux I__924 (
            .O(N__4412),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5));
    InMux I__923 (
            .O(N__4409),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__922 (
            .O(N__4406),
            .I(N__4403));
    LocalMux I__921 (
            .O(N__4403),
            .I(Pixel_1_RNOZ0Z_8));
    InMux I__920 (
            .O(N__4400),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__919 (
            .O(N__4397),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__918 (
            .O(N__4394),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__917 (
            .O(N__4391),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__916 (
            .O(N__4388),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__915 (
            .O(N__4385),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_));
    InMux I__914 (
            .O(N__4382),
            .I(N__4376));
    InMux I__913 (
            .O(N__4381),
            .I(N__4376));
    LocalMux I__912 (
            .O(N__4376),
            .I(N__4373));
    Span4Mux_s1_h I__911 (
            .O(N__4373),
            .I(N__4370));
    Odrv4 I__910 (
            .O(N__4370),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum));
    InMux I__909 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__908 (
            .O(N__4364),
            .I(N__4361));
    Odrv4 I__907 (
            .O(N__4361),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i));
    CascadeMux I__906 (
            .O(N__4358),
            .I(N__4355));
    InMux I__905 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__904 (
            .O(N__4352),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0));
    InMux I__903 (
            .O(N__4349),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__902 (
            .O(N__4346),
            .I(N__4343));
    LocalMux I__901 (
            .O(N__4343),
            .I(N__4340));
    Odrv4 I__900 (
            .O(N__4340),
            .I(un5_visiblex_cry_8_c_RNI1D62Z0Z_0));
    CascadeMux I__899 (
            .O(N__4337),
            .I(N__4333));
    IoInMux I__898 (
            .O(N__4336),
            .I(N__4327));
    InMux I__897 (
            .O(N__4333),
            .I(N__4324));
    CascadeMux I__896 (
            .O(N__4332),
            .I(N__4321));
    CascadeMux I__895 (
            .O(N__4331),
            .I(N__4318));
    CascadeMux I__894 (
            .O(N__4330),
            .I(N__4315));
    LocalMux I__893 (
            .O(N__4327),
            .I(N__4312));
    LocalMux I__892 (
            .O(N__4324),
            .I(N__4309));
    InMux I__891 (
            .O(N__4321),
            .I(N__4306));
    InMux I__890 (
            .O(N__4318),
            .I(N__4303));
    InMux I__889 (
            .O(N__4315),
            .I(N__4300));
    Span4Mux_s1_v I__888 (
            .O(N__4312),
            .I(N__4291));
    Span4Mux_v I__887 (
            .O(N__4309),
            .I(N__4286));
    LocalMux I__886 (
            .O(N__4306),
            .I(N__4279));
    LocalMux I__885 (
            .O(N__4303),
            .I(N__4279));
    LocalMux I__884 (
            .O(N__4300),
            .I(N__4279));
    InMux I__883 (
            .O(N__4299),
            .I(N__4276));
    InMux I__882 (
            .O(N__4298),
            .I(N__4271));
    InMux I__881 (
            .O(N__4297),
            .I(N__4271));
    CascadeMux I__880 (
            .O(N__4296),
            .I(N__4268));
    CascadeMux I__879 (
            .O(N__4295),
            .I(N__4265));
    CascadeMux I__878 (
            .O(N__4294),
            .I(N__4262));
    Span4Mux_h I__877 (
            .O(N__4291),
            .I(N__4257));
    InMux I__876 (
            .O(N__4290),
            .I(N__4252));
    InMux I__875 (
            .O(N__4289),
            .I(N__4252));
    Span4Mux_h I__874 (
            .O(N__4286),
            .I(N__4243));
    Span4Mux_v I__873 (
            .O(N__4279),
            .I(N__4243));
    LocalMux I__872 (
            .O(N__4276),
            .I(N__4243));
    LocalMux I__871 (
            .O(N__4271),
            .I(N__4243));
    InMux I__870 (
            .O(N__4268),
            .I(N__4240));
    InMux I__869 (
            .O(N__4265),
            .I(N__4235));
    InMux I__868 (
            .O(N__4262),
            .I(N__4235));
    InMux I__867 (
            .O(N__4261),
            .I(N__4232));
    InMux I__866 (
            .O(N__4260),
            .I(N__4229));
    Odrv4 I__865 (
            .O(N__4257),
            .I(CONSTANT_ONE_NET));
    LocalMux I__864 (
            .O(N__4252),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__863 (
            .O(N__4243),
            .I(CONSTANT_ONE_NET));
    LocalMux I__862 (
            .O(N__4240),
            .I(CONSTANT_ONE_NET));
    LocalMux I__861 (
            .O(N__4235),
            .I(CONSTANT_ONE_NET));
    LocalMux I__860 (
            .O(N__4232),
            .I(CONSTANT_ONE_NET));
    LocalMux I__859 (
            .O(N__4229),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__858 (
            .O(N__4214),
            .I(N__4211));
    InMux I__857 (
            .O(N__4211),
            .I(N__4208));
    LocalMux I__856 (
            .O(N__4208),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0));
    InMux I__855 (
            .O(N__4205),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__854 (
            .O(N__4202),
            .I(N__4198));
    InMux I__853 (
            .O(N__4201),
            .I(N__4195));
    LocalMux I__852 (
            .O(N__4198),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59));
    LocalMux I__851 (
            .O(N__4195),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59));
    InMux I__850 (
            .O(N__4190),
            .I(N__4186));
    InMux I__849 (
            .O(N__4189),
            .I(N__4183));
    LocalMux I__848 (
            .O(N__4186),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0));
    LocalMux I__847 (
            .O(N__4183),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0));
    CascadeMux I__846 (
            .O(N__4178),
            .I(N__4174));
    InMux I__845 (
            .O(N__4177),
            .I(N__4170));
    InMux I__844 (
            .O(N__4174),
            .I(N__4167));
    InMux I__843 (
            .O(N__4173),
            .I(N__4164));
    LocalMux I__842 (
            .O(N__4170),
            .I(un5_visibley_i));
    LocalMux I__841 (
            .O(N__4167),
            .I(un5_visibley_i));
    LocalMux I__840 (
            .O(N__4164),
            .I(un5_visibley_i));
    InMux I__839 (
            .O(N__4157),
            .I(N__4154));
    LocalMux I__838 (
            .O(N__4154),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0));
    CascadeMux I__837 (
            .O(N__4151),
            .I(N__4147));
    InMux I__836 (
            .O(N__4150),
            .I(N__4142));
    InMux I__835 (
            .O(N__4147),
            .I(N__4138));
    InMux I__834 (
            .O(N__4146),
            .I(N__4135));
    InMux I__833 (
            .O(N__4145),
            .I(N__4132));
    LocalMux I__832 (
            .O(N__4142),
            .I(N__4129));
    InMux I__831 (
            .O(N__4141),
            .I(N__4125));
    LocalMux I__830 (
            .O(N__4138),
            .I(N__4118));
    LocalMux I__829 (
            .O(N__4135),
            .I(N__4118));
    LocalMux I__828 (
            .O(N__4132),
            .I(N__4118));
    Span4Mux_v I__827 (
            .O(N__4129),
            .I(N__4115));
    InMux I__826 (
            .O(N__4128),
            .I(N__4112));
    LocalMux I__825 (
            .O(N__4125),
            .I(N__4107));
    Span4Mux_h I__824 (
            .O(N__4118),
            .I(N__4107));
    Odrv4 I__823 (
            .O(N__4115),
            .I(beamYZ0Z_1));
    LocalMux I__822 (
            .O(N__4112),
            .I(beamYZ0Z_1));
    Odrv4 I__821 (
            .O(N__4107),
            .I(beamYZ0Z_1));
    InMux I__820 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__819 (
            .O(N__4097),
            .I(Pixel_1_RNOZ0Z_12));
    CascadeMux I__818 (
            .O(N__4094),
            .I(N_8_cascade_));
    InMux I__817 (
            .O(N__4091),
            .I(N__4088));
    LocalMux I__816 (
            .O(N__4088),
            .I(N_11));
    CascadeMux I__815 (
            .O(N__4085),
            .I(un15_0_1_cascade_));
    IoInMux I__814 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__813 (
            .O(N__4079),
            .I(N__4076));
    IoSpan4Mux I__812 (
            .O(N__4076),
            .I(N__4073));
    Span4Mux_s3_h I__811 (
            .O(N__4073),
            .I(N__4070));
    Span4Mux_v I__810 (
            .O(N__4070),
            .I(N__4066));
    IoInMux I__809 (
            .O(N__4069),
            .I(N__4063));
    Sp12to4 I__808 (
            .O(N__4066),
            .I(N__4058));
    LocalMux I__807 (
            .O(N__4063),
            .I(N__4058));
    Odrv12 I__806 (
            .O(N__4058),
            .I(Pixel_c));
    ClkMux I__805 (
            .O(N__4055),
            .I(N__4025));
    ClkMux I__804 (
            .O(N__4054),
            .I(N__4025));
    ClkMux I__803 (
            .O(N__4053),
            .I(N__4025));
    ClkMux I__802 (
            .O(N__4052),
            .I(N__4025));
    ClkMux I__801 (
            .O(N__4051),
            .I(N__4025));
    ClkMux I__800 (
            .O(N__4050),
            .I(N__4025));
    ClkMux I__799 (
            .O(N__4049),
            .I(N__4025));
    ClkMux I__798 (
            .O(N__4048),
            .I(N__4025));
    ClkMux I__797 (
            .O(N__4047),
            .I(N__4025));
    ClkMux I__796 (
            .O(N__4046),
            .I(N__4025));
    GlobalMux I__795 (
            .O(N__4025),
            .I(N__4022));
    gio2CtrlBuf I__794 (
            .O(N__4022),
            .I(PixelClock_g));
    InMux I__793 (
            .O(N__4019),
            .I(N__4016));
    LocalMux I__792 (
            .O(N__4016),
            .I(un13_beamy));
    InMux I__791 (
            .O(N__4013),
            .I(N__4010));
    LocalMux I__790 (
            .O(N__4010),
            .I(un4_beamy_0));
    CascadeMux I__789 (
            .O(N__4007),
            .I(N__4004));
    InMux I__788 (
            .O(N__4004),
            .I(N__4001));
    LocalMux I__787 (
            .O(N__4001),
            .I(N__3998));
    Odrv4 I__786 (
            .O(N__3998),
            .I(un18_beamylt10_0));
    InMux I__785 (
            .O(N__3995),
            .I(N__3992));
    LocalMux I__784 (
            .O(N__3992),
            .I(N__3989));
    Odrv4 I__783 (
            .O(N__3989),
            .I(Pixel_0_sqmuxa_0));
    InMux I__782 (
            .O(N__3986),
            .I(N__3983));
    LocalMux I__781 (
            .O(N__3983),
            .I(Pixel_0_sqmuxa_3));
    CascadeMux I__780 (
            .O(N__3980),
            .I(N__3977));
    InMux I__779 (
            .O(N__3977),
            .I(N__3974));
    LocalMux I__778 (
            .O(N__3974),
            .I(N__3971));
    Span4Mux_s3_h I__777 (
            .O(N__3971),
            .I(N__3968));
    Odrv4 I__776 (
            .O(N__3968),
            .I(un1_visiblex_24));
    InMux I__775 (
            .O(N__3965),
            .I(N__3962));
    LocalMux I__774 (
            .O(N__3962),
            .I(N__3959));
    Odrv12 I__773 (
            .O(N__3959),
            .I(un14lt10));
    InMux I__772 (
            .O(N__3956),
            .I(N__3953));
    LocalMux I__771 (
            .O(N__3953),
            .I(N__3950));
    Odrv4 I__770 (
            .O(N__3950),
            .I(un1_visiblex_27));
    InMux I__769 (
            .O(N__3947),
            .I(N__3943));
    InMux I__768 (
            .O(N__3946),
            .I(N__3940));
    LocalMux I__767 (
            .O(N__3943),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    LocalMux I__766 (
            .O(N__3940),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    CascadeMux I__765 (
            .O(N__3935),
            .I(N__3932));
    InMux I__764 (
            .O(N__3932),
            .I(N__3929));
    LocalMux I__763 (
            .O(N__3929),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__762 (
            .O(N__3926),
            .I(N__3923));
    LocalMux I__761 (
            .O(N__3923),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__760 (
            .O(N__3920),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__759 (
            .O(N__3917),
            .I(N__3914));
    InMux I__758 (
            .O(N__3914),
            .I(N__3911));
    LocalMux I__757 (
            .O(N__3911),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4));
    InMux I__756 (
            .O(N__3908),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__755 (
            .O(N__3905),
            .I(N__3902));
    LocalMux I__754 (
            .O(N__3902),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7));
    InMux I__753 (
            .O(N__3899),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__752 (
            .O(N__3896),
            .I(N__3893));
    LocalMux I__751 (
            .O(N__3893),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7));
    CascadeMux I__750 (
            .O(N__3890),
            .I(N__3885));
    CascadeMux I__749 (
            .O(N__3889),
            .I(N__3881));
    InMux I__748 (
            .O(N__3888),
            .I(N__3877));
    InMux I__747 (
            .O(N__3885),
            .I(N__3868));
    InMux I__746 (
            .O(N__3884),
            .I(N__3868));
    InMux I__745 (
            .O(N__3881),
            .I(N__3868));
    InMux I__744 (
            .O(N__3880),
            .I(N__3868));
    LocalMux I__743 (
            .O(N__3877),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8));
    LocalMux I__742 (
            .O(N__3868),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8));
    CascadeMux I__741 (
            .O(N__3863),
            .I(N__3860));
    InMux I__740 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__739 (
            .O(N__3857),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__738 (
            .O(N__3854),
            .I(N__3851));
    LocalMux I__737 (
            .O(N__3851),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__736 (
            .O(N__3848),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__735 (
            .O(N__3845),
            .I(N__3842));
    LocalMux I__734 (
            .O(N__3842),
            .I(G_6_i_a4_0_0));
    CascadeMux I__733 (
            .O(N__3839),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_));
    CascadeMux I__732 (
            .O(N__3836),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_));
    InMux I__731 (
            .O(N__3833),
            .I(N__3829));
    InMux I__730 (
            .O(N__3832),
            .I(N__3826));
    LocalMux I__729 (
            .O(N__3829),
            .I(N__3823));
    LocalMux I__728 (
            .O(N__3826),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    Odrv4 I__727 (
            .O(N__3823),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    CascadeMux I__726 (
            .O(N__3818),
            .I(N__3815));
    InMux I__725 (
            .O(N__3815),
            .I(N__3812));
    LocalMux I__724 (
            .O(N__3812),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__723 (
            .O(N__3809),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__722 (
            .O(N__3806),
            .I(N__3803));
    LocalMux I__721 (
            .O(N__3803),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2));
    InMux I__720 (
            .O(N__3800),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__719 (
            .O(N__3797),
            .I(N__3793));
    InMux I__718 (
            .O(N__3796),
            .I(N__3784));
    InMux I__717 (
            .O(N__3793),
            .I(N__3784));
    InMux I__716 (
            .O(N__3792),
            .I(N__3784));
    InMux I__715 (
            .O(N__3791),
            .I(N__3781));
    LocalMux I__714 (
            .O(N__3784),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4));
    LocalMux I__713 (
            .O(N__3781),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4));
    CascadeMux I__712 (
            .O(N__3776),
            .I(N__3773));
    InMux I__711 (
            .O(N__3773),
            .I(N__3770));
    LocalMux I__710 (
            .O(N__3770),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3));
    InMux I__709 (
            .O(N__3767),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__708 (
            .O(N__3764),
            .I(N__3761));
    LocalMux I__707 (
            .O(N__3761),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3));
    CascadeMux I__706 (
            .O(N__3758),
            .I(N__3755));
    InMux I__705 (
            .O(N__3755),
            .I(N__3752));
    LocalMux I__704 (
            .O(N__3752),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__703 (
            .O(N__3749),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__702 (
            .O(N__3746),
            .I(N__3743));
    LocalMux I__701 (
            .O(N__3743),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__700 (
            .O(N__3740),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__699 (
            .O(N__3737),
            .I(N__3733));
    InMux I__698 (
            .O(N__3736),
            .I(N__3728));
    InMux I__697 (
            .O(N__3733),
            .I(N__3728));
    LocalMux I__696 (
            .O(N__3728),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    InMux I__695 (
            .O(N__3725),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__694 (
            .O(N__3722),
            .I(N__3719));
    LocalMux I__693 (
            .O(N__3719),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__692 (
            .O(N__3716),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__691 (
            .O(N__3713),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_));
    InMux I__690 (
            .O(N__3710),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__689 (
            .O(N__3707),
            .I(N__3704));
    LocalMux I__688 (
            .O(N__3704),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0));
    InMux I__687 (
            .O(N__3701),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__686 (
            .O(N__3698),
            .I(N__3694));
    InMux I__685 (
            .O(N__3697),
            .I(N__3685));
    InMux I__684 (
            .O(N__3694),
            .I(N__3685));
    InMux I__683 (
            .O(N__3693),
            .I(N__3685));
    InMux I__682 (
            .O(N__3692),
            .I(N__3682));
    LocalMux I__681 (
            .O(N__3685),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02));
    LocalMux I__680 (
            .O(N__3682),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02));
    CascadeMux I__679 (
            .O(N__3677),
            .I(N__3674));
    InMux I__678 (
            .O(N__3674),
            .I(N__3671));
    LocalMux I__677 (
            .O(N__3671),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1));
    InMux I__676 (
            .O(N__3668),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__675 (
            .O(N__3665),
            .I(N__3662));
    LocalMux I__674 (
            .O(N__3662),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1));
    CascadeMux I__673 (
            .O(N__3659),
            .I(N__3656));
    InMux I__672 (
            .O(N__3656),
            .I(N__3653));
    LocalMux I__671 (
            .O(N__3653),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__670 (
            .O(N__3650),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__669 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__668 (
            .O(N__3644),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__667 (
            .O(N__3641),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__666 (
            .O(N__3638),
            .I(N__3635));
    InMux I__665 (
            .O(N__3635),
            .I(N__3628));
    InMux I__664 (
            .O(N__3634),
            .I(N__3623));
    InMux I__663 (
            .O(N__3633),
            .I(N__3623));
    InMux I__662 (
            .O(N__3632),
            .I(N__3619));
    InMux I__661 (
            .O(N__3631),
            .I(N__3616));
    LocalMux I__660 (
            .O(N__3628),
            .I(N__3613));
    LocalMux I__659 (
            .O(N__3623),
            .I(N__3610));
    InMux I__658 (
            .O(N__3622),
            .I(N__3607));
    LocalMux I__657 (
            .O(N__3619),
            .I(beamXZ0Z_5));
    LocalMux I__656 (
            .O(N__3616),
            .I(beamXZ0Z_5));
    Odrv4 I__655 (
            .O(N__3613),
            .I(beamXZ0Z_5));
    Odrv4 I__654 (
            .O(N__3610),
            .I(beamXZ0Z_5));
    LocalMux I__653 (
            .O(N__3607),
            .I(beamXZ0Z_5));
    InMux I__652 (
            .O(N__3596),
            .I(N__3589));
    InMux I__651 (
            .O(N__3595),
            .I(N__3584));
    InMux I__650 (
            .O(N__3594),
            .I(N__3584));
    InMux I__649 (
            .O(N__3593),
            .I(N__3580));
    InMux I__648 (
            .O(N__3592),
            .I(N__3577));
    LocalMux I__647 (
            .O(N__3589),
            .I(N__3574));
    LocalMux I__646 (
            .O(N__3584),
            .I(N__3571));
    InMux I__645 (
            .O(N__3583),
            .I(N__3568));
    LocalMux I__644 (
            .O(N__3580),
            .I(beamXZ0Z_4));
    LocalMux I__643 (
            .O(N__3577),
            .I(beamXZ0Z_4));
    Odrv4 I__642 (
            .O(N__3574),
            .I(beamXZ0Z_4));
    Odrv4 I__641 (
            .O(N__3571),
            .I(beamXZ0Z_4));
    LocalMux I__640 (
            .O(N__3568),
            .I(beamXZ0Z_4));
    CascadeMux I__639 (
            .O(N__3557),
            .I(N__3553));
    InMux I__638 (
            .O(N__3556),
            .I(N__3548));
    InMux I__637 (
            .O(N__3553),
            .I(N__3545));
    InMux I__636 (
            .O(N__3552),
            .I(N__3541));
    InMux I__635 (
            .O(N__3551),
            .I(N__3538));
    LocalMux I__634 (
            .O(N__3548),
            .I(N__3533));
    LocalMux I__633 (
            .O(N__3545),
            .I(N__3533));
    InMux I__632 (
            .O(N__3544),
            .I(N__3530));
    LocalMux I__631 (
            .O(N__3541),
            .I(beamXZ0Z_3));
    LocalMux I__630 (
            .O(N__3538),
            .I(beamXZ0Z_3));
    Odrv4 I__629 (
            .O(N__3533),
            .I(beamXZ0Z_3));
    LocalMux I__628 (
            .O(N__3530),
            .I(beamXZ0Z_3));
    CascadeMux I__627 (
            .O(N__3521),
            .I(N__3516));
    InMux I__626 (
            .O(N__3520),
            .I(N__3511));
    InMux I__625 (
            .O(N__3519),
            .I(N__3511));
    InMux I__624 (
            .O(N__3516),
            .I(N__3508));
    LocalMux I__623 (
            .O(N__3511),
            .I(N__3501));
    LocalMux I__622 (
            .O(N__3508),
            .I(N__3501));
    InMux I__621 (
            .O(N__3507),
            .I(N__3498));
    InMux I__620 (
            .O(N__3506),
            .I(N__3495));
    Span4Mux_h I__619 (
            .O(N__3501),
            .I(N__3492));
    LocalMux I__618 (
            .O(N__3498),
            .I(beamXZ0Z_10));
    LocalMux I__617 (
            .O(N__3495),
            .I(beamXZ0Z_10));
    Odrv4 I__616 (
            .O(N__3492),
            .I(beamXZ0Z_10));
    CascadeMux I__615 (
            .O(N__3485),
            .I(un1_beamxlt10_0_cascade_));
    IoInMux I__614 (
            .O(N__3482),
            .I(N__3478));
    IoInMux I__613 (
            .O(N__3481),
            .I(N__3475));
    LocalMux I__612 (
            .O(N__3478),
            .I(N__3472));
    LocalMux I__611 (
            .O(N__3475),
            .I(N__3469));
    Span12Mux_s9_v I__610 (
            .O(N__3472),
            .I(N__3466));
    Span4Mux_s2_v I__609 (
            .O(N__3469),
            .I(N__3463));
    Odrv12 I__608 (
            .O(N__3466),
            .I(HSync_c));
    Odrv4 I__607 (
            .O(N__3463),
            .I(HSync_c));
    InMux I__606 (
            .O(N__3458),
            .I(N__3454));
    InMux I__605 (
            .O(N__3457),
            .I(N__3450));
    LocalMux I__604 (
            .O(N__3454),
            .I(N__3444));
    InMux I__603 (
            .O(N__3453),
            .I(N__3441));
    LocalMux I__602 (
            .O(N__3450),
            .I(N__3438));
    InMux I__601 (
            .O(N__3449),
            .I(N__3433));
    InMux I__600 (
            .O(N__3448),
            .I(N__3433));
    InMux I__599 (
            .O(N__3447),
            .I(N__3430));
    Odrv4 I__598 (
            .O(N__3444),
            .I(beamXZ0Z_7));
    LocalMux I__597 (
            .O(N__3441),
            .I(beamXZ0Z_7));
    Odrv4 I__596 (
            .O(N__3438),
            .I(beamXZ0Z_7));
    LocalMux I__595 (
            .O(N__3433),
            .I(beamXZ0Z_7));
    LocalMux I__594 (
            .O(N__3430),
            .I(beamXZ0Z_7));
    InMux I__593 (
            .O(N__3419),
            .I(N__3415));
    InMux I__592 (
            .O(N__3418),
            .I(N__3412));
    LocalMux I__591 (
            .O(N__3415),
            .I(N__3405));
    LocalMux I__590 (
            .O(N__3412),
            .I(N__3405));
    CascadeMux I__589 (
            .O(N__3411),
            .I(N__3402));
    InMux I__588 (
            .O(N__3410),
            .I(N__3397));
    Span4Mux_h I__587 (
            .O(N__3405),
            .I(N__3394));
    InMux I__586 (
            .O(N__3402),
            .I(N__3389));
    InMux I__585 (
            .O(N__3401),
            .I(N__3389));
    InMux I__584 (
            .O(N__3400),
            .I(N__3386));
    LocalMux I__583 (
            .O(N__3397),
            .I(beamXZ0Z_6));
    Odrv4 I__582 (
            .O(N__3394),
            .I(beamXZ0Z_6));
    LocalMux I__581 (
            .O(N__3389),
            .I(beamXZ0Z_6));
    LocalMux I__580 (
            .O(N__3386),
            .I(beamXZ0Z_6));
    CascadeMux I__579 (
            .O(N__3377),
            .I(N__3374));
    InMux I__578 (
            .O(N__3374),
            .I(N__3371));
    LocalMux I__577 (
            .O(N__3371),
            .I(N__3368));
    Odrv4 I__576 (
            .O(N__3368),
            .I(un18_beamylto9_2));
    InMux I__575 (
            .O(N__3365),
            .I(N__3359));
    InMux I__574 (
            .O(N__3364),
            .I(N__3356));
    InMux I__573 (
            .O(N__3363),
            .I(N__3351));
    InMux I__572 (
            .O(N__3362),
            .I(N__3351));
    LocalMux I__571 (
            .O(N__3359),
            .I(beamXZ0Z_8));
    LocalMux I__570 (
            .O(N__3356),
            .I(beamXZ0Z_8));
    LocalMux I__569 (
            .O(N__3351),
            .I(beamXZ0Z_8));
    CascadeMux I__568 (
            .O(N__3344),
            .I(N__3340));
    InMux I__567 (
            .O(N__3343),
            .I(N__3335));
    InMux I__566 (
            .O(N__3340),
            .I(N__3328));
    InMux I__565 (
            .O(N__3339),
            .I(N__3328));
    InMux I__564 (
            .O(N__3338),
            .I(N__3328));
    LocalMux I__563 (
            .O(N__3335),
            .I(beamXZ0Z_9));
    LocalMux I__562 (
            .O(N__3328),
            .I(beamXZ0Z_9));
    InMux I__561 (
            .O(N__3323),
            .I(N__3318));
    InMux I__560 (
            .O(N__3322),
            .I(N__3315));
    InMux I__559 (
            .O(N__3321),
            .I(N__3312));
    LocalMux I__558 (
            .O(N__3318),
            .I(N__3307));
    LocalMux I__557 (
            .O(N__3315),
            .I(N__3307));
    LocalMux I__556 (
            .O(N__3312),
            .I(un1_beamx_2));
    Odrv4 I__555 (
            .O(N__3307),
            .I(un1_beamx_2));
    CascadeMux I__554 (
            .O(N__3302),
            .I(N__3299));
    InMux I__553 (
            .O(N__3299),
            .I(N__3296));
    LocalMux I__552 (
            .O(N__3296),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__551 (
            .O(N__3293),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__550 (
            .O(N__3290),
            .I(N__3287));
    LocalMux I__549 (
            .O(N__3287),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0));
    InMux I__548 (
            .O(N__3284),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__547 (
            .O(N__3281),
            .I(N__3277));
    InMux I__546 (
            .O(N__3280),
            .I(N__3268));
    InMux I__545 (
            .O(N__3277),
            .I(N__3268));
    InMux I__544 (
            .O(N__3276),
            .I(N__3268));
    InMux I__543 (
            .O(N__3275),
            .I(N__3265));
    LocalMux I__542 (
            .O(N__3268),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    LocalMux I__541 (
            .O(N__3265),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    CascadeMux I__540 (
            .O(N__3260),
            .I(N__3257));
    InMux I__539 (
            .O(N__3257),
            .I(N__3254));
    LocalMux I__538 (
            .O(N__3254),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0));
    InMux I__537 (
            .O(N__3251),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__536 (
            .O(N__3248),
            .I(N__3245));
    LocalMux I__535 (
            .O(N__3245),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61));
    CascadeMux I__534 (
            .O(N__3242),
            .I(N__3239));
    InMux I__533 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__532 (
            .O(N__3236),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_7));
    InMux I__531 (
            .O(N__3233),
            .I(N__3227));
    InMux I__530 (
            .O(N__3232),
            .I(N__3224));
    InMux I__529 (
            .O(N__3231),
            .I(N__3221));
    InMux I__528 (
            .O(N__3230),
            .I(N__3218));
    LocalMux I__527 (
            .O(N__3227),
            .I(N__3213));
    LocalMux I__526 (
            .O(N__3224),
            .I(N__3213));
    LocalMux I__525 (
            .O(N__3221),
            .I(N__3210));
    LocalMux I__524 (
            .O(N__3218),
            .I(beamXZ0Z_2));
    Odrv4 I__523 (
            .O(N__3213),
            .I(beamXZ0Z_2));
    Odrv4 I__522 (
            .O(N__3210),
            .I(beamXZ0Z_2));
    InMux I__521 (
            .O(N__3203),
            .I(un5_visiblex_cry_2));
    InMux I__520 (
            .O(N__3200),
            .I(un5_visiblex_cry_3));
    InMux I__519 (
            .O(N__3197),
            .I(un5_visiblex_cry_4));
    InMux I__518 (
            .O(N__3194),
            .I(un5_visiblex_cry_5));
    InMux I__517 (
            .O(N__3191),
            .I(un5_visiblex_cry_6));
    InMux I__516 (
            .O(N__3188),
            .I(bfn_8_7_0_));
    InMux I__515 (
            .O(N__3185),
            .I(un5_visiblex_cry_8));
    CascadeMux I__514 (
            .O(N__3182),
            .I(un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_));
    InMux I__513 (
            .O(N__3179),
            .I(N__3176));
    LocalMux I__512 (
            .O(N__3176),
            .I(un18_beamylt4));
    CascadeMux I__511 (
            .O(N__3173),
            .I(un18_beamylt4_cascade_));
    CascadeMux I__510 (
            .O(N__3170),
            .I(un13_beamylt7_cascade_));
    InMux I__509 (
            .O(N__3167),
            .I(N__3164));
    LocalMux I__508 (
            .O(N__3164),
            .I(N__3160));
    InMux I__507 (
            .O(N__3163),
            .I(N__3157));
    Odrv4 I__506 (
            .O(N__3160),
            .I(un8_beamy_2));
    LocalMux I__505 (
            .O(N__3157),
            .I(un8_beamy_2));
    CascadeMux I__504 (
            .O(N__3152),
            .I(N__3147));
    InMux I__503 (
            .O(N__3151),
            .I(N__3144));
    InMux I__502 (
            .O(N__3150),
            .I(N__3141));
    InMux I__501 (
            .O(N__3147),
            .I(N__3138));
    LocalMux I__500 (
            .O(N__3144),
            .I(N__3135));
    LocalMux I__499 (
            .O(N__3141),
            .I(un1_beamy_4));
    LocalMux I__498 (
            .O(N__3138),
            .I(un1_beamy_4));
    Odrv4 I__497 (
            .O(N__3135),
            .I(un1_beamy_4));
    InMux I__496 (
            .O(N__3128),
            .I(N__3124));
    InMux I__495 (
            .O(N__3127),
            .I(N__3121));
    LocalMux I__494 (
            .O(N__3124),
            .I(N__3112));
    LocalMux I__493 (
            .O(N__3121),
            .I(N__3112));
    CascadeMux I__492 (
            .O(N__3120),
            .I(N__3109));
    InMux I__491 (
            .O(N__3119),
            .I(N__3106));
    InMux I__490 (
            .O(N__3118),
            .I(N__3103));
    InMux I__489 (
            .O(N__3117),
            .I(N__3100));
    Span4Mux_v I__488 (
            .O(N__3112),
            .I(N__3097));
    InMux I__487 (
            .O(N__3109),
            .I(N__3094));
    LocalMux I__486 (
            .O(N__3106),
            .I(beamYZ0Z_7));
    LocalMux I__485 (
            .O(N__3103),
            .I(beamYZ0Z_7));
    LocalMux I__484 (
            .O(N__3100),
            .I(beamYZ0Z_7));
    Odrv4 I__483 (
            .O(N__3097),
            .I(beamYZ0Z_7));
    LocalMux I__482 (
            .O(N__3094),
            .I(beamYZ0Z_7));
    InMux I__481 (
            .O(N__3083),
            .I(N__3073));
    InMux I__480 (
            .O(N__3082),
            .I(N__3073));
    InMux I__479 (
            .O(N__3081),
            .I(N__3063));
    InMux I__478 (
            .O(N__3080),
            .I(N__3063));
    InMux I__477 (
            .O(N__3079),
            .I(N__3063));
    InMux I__476 (
            .O(N__3078),
            .I(N__3063));
    LocalMux I__475 (
            .O(N__3073),
            .I(N__3060));
    InMux I__474 (
            .O(N__3072),
            .I(N__3057));
    LocalMux I__473 (
            .O(N__3063),
            .I(un5_beamx_3));
    Odrv4 I__472 (
            .O(N__3060),
            .I(un5_beamx_3));
    LocalMux I__471 (
            .O(N__3057),
            .I(un5_beamx_3));
    CascadeMux I__470 (
            .O(N__3050),
            .I(un8_beamylto9_1_cascade_));
    CascadeMux I__469 (
            .O(N__3047),
            .I(N__3043));
    CascadeMux I__468 (
            .O(N__3046),
            .I(N__3035));
    InMux I__467 (
            .O(N__3043),
            .I(N__3032));
    InMux I__466 (
            .O(N__3042),
            .I(N__3029));
    InMux I__465 (
            .O(N__3041),
            .I(N__3026));
    InMux I__464 (
            .O(N__3040),
            .I(N__3019));
    InMux I__463 (
            .O(N__3039),
            .I(N__3019));
    InMux I__462 (
            .O(N__3038),
            .I(N__3019));
    InMux I__461 (
            .O(N__3035),
            .I(N__3016));
    LocalMux I__460 (
            .O(N__3032),
            .I(beamYZ0Z_2));
    LocalMux I__459 (
            .O(N__3029),
            .I(beamYZ0Z_2));
    LocalMux I__458 (
            .O(N__3026),
            .I(beamYZ0Z_2));
    LocalMux I__457 (
            .O(N__3019),
            .I(beamYZ0Z_2));
    LocalMux I__456 (
            .O(N__3016),
            .I(beamYZ0Z_2));
    InMux I__455 (
            .O(N__3005),
            .I(N__3002));
    LocalMux I__454 (
            .O(N__3002),
            .I(N__2994));
    InMux I__453 (
            .O(N__3001),
            .I(N__2989));
    InMux I__452 (
            .O(N__3000),
            .I(N__2989));
    InMux I__451 (
            .O(N__2999),
            .I(N__2986));
    InMux I__450 (
            .O(N__2998),
            .I(N__2981));
    InMux I__449 (
            .O(N__2997),
            .I(N__2981));
    Odrv4 I__448 (
            .O(N__2994),
            .I(beamXZ0Z_0));
    LocalMux I__447 (
            .O(N__2989),
            .I(beamXZ0Z_0));
    LocalMux I__446 (
            .O(N__2986),
            .I(beamXZ0Z_0));
    LocalMux I__445 (
            .O(N__2981),
            .I(beamXZ0Z_0));
    CascadeMux I__444 (
            .O(N__2972),
            .I(N__2969));
    InMux I__443 (
            .O(N__2969),
            .I(N__2963));
    InMux I__442 (
            .O(N__2968),
            .I(N__2960));
    InMux I__441 (
            .O(N__2967),
            .I(N__2957));
    InMux I__440 (
            .O(N__2966),
            .I(N__2954));
    LocalMux I__439 (
            .O(N__2963),
            .I(beamXZ0Z_1));
    LocalMux I__438 (
            .O(N__2960),
            .I(beamXZ0Z_1));
    LocalMux I__437 (
            .O(N__2957),
            .I(beamXZ0Z_1));
    LocalMux I__436 (
            .O(N__2954),
            .I(beamXZ0Z_1));
    CascadeMux I__435 (
            .O(N__2945),
            .I(N__2939));
    InMux I__434 (
            .O(N__2944),
            .I(N__2936));
    InMux I__433 (
            .O(N__2943),
            .I(N__2933));
    InMux I__432 (
            .O(N__2942),
            .I(N__2930));
    InMux I__431 (
            .O(N__2939),
            .I(N__2927));
    LocalMux I__430 (
            .O(N__2936),
            .I(beamYZ0Z_6));
    LocalMux I__429 (
            .O(N__2933),
            .I(beamYZ0Z_6));
    LocalMux I__428 (
            .O(N__2930),
            .I(beamYZ0Z_6));
    LocalMux I__427 (
            .O(N__2927),
            .I(beamYZ0Z_6));
    CascadeMux I__426 (
            .O(N__2918),
            .I(N__2912));
    InMux I__425 (
            .O(N__2917),
            .I(N__2909));
    InMux I__424 (
            .O(N__2916),
            .I(N__2904));
    InMux I__423 (
            .O(N__2915),
            .I(N__2904));
    InMux I__422 (
            .O(N__2912),
            .I(N__2901));
    LocalMux I__421 (
            .O(N__2909),
            .I(beamYZ0Z_5));
    LocalMux I__420 (
            .O(N__2904),
            .I(beamYZ0Z_5));
    LocalMux I__419 (
            .O(N__2901),
            .I(beamYZ0Z_5));
    CascadeMux I__418 (
            .O(N__2894),
            .I(un4_beamylt6_cascade_));
    CascadeMux I__417 (
            .O(N__2891),
            .I(un4_beamylt8_0_cascade_));
    CascadeMux I__416 (
            .O(N__2888),
            .I(N__2881));
    InMux I__415 (
            .O(N__2887),
            .I(N__2878));
    InMux I__414 (
            .O(N__2886),
            .I(N__2871));
    InMux I__413 (
            .O(N__2885),
            .I(N__2871));
    InMux I__412 (
            .O(N__2884),
            .I(N__2871));
    InMux I__411 (
            .O(N__2881),
            .I(N__2868));
    LocalMux I__410 (
            .O(N__2878),
            .I(beamYZ0Z_3));
    LocalMux I__409 (
            .O(N__2871),
            .I(beamYZ0Z_3));
    LocalMux I__408 (
            .O(N__2868),
            .I(beamYZ0Z_3));
    CascadeMux I__407 (
            .O(N__2861),
            .I(un1_beamylto9_2_cascade_));
    CascadeMux I__406 (
            .O(N__2858),
            .I(N__2851));
    InMux I__405 (
            .O(N__2857),
            .I(N__2848));
    InMux I__404 (
            .O(N__2856),
            .I(N__2841));
    InMux I__403 (
            .O(N__2855),
            .I(N__2841));
    InMux I__402 (
            .O(N__2854),
            .I(N__2841));
    InMux I__401 (
            .O(N__2851),
            .I(N__2838));
    LocalMux I__400 (
            .O(N__2848),
            .I(beamYZ0Z_4));
    LocalMux I__399 (
            .O(N__2841),
            .I(beamYZ0Z_4));
    LocalMux I__398 (
            .O(N__2838),
            .I(beamYZ0Z_4));
    IoInMux I__397 (
            .O(N__2831),
            .I(N__2828));
    LocalMux I__396 (
            .O(N__2828),
            .I(N__2825));
    IoSpan4Mux I__395 (
            .O(N__2825),
            .I(N__2822));
    Sp12to4 I__394 (
            .O(N__2822),
            .I(N__2818));
    IoInMux I__393 (
            .O(N__2821),
            .I(N__2815));
    Span12Mux_v I__392 (
            .O(N__2818),
            .I(N__2812));
    LocalMux I__391 (
            .O(N__2815),
            .I(N__2809));
    Odrv12 I__390 (
            .O(N__2812),
            .I(VSync_c));
    Odrv12 I__389 (
            .O(N__2809),
            .I(VSync_c));
    InMux I__388 (
            .O(N__2804),
            .I(N__2796));
    InMux I__387 (
            .O(N__2803),
            .I(N__2796));
    InMux I__386 (
            .O(N__2802),
            .I(N__2793));
    InMux I__385 (
            .O(N__2801),
            .I(N__2789));
    LocalMux I__384 (
            .O(N__2796),
            .I(N__2784));
    LocalMux I__383 (
            .O(N__2793),
            .I(N__2784));
    InMux I__382 (
            .O(N__2792),
            .I(N__2781));
    LocalMux I__381 (
            .O(N__2789),
            .I(beamYZ0Z_9));
    Odrv4 I__380 (
            .O(N__2784),
            .I(beamYZ0Z_9));
    LocalMux I__379 (
            .O(N__2781),
            .I(beamYZ0Z_9));
    CascadeMux I__378 (
            .O(N__2774),
            .I(N__2767));
    InMux I__377 (
            .O(N__2773),
            .I(N__2764));
    InMux I__376 (
            .O(N__2772),
            .I(N__2761));
    InMux I__375 (
            .O(N__2771),
            .I(N__2758));
    InMux I__374 (
            .O(N__2770),
            .I(N__2755));
    InMux I__373 (
            .O(N__2767),
            .I(N__2752));
    LocalMux I__372 (
            .O(N__2764),
            .I(beamYZ0Z_8));
    LocalMux I__371 (
            .O(N__2761),
            .I(beamYZ0Z_8));
    LocalMux I__370 (
            .O(N__2758),
            .I(beamYZ0Z_8));
    LocalMux I__369 (
            .O(N__2755),
            .I(beamYZ0Z_8));
    LocalMux I__368 (
            .O(N__2752),
            .I(beamYZ0Z_8));
    InMux I__367 (
            .O(N__2741),
            .I(un5_visibley_cry_2));
    InMux I__366 (
            .O(N__2738),
            .I(un5_visibley_cry_3));
    InMux I__365 (
            .O(N__2735),
            .I(un5_visibley_cry_4));
    InMux I__364 (
            .O(N__2732),
            .I(N__2728));
    InMux I__363 (
            .O(N__2731),
            .I(N__2725));
    LocalMux I__362 (
            .O(N__2728),
            .I(N__2722));
    LocalMux I__361 (
            .O(N__2725),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__360 (
            .O(N__2722),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    InMux I__359 (
            .O(N__2717),
            .I(un5_visibley_cry_5));
    CascadeMux I__358 (
            .O(N__2714),
            .I(N__2711));
    InMux I__357 (
            .O(N__2711),
            .I(N__2707));
    InMux I__356 (
            .O(N__2710),
            .I(N__2704));
    LocalMux I__355 (
            .O(N__2707),
            .I(N__2701));
    LocalMux I__354 (
            .O(N__2704),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    Odrv4 I__353 (
            .O(N__2701),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    InMux I__352 (
            .O(N__2696),
            .I(un5_visibley_cry_6));
    InMux I__351 (
            .O(N__2693),
            .I(N__2687));
    InMux I__350 (
            .O(N__2692),
            .I(N__2687));
    LocalMux I__349 (
            .O(N__2687),
            .I(un5_visibley_cry_7_c_RNI1L4CZ0));
    InMux I__348 (
            .O(N__2684),
            .I(un5_visibley_cry_7));
    InMux I__347 (
            .O(N__2681),
            .I(un5_visibley_cry_8));
    CascadeMux I__346 (
            .O(N__2678),
            .I(N__2675));
    InMux I__345 (
            .O(N__2675),
            .I(N__2669));
    InMux I__344 (
            .O(N__2674),
            .I(N__2669));
    LocalMux I__343 (
            .O(N__2669),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3));
    CEMux I__342 (
            .O(N__2666),
            .I(N__2661));
    InMux I__341 (
            .O(N__2665),
            .I(N__2656));
    InMux I__340 (
            .O(N__2664),
            .I(N__2653));
    LocalMux I__339 (
            .O(N__2661),
            .I(N__2650));
    CEMux I__338 (
            .O(N__2660),
            .I(N__2647));
    CEMux I__337 (
            .O(N__2659),
            .I(N__2643));
    LocalMux I__336 (
            .O(N__2656),
            .I(N__2634));
    LocalMux I__335 (
            .O(N__2653),
            .I(N__2634));
    Span4Mux_v I__334 (
            .O(N__2650),
            .I(N__2634));
    LocalMux I__333 (
            .O(N__2647),
            .I(N__2634));
    InMux I__332 (
            .O(N__2646),
            .I(N__2631));
    LocalMux I__331 (
            .O(N__2643),
            .I(N__2626));
    Span4Mux_v I__330 (
            .O(N__2634),
            .I(N__2626));
    LocalMux I__329 (
            .O(N__2631),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__328 (
            .O(N__2626),
            .I(beamX_RNI5457Z0Z_5));
    InMux I__327 (
            .O(N__2621),
            .I(un8_beamx_cry_9));
    InMux I__326 (
            .O(N__2618),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__325 (
            .O(N__2615),
            .I(N__2612));
    InMux I__324 (
            .O(N__2612),
            .I(N__2609));
    LocalMux I__323 (
            .O(N__2609),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0));
    InMux I__322 (
            .O(N__2606),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__321 (
            .O(N__2603),
            .I(N__2600));
    LocalMux I__320 (
            .O(N__2600),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0));
    InMux I__319 (
            .O(N__2597),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__318 (
            .O(N__2594),
            .I(N__2591));
    LocalMux I__317 (
            .O(N__2591),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0));
    CascadeMux I__316 (
            .O(N__2588),
            .I(N__2585));
    InMux I__315 (
            .O(N__2585),
            .I(N__2582));
    LocalMux I__314 (
            .O(N__2582),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__313 (
            .O(N__2579),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__312 (
            .O(N__2576),
            .I(N__2573));
    LocalMux I__311 (
            .O(N__2573),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    CascadeMux I__310 (
            .O(N__2570),
            .I(N__2565));
    InMux I__309 (
            .O(N__2569),
            .I(N__2562));
    InMux I__308 (
            .O(N__2568),
            .I(N__2559));
    InMux I__307 (
            .O(N__2565),
            .I(N__2556));
    LocalMux I__306 (
            .O(N__2562),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__305 (
            .O(N__2559),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__304 (
            .O(N__2556),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    CascadeMux I__303 (
            .O(N__2549),
            .I(N__2544));
    CascadeMux I__302 (
            .O(N__2548),
            .I(N__2541));
    CascadeMux I__301 (
            .O(N__2547),
            .I(N__2537));
    InMux I__300 (
            .O(N__2544),
            .I(N__2528));
    InMux I__299 (
            .O(N__2541),
            .I(N__2528));
    InMux I__298 (
            .O(N__2540),
            .I(N__2528));
    InMux I__297 (
            .O(N__2537),
            .I(N__2528));
    LocalMux I__296 (
            .O(N__2528),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0));
    InMux I__295 (
            .O(N__2525),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__294 (
            .O(N__2522),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_));
    InMux I__293 (
            .O(N__2519),
            .I(N__2516));
    LocalMux I__292 (
            .O(N__2516),
            .I(N__2513));
    Odrv4 I__291 (
            .O(N__2513),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__290 (
            .O(N__2510),
            .I(un8_beamx_cry_1));
    InMux I__289 (
            .O(N__2507),
            .I(un8_beamx_cry_2));
    InMux I__288 (
            .O(N__2504),
            .I(un8_beamx_cry_3));
    InMux I__287 (
            .O(N__2501),
            .I(un8_beamx_cry_4));
    InMux I__286 (
            .O(N__2498),
            .I(un8_beamx_cry_5));
    InMux I__285 (
            .O(N__2495),
            .I(un8_beamx_cry_6));
    InMux I__284 (
            .O(N__2492),
            .I(un8_beamx_cry_7));
    InMux I__283 (
            .O(N__2489),
            .I(bfn_7_8_0_));
    InMux I__282 (
            .O(N__2486),
            .I(bfn_7_5_0_));
    InMux I__281 (
            .O(N__2483),
            .I(N__2480));
    LocalMux I__280 (
            .O(N__2480),
            .I(N__2477));
    Odrv4 I__279 (
            .O(N__2477),
            .I(beamY_RNO_0Z0Z_9));
    CascadeMux I__278 (
            .O(N__2474),
            .I(un3_beamx_5_cascade_));
    InMux I__277 (
            .O(N__2471),
            .I(N__2468));
    LocalMux I__276 (
            .O(N__2468),
            .I(un3_beamx_7));
    InMux I__275 (
            .O(N__2465),
            .I(N__2462));
    LocalMux I__274 (
            .O(N__2462),
            .I(beamY_RNO_0Z0Z_1));
    CascadeMux I__273 (
            .O(N__2459),
            .I(N__2456));
    InMux I__272 (
            .O(N__2456),
            .I(N__2444));
    InMux I__271 (
            .O(N__2455),
            .I(N__2444));
    InMux I__270 (
            .O(N__2454),
            .I(N__2444));
    InMux I__269 (
            .O(N__2453),
            .I(N__2444));
    LocalMux I__268 (
            .O(N__2444),
            .I(N__2439));
    InMux I__267 (
            .O(N__2443),
            .I(N__2434));
    InMux I__266 (
            .O(N__2442),
            .I(N__2434));
    Odrv4 I__265 (
            .O(N__2439),
            .I(un5_beamx_3_0));
    LocalMux I__264 (
            .O(N__2434),
            .I(un5_beamx_3_0));
    CascadeMux I__263 (
            .O(N__2429),
            .I(N__2423));
    InMux I__262 (
            .O(N__2428),
            .I(N__2413));
    InMux I__261 (
            .O(N__2427),
            .I(N__2413));
    InMux I__260 (
            .O(N__2426),
            .I(N__2413));
    InMux I__259 (
            .O(N__2423),
            .I(N__2413));
    CascadeMux I__258 (
            .O(N__2422),
            .I(N__2410));
    LocalMux I__257 (
            .O(N__2413),
            .I(N__2406));
    InMux I__256 (
            .O(N__2410),
            .I(N__2401));
    InMux I__255 (
            .O(N__2409),
            .I(N__2401));
    Odrv4 I__254 (
            .O(N__2406),
            .I(un5_beamx_4));
    LocalMux I__253 (
            .O(N__2401),
            .I(un5_beamx_4));
    CascadeMux I__252 (
            .O(N__2396),
            .I(N__2392));
    CascadeMux I__251 (
            .O(N__2395),
            .I(N__2389));
    InMux I__250 (
            .O(N__2392),
            .I(N__2384));
    InMux I__249 (
            .O(N__2389),
            .I(N__2381));
    InMux I__248 (
            .O(N__2388),
            .I(N__2378));
    InMux I__247 (
            .O(N__2387),
            .I(N__2375));
    LocalMux I__246 (
            .O(N__2384),
            .I(N__2372));
    LocalMux I__245 (
            .O(N__2381),
            .I(beamYZ0Z_0));
    LocalMux I__244 (
            .O(N__2378),
            .I(beamYZ0Z_0));
    LocalMux I__243 (
            .O(N__2375),
            .I(beamYZ0Z_0));
    Odrv4 I__242 (
            .O(N__2372),
            .I(beamYZ0Z_0));
    InMux I__241 (
            .O(N__2363),
            .I(un21_beamy_cry_1));
    InMux I__240 (
            .O(N__2360),
            .I(N__2357));
    LocalMux I__239 (
            .O(N__2357),
            .I(beamY_RNO_0Z0Z_3));
    InMux I__238 (
            .O(N__2354),
            .I(un21_beamy_cry_2));
    CascadeMux I__237 (
            .O(N__2351),
            .I(N__2348));
    InMux I__236 (
            .O(N__2348),
            .I(N__2345));
    LocalMux I__235 (
            .O(N__2345),
            .I(beamY_RNO_0Z0Z_4));
    InMux I__234 (
            .O(N__2342),
            .I(un21_beamy_cry_3));
    InMux I__233 (
            .O(N__2339),
            .I(un21_beamy_cry_4));
    InMux I__232 (
            .O(N__2336),
            .I(un21_beamy_cry_5));
    CascadeMux I__231 (
            .O(N__2333),
            .I(N__2330));
    InMux I__230 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__229 (
            .O(N__2327),
            .I(beamY_RNO_0Z0Z_7));
    InMux I__228 (
            .O(N__2324),
            .I(un21_beamy_cry_6));
    InMux I__227 (
            .O(N__2321),
            .I(un21_beamy_cry_7));
    InMux I__226 (
            .O(N__2318),
            .I(N__2315));
    LocalMux I__225 (
            .O(N__2315),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0));
    InMux I__224 (
            .O(N__2312),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__223 (
            .O(N__2309),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__222 (
            .O(N__2306),
            .I(N__2303));
    LocalMux I__221 (
            .O(N__2303),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    CascadeMux I__220 (
            .O(N__2300),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    CascadeMux I__219 (
            .O(N__2297),
            .I(N__2294));
    InMux I__218 (
            .O(N__2294),
            .I(N__2291));
    LocalMux I__217 (
            .O(N__2291),
            .I(un5_visibley_cry_8_c_RNI3O5CZ0Z_0));
    InMux I__216 (
            .O(N__2288),
            .I(N__2285));
    LocalMux I__215 (
            .O(N__2285),
            .I(un5_visibley_cry_7_c_RNI1L4CZ0Z_0));
    InMux I__214 (
            .O(N__2282),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__213 (
            .O(N__2279),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__212 (
            .O(N__2276),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__211 (
            .O(N__2273),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__210 (
            .O(N__2270),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__209 (
            .O(N__2267),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_));
    InMux I__208 (
            .O(N__2264),
            .I(N__2261));
    LocalMux I__207 (
            .O(N__2261),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0));
    InMux I__206 (
            .O(N__2258),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2));
    IoInMux I__205 (
            .O(N__2255),
            .I(N__2252));
    LocalMux I__204 (
            .O(N__2252),
            .I(N__2249));
    Span4Mux_s1_h I__203 (
            .O(N__2249),
            .I(N__2246));
    Span4Mux_h I__202 (
            .O(N__2246),
            .I(N__2243));
    Sp12to4 I__201 (
            .O(N__2243),
            .I(N__2240));
    Odrv12 I__200 (
            .O(N__2240),
            .I(\Clock50MHz.PixelClock ));
    IoInMux I__199 (
            .O(N__2237),
            .I(N__2234));
    LocalMux I__198 (
            .O(N__2234),
            .I(N__2231));
    IoSpan4Mux I__197 (
            .O(N__2231),
            .I(N__2228));
    Odrv4 I__196 (
            .O(N__2228),
            .I(Clock12MHz_c));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_7_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_1_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__2255),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam beamY_RNO_0_1_LC_6_6_4.C_ON=1'b0;
    defparam beamY_RNO_0_1_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNO_0_1_LC_6_6_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamY_RNO_0_1_LC_6_6_4 (
            .in0(_gnd_net_),
            .in1(N__2388),
            .in2(_gnd_net_),
            .in3(N__4128),
            .lcout(beamY_RNO_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2714),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUC_LC_7_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUC_LC_7_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUC_LC_7_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUC_LC_7_1_1 (
            .in0(_gnd_net_),
            .in1(N__2288),
            .in2(N__4294),
            .in3(N__2282),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJN_LC_7_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJN_LC_7_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJN_LC_7_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJN_LC_7_1_2 (
            .in0(_gnd_net_),
            .in1(N__2264),
            .in2(N__4296),
            .in3(N__2279),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MN_LC_7_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MN_LC_7_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MN_LC_7_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MN_LC_7_1_3 (
            .in0(_gnd_net_),
            .in1(N__2318),
            .in2(N__4295),
            .in3(N__2276),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_1_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2570),
            .in3(N__2273),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(N__2306),
            .in2(_gnd_net_),
            .in3(N__2270),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2267),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(N__2692),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOM_LC_7_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOM_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOM_LC_7_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOM_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(N__4260),
            .in2(N__2297),
            .in3(N__2258),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPM_LC_7_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPM_LC_7_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPM_LC_7_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPM_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(N__4261),
            .in2(N__2678),
            .in3(N__2312),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2309),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2300),
            .in3(N__2569),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_7_2_5.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_0_LC_7_2_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_0_LC_7_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2674),
            .lcout(un5_visibley_cry_8_c_RNI3O5CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_7_2_6.C_ON=1'b0;
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_7_c_RNI1L4C_0_LC_7_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visibley_cry_7_c_RNI1L4C_0_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2693),
            .lcout(un5_visibley_cry_7_c_RNI1L4CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_2_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_2_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_2_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_7_LC_7_3_2.C_ON=1'b0;
    defparam beamY_7_LC_7_3_2.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_7_3_2.LUT_INIT=16'b0111000011110000;
    LogicCell40 beamY_7_LC_7_3_2 (
            .in0(N__2427),
            .in1(N__3081),
            .in2(N__2333),
            .in3(N__2455),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4053),
            .ce(N__2659),
            .sr(_gnd_net_));
    defparam beamY_3_LC_7_3_4.C_ON=1'b0;
    defparam beamY_3_LC_7_3_4.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_7_3_4.LUT_INIT=16'b0010101010101010;
    LogicCell40 beamY_3_LC_7_3_4 (
            .in0(N__2360),
            .in1(N__2453),
            .in2(N__2429),
            .in3(N__3079),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4053),
            .ce(N__2659),
            .sr(_gnd_net_));
    defparam beamY_4_LC_7_3_6.C_ON=1'b0;
    defparam beamY_4_LC_7_3_6.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_7_3_6.LUT_INIT=16'b0111000011110000;
    LogicCell40 beamY_4_LC_7_3_6 (
            .in0(N__2426),
            .in1(N__3080),
            .in2(N__2351),
            .in3(N__2454),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4053),
            .ce(N__2659),
            .sr(_gnd_net_));
    defparam beamY_9_LC_7_3_7.C_ON=1'b0;
    defparam beamY_9_LC_7_3_7.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_7_3_7.LUT_INIT=16'b0111111100000000;
    LogicCell40 beamY_9_LC_7_3_7 (
            .in0(N__3078),
            .in1(N__2428),
            .in2(N__2459),
            .in3(N__2483),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4053),
            .ce(N__2659),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_7_4_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_7_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(N__4146),
            .in2(N__2396),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_7_4_1.C_ON=1'b1;
    defparam beamY_2_LC_7_4_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_7_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_2_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(N__3041),
            .in2(_gnd_net_),
            .in3(N__2363),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(N__4052),
            .ce(N__2666),
            .sr(_gnd_net_));
    defparam beamY_RNO_0_3_LC_7_4_2.C_ON=1'b1;
    defparam beamY_RNO_0_3_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNO_0_3_LC_7_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNO_0_3_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__2887),
            .in2(_gnd_net_),
            .in3(N__2354),
            .lcout(beamY_RNO_0Z0Z_3),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNO_0_4_LC_7_4_3.C_ON=1'b1;
    defparam beamY_RNO_0_4_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNO_0_4_LC_7_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNO_0_4_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__2857),
            .in2(_gnd_net_),
            .in3(N__2342),
            .lcout(beamY_RNO_0Z0Z_4),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_5_LC_7_4_4.C_ON=1'b1;
    defparam beamY_5_LC_7_4_4.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_7_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(N__2917),
            .in2(_gnd_net_),
            .in3(N__2339),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(N__4052),
            .ce(N__2666),
            .sr(_gnd_net_));
    defparam beamY_6_LC_7_4_5.C_ON=1'b1;
    defparam beamY_6_LC_7_4_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_7_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_7_4_5 (
            .in0(_gnd_net_),
            .in1(N__2944),
            .in2(_gnd_net_),
            .in3(N__2336),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(N__4052),
            .ce(N__2666),
            .sr(_gnd_net_));
    defparam beamY_RNO_0_7_LC_7_4_6.C_ON=1'b1;
    defparam beamY_RNO_0_7_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNO_0_7_LC_7_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNO_0_7_LC_7_4_6 (
            .in0(_gnd_net_),
            .in1(N__3117),
            .in2(_gnd_net_),
            .in3(N__2324),
            .lcout(beamY_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_8_LC_7_4_7.C_ON=1'b1;
    defparam beamY_8_LC_7_4_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_7_4_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_7_4_7 (
            .in0(_gnd_net_),
            .in1(N__2772),
            .in2(_gnd_net_),
            .in3(N__2321),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(N__4052),
            .ce(N__2666),
            .sr(_gnd_net_));
    defparam beamY_RNO_0_9_LC_7_5_0.C_ON=1'b0;
    defparam beamY_RNO_0_9_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNO_0_9_LC_7_5_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 beamY_RNO_0_9_LC_7_5_0 (
            .in0(N__2803),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2486),
            .lcout(beamY_RNO_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_7_5_1.C_ON=1'b0;
    defparam beamX_0_LC_7_5_1.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_7_5_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_0_LC_7_5_1 (
            .in0(N__3001),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2646),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4050),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIA525_0_LC_7_5_2.C_ON=1'b0;
    defparam beamY_RNIA525_0_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIA525_0_LC_7_5_2.LUT_INIT=16'b0101000000000000;
    LogicCell40 beamY_RNIA525_0_LC_7_5_2 (
            .in0(N__2387),
            .in1(_gnd_net_),
            .in2(N__3152),
            .in3(N__3128),
            .lcout(un5_beamx_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_1_LC_7_5_3.C_ON=1'b0;
    defparam beamX_RNICPU5_1_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_1_LC_7_5_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNICPU5_1_LC_7_5_3 (
            .in0(N__3596),
            .in1(N__3233),
            .in2(N__3521),
            .in3(N__2968),
            .lcout(),
            .ltout(un3_beamx_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_0_LC_7_5_4.C_ON=1'b0;
    defparam beamX_RNIKVE6_0_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_0_LC_7_5_4.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNIKVE6_0_LC_7_5_4 (
            .in0(N__3556),
            .in1(N__3419),
            .in2(N__2474),
            .in3(N__3000),
            .lcout(un3_beamx_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_7_5_5.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_7_5_5.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_7_5_5.LUT_INIT=16'b0000001000000000;
    LogicCell40 beamX_RNI5457_5_LC_7_5_5 (
            .in0(N__2471),
            .in1(N__3458),
            .in2(N__3638),
            .in3(N__3323),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC725_9_LC_7_5_7.C_ON=1'b0;
    defparam beamY_RNIC725_9_LC_7_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIC725_9_LC_7_5_7.LUT_INIT=16'b0000001000000000;
    LogicCell40 beamY_RNIC725_9_LC_7_5_7 (
            .in0(N__4141),
            .in1(N__2773),
            .in2(N__3047),
            .in3(N__2804),
            .lcout(un5_beamx_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_7_6_1.C_ON=1'b0;
    defparam beamY_1_LC_7_6_1.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_7_6_1.LUT_INIT=16'b0100110011001100;
    LogicCell40 beamY_1_LC_7_6_1 (
            .in0(N__3082),
            .in1(N__2465),
            .in2(N__2422),
            .in3(N__2443),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4048),
            .ce(N__2660),
            .sr(_gnd_net_));
    defparam beamY_0_LC_7_6_4.C_ON=1'b0;
    defparam beamY_0_LC_7_6_4.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_7_6_4.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamY_0_LC_7_6_4 (
            .in0(N__2442),
            .in1(N__2409),
            .in2(N__2395),
            .in3(N__3083),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4048),
            .ce(N__2660),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_7_7_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_7_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__3005),
            .in2(N__2972),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_7_7_1.C_ON=1'b1;
    defparam beamX_2_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_7_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__3230),
            .in2(_gnd_net_),
            .in3(N__2510),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_7_7_2.C_ON=1'b1;
    defparam beamX_3_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_7_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(N__3551),
            .in2(_gnd_net_),
            .in3(N__2507),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_7_7_3.C_ON=1'b1;
    defparam beamX_4_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_7_7_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_7_7_3 (
            .in0(N__2664),
            .in1(N__3592),
            .in2(_gnd_net_),
            .in3(N__2504),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_7_7_4.C_ON=1'b1;
    defparam beamX_5_LC_7_7_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_7_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__3631),
            .in2(_gnd_net_),
            .in3(N__2501),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_7_7_5.C_ON=1'b1;
    defparam beamX_6_LC_7_7_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_7_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(N__3410),
            .in2(_gnd_net_),
            .in3(N__2498),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_7_7_6.C_ON=1'b1;
    defparam beamX_7_LC_7_7_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_7_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_7_7_6 (
            .in0(_gnd_net_),
            .in1(N__3453),
            .in2(_gnd_net_),
            .in3(N__2495),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_7_7_7.C_ON=1'b1;
    defparam beamX_8_LC_7_7_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_7_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(N__3365),
            .in2(_gnd_net_),
            .in3(N__2492),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__4047),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_7_8_0.C_ON=1'b1;
    defparam beamX_9_LC_7_8_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_7_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__3343),
            .in2(_gnd_net_),
            .in3(N__2489),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__4046),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_7_8_1.C_ON=1'b0;
    defparam beamX_10_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_7_8_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_10_LC_7_8_1 (
            .in0(N__2665),
            .in1(N__3506),
            .in2(_gnd_net_),
            .in3(N__2621),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4046),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_1_0 (
            .in0(_gnd_net_),
            .in1(N__2732),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_1_1 (
            .in0(_gnd_net_),
            .in1(N__2519),
            .in2(N__2547),
            .in3(N__2618),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5UR_LC_8_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5UR_LC_8_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5UR_LC_8_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5UR_LC_8_1_2 (
            .in0(_gnd_net_),
            .in1(N__2540),
            .in2(N__2615),
            .in3(N__2606),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9K61_LC_8_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9K61_LC_8_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9K61_LC_8_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9K61_LC_8_1_3 (
            .in0(_gnd_net_),
            .in1(N__2603),
            .in2(N__2548),
            .in3(N__2597),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIVBNM1_LC_8_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIVBNM1_LC_8_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIVBNM1_LC_8_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIVBNM1_LC_8_1_4 (
            .in0(N__3275),
            .in1(N__2594),
            .in2(N__2588),
            .in3(N__2579),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_1_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_1_5 (
            .in0(N__2576),
            .in1(N__2568),
            .in2(N__2549),
            .in3(N__2525),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_8_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_8_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_8_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_8_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2522),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_2_2.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_2_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2710),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_8_2_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_8_2_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_8_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2731),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_2_c_LC_8_3_0.C_ON=1'b1;
    defparam un5_visibley_cry_2_c_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_2_c_LC_8_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visibley_cry_2_c_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3046),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(un5_visibley_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_3_1.C_ON=1'b1;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_2_c_RNIN5VB_LC_8_3_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_2_c_RNIN5VB_LC_8_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2888),
            .in3(N__2741),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visibley_cry_2),
            .carryout(un5_visibley_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_3_2.C_ON=1'b1;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_3_c_RNIP80C_LC_8_3_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visibley_cry_3_c_RNIP80C_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2858),
            .in3(N__2738),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visibley_cry_3),
            .carryout(un5_visibley_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_3_3.C_ON=1'b1;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_4_c_RNIRB1C_LC_8_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_4_c_RNIRB1C_LC_8_3_3 (
            .in0(_gnd_net_),
            .in1(N__4297),
            .in2(N__2918),
            .in3(N__2735),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visibley_cry_4),
            .carryout(un5_visibley_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_3_4.C_ON=1'b1;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_5_c_RNITE2C_LC_8_3_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_5_c_RNITE2C_LC_8_3_4 (
            .in0(_gnd_net_),
            .in1(N__4289),
            .in2(N__2945),
            .in3(N__2717),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visibley_cry_5),
            .carryout(un5_visibley_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_3_5.C_ON=1'b1;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_6_c_RNIVH3C_LC_8_3_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_6_c_RNIVH3C_LC_8_3_5 (
            .in0(_gnd_net_),
            .in1(N__4298),
            .in2(N__3120),
            .in3(N__2696),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visibley_cry_6),
            .carryout(un5_visibley_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_3_6.C_ON=1'b1;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_7_c_RNI1L4C_LC_8_3_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visibley_cry_7_c_RNI1L4C_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(N__4290),
            .in2(N__2774),
            .in3(N__2684),
            .lcout(un5_visibley_cry_7_c_RNI1L4CZ0),
            .ltout(),
            .carryin(un5_visibley_cry_7),
            .carryout(un5_visibley_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_3_7.C_ON=1'b0;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam un5_visibley_cry_8_c_RNI3O5C_LC_8_3_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visibley_cry_8_c_RNI3O5C_LC_8_3_7 (
            .in0(_gnd_net_),
            .in1(N__2792),
            .in2(_gnd_net_),
            .in3(N__2681),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_axb_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_4_0.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_4_0.LUT_INIT=16'b0011001100110011;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_4_0 (
            .in0(N__4299),
            .in1(N__3038),
            .in2(_gnd_net_),
            .in3(N__4177),
            .lcout(un5_visibley_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4H2_5_LC_8_4_1.C_ON=1'b0;
    defparam beamY_RNIN4H2_5_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4H2_5_LC_8_4_1.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIN4H2_5_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__2942),
            .in2(_gnd_net_),
            .in3(N__2915),
            .lcout(un1_beamy_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_18_LC_8_4_2.C_ON=1'b0;
    defparam Pixel_1_RNO_18_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_18_LC_8_4_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 Pixel_1_RNO_18_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(N__3039),
            .in2(_gnd_net_),
            .in3(N__2884),
            .lcout(),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_14_LC_8_4_3.C_ON=1'b0;
    defparam Pixel_1_RNO_14_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_14_LC_8_4_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_14_LC_8_4_3 (
            .in0(N__2943),
            .in1(N__2916),
            .in2(N__2894),
            .in3(N__2855),
            .lcout(),
            .ltout(un4_beamylt8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_5_LC_8_4_4.C_ON=1'b0;
    defparam Pixel_1_RNO_5_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_5_LC_8_4_4.LUT_INIT=16'b1010101010101000;
    LogicCell40 Pixel_1_RNO_5_LC_8_4_4 (
            .in0(N__2801),
            .in1(N__2771),
            .in2(N__2891),
            .in3(N__3118),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0H2_3_LC_8_4_5.C_ON=1'b0;
    defparam beamY_RNIJ0H2_3_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0H2_3_LC_8_4_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 beamY_RNIJ0H2_3_LC_8_4_5 (
            .in0(N__2885),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2854),
            .lcout(un5_beamx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_RNO_0_LC_8_4_6.C_ON=1'b0;
    defparam VSync_1_RNO_0_LC_8_4_6.SEQ_MODE=4'b0000;
    defparam VSync_1_RNO_0_LC_8_4_6.LUT_INIT=16'b0000000000010101;
    LogicCell40 VSync_1_RNO_0_LC_8_4_6 (
            .in0(N__3119),
            .in1(N__3040),
            .in2(N__4151),
            .in3(N__2886),
            .lcout(),
            .ltout(un1_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_8_4_7.C_ON=1'b0;
    defparam VSync_1_LC_8_4_7.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_8_4_7.LUT_INIT=16'b1111111101111111;
    LogicCell40 VSync_1_LC_8_4_7 (
            .in0(N__3167),
            .in1(N__3150),
            .in2(N__2861),
            .in3(N__2856),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4054),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITAH2_9_LC_8_5_0.C_ON=1'b0;
    defparam beamY_RNITAH2_9_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNITAH2_9_LC_8_5_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNITAH2_9_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(N__2802),
            .in2(_gnd_net_),
            .in3(N__2770),
            .lcout(un8_beamy_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_7_LC_8_5_1.C_ON=1'b0;
    defparam Pixel_1_RNO_7_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_7_LC_8_5_1.LUT_INIT=16'b1101000011000000;
    LogicCell40 Pixel_1_RNO_7_LC_8_5_1 (
            .in0(N__3179),
            .in1(N__3634),
            .in2(N__3377),
            .in3(N__3595),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_8_5_2.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_8_5_2.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamX_RNIQCL_1_LC_8_5_2 (
            .in0(N__2967),
            .in1(N__2999),
            .in2(N__3557),
            .in3(N__3232),
            .lcout(un18_beamylt4),
            .ltout(un18_beamylt4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_15_LC_8_5_3.C_ON=1'b0;
    defparam Pixel_1_RNO_15_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_15_LC_8_5_3.LUT_INIT=16'b0101000101010101;
    LogicCell40 Pixel_1_RNO_15_LC_8_5_3 (
            .in0(N__3418),
            .in1(N__3633),
            .in2(N__3173),
            .in3(N__3594),
            .lcout(),
            .ltout(un13_beamylt7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_6_LC_8_5_4.C_ON=1'b0;
    defparam Pixel_1_RNO_6_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_6_LC_8_5_4.LUT_INIT=16'b0100000001000100;
    LogicCell40 Pixel_1_RNO_6_LC_8_5_4 (
            .in0(N__3520),
            .in1(N__3322),
            .in2(N__3170),
            .in3(N__3457),
            .lcout(un13_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_13_LC_8_5_5.C_ON=1'b0;
    defparam Pixel_1_RNO_13_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_13_LC_8_5_5.LUT_INIT=16'b0000000010001000;
    LogicCell40 Pixel_1_RNO_13_LC_8_5_5 (
            .in0(N__3163),
            .in1(N__3151),
            .in2(_gnd_net_),
            .in3(N__3127),
            .lcout(),
            .ltout(un8_beamylto9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_4_LC_8_5_6.C_ON=1'b0;
    defparam Pixel_1_RNO_4_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_4_LC_8_5_6.LUT_INIT=16'b0100010100000101;
    LogicCell40 Pixel_1_RNO_4_LC_8_5_6 (
            .in0(N__3519),
            .in1(N__3072),
            .in2(N__3050),
            .in3(N__3042),
            .lcout(Pixel_0_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_8_6_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__2997),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_8_6_1.C_ON=1'b1;
    defparam beamX_1_LC_8_6_1.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_8_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_1_LC_8_6_1 (
            .in0(N__2998),
            .in1(N__2966),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(N__4051),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_LC_8_6_2.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_LC_8_6_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_2_c_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(N__3231),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_9_LC_8_6_3.C_ON=1'b1;
    defparam Pixel_1_RNO_9_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_9_LC_8_6_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_9_LC_8_6_3 (
            .in0(_gnd_net_),
            .in1(N__3544),
            .in2(N__4330),
            .in3(N__3203),
            .lcout(un1_visiblex_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_6_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_8_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(N__3583),
            .in2(_gnd_net_),
            .in3(N__3200),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_6_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_8_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(N__3622),
            .in2(_gnd_net_),
            .in3(N__3197),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_6_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_8_6_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(N__3400),
            .in2(N__4331),
            .in3(N__3194),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_6_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_8_6_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_8_6_7 (
            .in0(_gnd_net_),
            .in1(N__3447),
            .in2(_gnd_net_),
            .in3(N__3191),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_7_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_8_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(N__3362),
            .in2(N__4332),
            .in3(N__3188),
            .lcout(un5_visiblex_cry_7_c_RNIVZ0Z952),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_7_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_8_7_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(N__3338),
            .in2(_gnd_net_),
            .in3(N__3185),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_c5),
            .ltout(un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_7_2.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_8_7_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3182),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_RNO_0_LC_8_7_3.C_ON=1'b0;
    defparam HSync_1_RNO_0_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam HSync_1_RNO_0_LC_8_7_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 HSync_1_RNO_0_LC_8_7_3 (
            .in0(N__3632),
            .in1(N__3593),
            .in2(N__3411),
            .in3(N__3552),
            .lcout(),
            .ltout(un1_beamxlt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_8_7_4.C_ON=1'b0;
    defparam HSync_1_LC_8_7_4.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_8_7_4.LUT_INIT=16'b1111111111111011;
    LogicCell40 HSync_1_LC_8_7_4 (
            .in0(N__3507),
            .in1(N__3321),
            .in2(N__3485),
            .in3(N__3449),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4049),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_16_LC_8_7_6.C_ON=1'b0;
    defparam Pixel_1_RNO_16_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_16_LC_8_7_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 Pixel_1_RNO_16_LC_8_7_6 (
            .in0(N__3364),
            .in1(N__3448),
            .in2(N__3344),
            .in3(N__3401),
            .lcout(un18_beamylto9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_8_7_7.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_8_7_7.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_RNIR4B_9_LC_8_7_7 (
            .in0(N__3363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3339),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_1_0 (
            .in0(_gnd_net_),
            .in1(N__3833),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_9_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_9_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_9_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_9_1_1 (
            .in0(_gnd_net_),
            .in1(N__3276),
            .in2(N__3302),
            .in3(N__3293),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_9_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_9_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_9_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(N__3290),
            .in2(N__3281),
            .in3(N__3284),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8IL1_LC_9_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8IL1_LC_9_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8IL1_LC_9_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8IL1_LC_9_1_3 (
            .in0(_gnd_net_),
            .in1(N__3280),
            .in2(N__3260),
            .in3(N__3251),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ5N04_LC_9_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ5N04_LC_9_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ5N04_LC_9_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ5N04_LC_9_1_4 (
            .in0(N__3692),
            .in1(N__3248),
            .in2(N__3242),
            .in3(N__3725),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_LC_9_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_LC_9_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_LC_9_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_LC_9_1_5 (
            .in0(_gnd_net_),
            .in1(N__3722),
            .in2(_gnd_net_),
            .in3(N__3716),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02),
            .ltout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_0_LC_9_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_0_LC_9_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_0_LC_9_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_0_LC_9_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3713),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_9_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_9_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_9_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_9_2_0 (
            .in0(_gnd_net_),
            .in1(N__3946),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFR2_LC_9_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFR2_LC_9_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFR2_LC_9_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFR2_LC_9_2_1 (
            .in0(_gnd_net_),
            .in1(N__3693),
            .in2(N__3818),
            .in3(N__3710),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6B3_LC_9_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6B3_LC_9_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6B3_LC_9_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6B3_LC_9_2_2 (
            .in0(_gnd_net_),
            .in1(N__3707),
            .in2(N__3698),
            .in3(N__3701),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3R3_LC_9_2_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3R3_LC_9_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3R3_LC_9_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3R3_LC_9_2_3 (
            .in0(_gnd_net_),
            .in1(N__3697),
            .in2(N__3677),
            .in3(N__3668),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHBHM8_LC_9_2_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHBHM8_LC_9_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHBHM8_LC_9_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHBHM8_LC_9_2_4 (
            .in0(N__3791),
            .in1(N__3665),
            .in2(N__3659),
            .in3(N__3650),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_LC_9_2_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_LC_9_2_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_LC_9_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_LC_9_2_5 (
            .in0(_gnd_net_),
            .in1(N__3647),
            .in2(_gnd_net_),
            .in3(N__3641),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4),
            .ltout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_0_LC_9_2_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_0_LC_9_2_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_0_LC_9_2_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_0_LC_9_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3836),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_2_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_2_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3832),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_3_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3O4_LC_9_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3O4_LC_9_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3O4_LC_9_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3O4_LC_9_3_1 (
            .in0(_gnd_net_),
            .in1(N__3792),
            .in2(N__3935),
            .in3(N__3809),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFE7_LC_9_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFE7_LC_9_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFE7_LC_9_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFE7_LC_9_3_2 (
            .in0(_gnd_net_),
            .in1(N__3806),
            .in2(N__3797),
            .in3(N__3800),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7U7_LC_9_3_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7U7_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7U7_LC_9_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7U7_LC_9_3_3 (
            .in0(_gnd_net_),
            .in1(N__3796),
            .in2(N__3776),
            .in3(N__3767),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIS657H_LC_9_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIS657H_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIS657H_LC_9_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIS657H_LC_9_3_4 (
            .in0(N__3888),
            .in1(N__3764),
            .in2(N__3758),
            .in3(N__3749),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVO8_LC_9_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVO8_LC_9_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVO8_LC_9_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVO8_LC_9_3_5 (
            .in0(_gnd_net_),
            .in1(N__3746),
            .in2(_gnd_net_),
            .in3(N__3740),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_9_3_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_9_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_9_3_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_9_3_6 (
            .in0(N__3736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_9_3_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_9_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_9_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_9_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3947),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_17_LC_9_4_0.C_ON=1'b1;
    defparam Pixel_1_RNO_17_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_17_LC_9_4_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 Pixel_1_RNO_17_LC_9_4_0 (
            .in0(_gnd_net_),
            .in1(N__4173),
            .in2(_gnd_net_),
            .in3(N__4145),
            .lcout(G_6_i_a4_0_0),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFP59_LC_9_4_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFP59_LC_9_4_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFP59_LC_9_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFP59_LC_9_4_1 (
            .in0(_gnd_net_),
            .in1(N__3926),
            .in2(N__3889),
            .in3(N__3920),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPD_LC_9_4_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPD_LC_9_4_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPD_LC_9_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPD_LC_9_4_2 (
            .in0(_gnd_net_),
            .in1(N__3884),
            .in2(N__3917),
            .in3(N__3908),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_12_LC_9_4_3.C_ON=1'b1;
    defparam Pixel_1_RNO_12_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_12_LC_9_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_12_LC_9_4_3 (
            .in0(_gnd_net_),
            .in1(N__3905),
            .in2(N__3890),
            .in3(N__3899),
            .lcout(Pixel_1_RNOZ0Z_12),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_4_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_4_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(N__3896),
            .in2(N__3863),
            .in3(N__3880),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFH_LC_9_4_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFH_LC_9_4_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFH_LC_9_4_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFH_LC_9_4_5 (
            .in0(_gnd_net_),
            .in1(N__3854),
            .in2(_gnd_net_),
            .in3(N__3848),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_11_LC_9_4_6.C_ON=1'b0;
    defparam Pixel_1_RNO_11_LC_9_4_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_11_LC_9_4_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_11_LC_9_4_6 (
            .in0(N__3845),
            .in1(N__4202),
            .in2(N__3839),
            .in3(N__4190),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_10_LC_9_5_2.C_ON=1'b0;
    defparam Pixel_1_RNO_10_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_10_LC_9_5_2.LUT_INIT=16'b1110111111111111;
    LogicCell40 Pixel_1_RNO_10_LC_9_5_2 (
            .in0(N__4201),
            .in1(N__4189),
            .in2(N__4178),
            .in3(N__4157),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_3_LC_9_5_3.C_ON=1'b0;
    defparam Pixel_1_RNO_3_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_3_LC_9_5_3.LUT_INIT=16'b0000000000110100;
    LogicCell40 Pixel_1_RNO_3_LC_9_5_3 (
            .in0(N__4150),
            .in1(N__4100),
            .in2(N__4094),
            .in3(N__4091),
            .lcout(),
            .ltout(un15_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_9_5_4.C_ON=1'b0;
    defparam Pixel_1_LC_9_5_4.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_9_5_4.LUT_INIT=16'b1100000010000100;
    LogicCell40 Pixel_1_LC_9_5_4 (
            .in0(N__3956),
            .in1(N__3986),
            .in2(N__4085),
            .in3(N__3965),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4055),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_0_LC_9_5_6.C_ON=1'b0;
    defparam Pixel_1_RNO_0_LC_9_5_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_0_LC_9_5_6.LUT_INIT=16'b0000000100000000;
    LogicCell40 Pixel_1_RNO_0_LC_9_5_6 (
            .in0(N__4019),
            .in1(N__4013),
            .in2(N__4007),
            .in3(N__3995),
            .lcout(Pixel_0_sqmuxa_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_7_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_9_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4530),
            .lcout(un5_visiblex_cry_8_c_RNI1D62Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_2_LC_11_5_1.C_ON=1'b0;
    defparam Pixel_1_RNO_2_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_2_LC_11_5_1.LUT_INIT=16'b1001100010100010;
    LogicCell40 Pixel_1_RNO_2_LC_11_5_1 (
            .in0(N__4418),
            .in1(N__4450),
            .in2(N__3980),
            .in3(N__4634),
            .lcout(un14lt10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_1_LC_11_5_5.C_ON=1'b0;
    defparam Pixel_1_RNO_1_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_1_LC_11_5_5.LUT_INIT=16'b0011100111001100;
    LogicCell40 Pixel_1_RNO_1_LC_11_5_5 (
            .in0(N__4417),
            .in1(N__4406),
            .in2(N__4451),
            .in3(N__4633),
            .lcout(un1_visiblex_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_11_6_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_11_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__4381),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_11_6_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_11_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__4502),
            .in2(N__4460),
            .in3(N__4397),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_11_6_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_11_6_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_11_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(N__4492),
            .in2(N__4358),
            .in3(N__4394),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_11_6_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_11_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_11_6_3 (
            .in0(N__4691),
            .in1(N__4478),
            .in2(N__4214),
            .in3(N__4391),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_11_6_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_11_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_11_6_4 (
            .in0(N__4493),
            .in1(N__4541),
            .in2(N__4517),
            .in3(N__4388),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31),
            .ltout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_11_6_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_11_6_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_11_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4385),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_11_6_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_11_6_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_11_6_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_11_6_7 (
            .in0(N__4382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_7_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(N__4471),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_11_7_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_11_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__4367),
            .in2(_gnd_net_),
            .in3(N__4349),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_11_7_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_11_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__4346),
            .in2(N__4337),
            .in3(N__4205),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_7_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_7_3 (
            .in0(_gnd_net_),
            .in1(N__4537),
            .in2(_gnd_net_),
            .in3(N__4508),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_7_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4505),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO),
            .ltout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_11_7_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_11_7_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_11_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_11_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4496),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0),
            .ltout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_11_7_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_11_7_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_11_7_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_11_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4481),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_11_7_7.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_11_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_11_7_7 (
            .in0(N__4472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_visiblex_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_12_4_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_12_4_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_12_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(N__4446),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_12_4_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_12_4_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_12_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__4645),
            .in2(N__4625),
            .in3(N__4409),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_8_LC_12_4_2.C_ON=1'b1;
    defparam Pixel_1_RNO_8_LC_12_4_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_8_LC_12_4_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_8_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(N__4592),
            .in2(N__4559),
            .in3(N__4400),
            .lcout(Pixel_1_RNOZ0Z_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_12_4_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_12_4_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_12_4_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(N__4646),
            .in2(N__4583),
            .in3(N__4554),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PB_LC_12_4_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PB_LC_12_4_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PB_LC_12_4_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PB_LC_12_4_4 (
            .in0(_gnd_net_),
            .in1(N__4571),
            .in2(_gnd_net_),
            .in3(N__4637),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_12_4_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_12_4_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_12_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4616),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_12_5_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_12_5_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_12_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_12_5_0 (
            .in0(_gnd_net_),
            .in1(N__4615),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_12_5_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_12_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(N__4711),
            .in2(N__4655),
            .in3(N__4586),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_12_5_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_12_5_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_12_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_12_5_2 (
            .in0(_gnd_net_),
            .in1(N__4727),
            .in2(N__4778),
            .in3(N__4574),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGQELB_LC_12_5_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGQELB_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGQELB_LC_12_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGQELB_LC_12_5_3 (
            .in0(N__4558),
            .in1(N__4712),
            .in2(N__4757),
            .in3(N__4565),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJ6_LC_12_5_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJ6_LC_12_5_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJ6_LC_12_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJ6_LC_12_5_4 (
            .in0(_gnd_net_),
            .in1(N__4745),
            .in2(_gnd_net_),
            .in3(N__4562),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_12_6_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_12_6_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_12_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_12_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_12_6_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_12_6_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_12_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_12_6_1 (
            .in0(_gnd_net_),
            .in1(N__4793),
            .in2(N__4787),
            .in3(N__4769),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_12_6_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_12_6_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_12_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_12_6_2 (
            .in0(_gnd_net_),
            .in1(N__4690),
            .in2(N__4766),
            .in3(N__4748),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNIEN766_LC_12_6_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNIEN766_LC_12_6_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNIEN766_LC_12_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNIEN766_LC_12_6_3 (
            .in0(N__4726),
            .in1(N__4676),
            .in2(N__4703),
            .in3(N__4739),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_12_6_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_12_6_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_12_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_12_6_4 (
            .in0(_gnd_net_),
            .in1(N__4736),
            .in2(_gnd_net_),
            .in3(N__4730),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2),
            .ltout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_12_6_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_12_6_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_12_6_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_12_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4715),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKL62_LC_12_6_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKL62_LC_12_6_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKL62_LC_12_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKL62_LC_12_6_6 (
            .in0(_gnd_net_),
            .in1(N__4702),
            .in2(_gnd_net_),
            .in3(N__4689),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_12_6_7.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_12_6_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_12_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_12_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4669),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
